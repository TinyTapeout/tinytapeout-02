* NGSPICE file created from user_project_wrapper.ext - technology: sky130B

* Black-box entry subcircuit for user_module_347688030570545747 abstract view
.subckt user_module_347688030570545747 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_339501025136214612 abstract view
.subckt user_module_339501025136214612 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for scanchain abstract view
.subckt scanchain clk_in clk_out data_in data_out latch_enable_in latch_enable_out
+ module_data_in[0] module_data_in[1] module_data_in[2] module_data_in[3] module_data_in[4]
+ module_data_in[5] module_data_in[6] module_data_in[7] module_data_out[0] module_data_out[1]
+ module_data_out[2] module_data_out[3] module_data_out[4] module_data_out[5] module_data_out[6]
+ module_data_out[7] scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for alu_top abstract view
.subckt alu_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for migcorre_pwm abstract view
.subckt migcorre_pwm io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347894637149553236 abstract view
.subckt user_module_347894637149553236 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for azdle_binary_clock abstract view
.subckt azdle_binary_clock io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for phasenoisepon_seven_segment_seconds abstract view
.subckt phasenoisepon_seven_segment_seconds io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for jar_sram_top abstract view
.subckt jar_sram_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341620484740219475 abstract view
.subckt user_module_341620484740219475 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for xor_shift32_evango abstract view
.subckt xor_shift32_evango io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for rc5_top abstract view
.subckt rc5_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for tt2_tholin_multiplier abstract view
.subckt tt2_tholin_multiplier io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_346916357828248146 abstract view
.subckt user_module_346916357828248146 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for chrisruk_matrix abstract view
.subckt chrisruk_matrix io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for yubex_egg_timer abstract view
.subckt yubex_egg_timer io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347619669052490324 abstract view
.subckt user_module_347619669052490324 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348121131386929746 abstract view
.subckt user_module_348121131386929746 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt2_tholin_multiplexed_counter abstract view
.subckt tt2_tholin_multiplexed_counter io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for jleightcap_top abstract view
.subckt jleightcap_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348195845106041428 abstract view
.subckt user_module_348195845106041428 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for xor_shift32_quantamhd abstract view
.subckt xor_shift32_quantamhd io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for mbikovitsky_top abstract view
.subckt mbikovitsky_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for meriac_tt02_play_tune abstract view
.subckt meriac_tt02_play_tune io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347690870424732244 abstract view
.subckt user_module_347690870424732244 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tholin_avalonsemi_5401 abstract view
.subckt tholin_avalonsemi_5401 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for mm21_LEDMatrixTop abstract view
.subckt mm21_LEDMatrixTop io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_346553315158393428 abstract view
.subckt user_module_346553315158393428 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341541108650607187 abstract view
.subckt user_module_341541108650607187 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tholin_avalonsemi_tbb1143 abstract view
.subckt tholin_avalonsemi_tbb1143 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tomkeddie_top_tto_a abstract view
.subckt tomkeddie_top_tto_a io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for top abstract view
.subckt top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348242239268323922 abstract view
.subckt user_module_348242239268323922 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for moyes0_top_module abstract view
.subckt moyes0_top_module io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for flygoat_tt02_play_tune abstract view
.subckt flygoat_tt02_play_tune io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348260124451668562 abstract view
.subckt user_module_348260124451668562 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tiny_fft abstract view
.subckt tiny_fft io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for tt2_tholin_namebadge abstract view
.subckt tt2_tholin_namebadge io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tomkeddie_top_tto abstract view
.subckt tomkeddie_top_tto io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for zoechip abstract view
.subckt zoechip io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for thezoq2_yafpga abstract view
.subckt thezoq2_yafpga io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347594509754827347 abstract view
.subckt user_module_347594509754827347 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for s4ga abstract view
.subckt s4ga io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for asic_multiplier_wrapper abstract view
.subckt asic_multiplier_wrapper io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for loxodes_sequencer abstract view
.subckt loxodes_sequencer io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for jar_illegal_logic abstract view
.subckt jar_illegal_logic io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for aidan_McCoy abstract view
.subckt aidan_McCoy io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341516949939814994 abstract view
.subckt user_module_341516949939814994 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for rolfmobile99_alu_fsm_top abstract view
.subckt rolfmobile99_alu_fsm_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341614374571475540 abstract view
.subckt user_module_341614374571475540 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347787021138264660 abstract view
.subckt user_module_347787021138264660 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_controller abstract view
.subckt scan_controller active_select[0] active_select[1] active_select[2] active_select[3]
+ active_select[4] active_select[5] active_select[6] active_select[7] active_select[8]
+ clk driver_sel[0] driver_sel[1] inputs[0] inputs[1] inputs[2] inputs[3] inputs[4]
+ inputs[5] inputs[6] inputs[7] la_scan_clk_in la_scan_data_in la_scan_data_out la_scan_latch_en
+ la_scan_select oeb[0] oeb[10] oeb[11] oeb[12] oeb[13] oeb[14] oeb[15] oeb[16] oeb[17]
+ oeb[18] oeb[19] oeb[1] oeb[20] oeb[21] oeb[22] oeb[23] oeb[24] oeb[25] oeb[26] oeb[27]
+ oeb[28] oeb[29] oeb[2] oeb[30] oeb[31] oeb[32] oeb[33] oeb[34] oeb[35] oeb[36] oeb[37]
+ oeb[3] oeb[4] oeb[5] oeb[6] oeb[7] oeb[8] oeb[9] outputs[0] outputs[1] outputs[2]
+ outputs[3] outputs[4] outputs[5] outputs[6] outputs[7] ready reset scan_clk_in scan_clk_out
+ scan_data_in scan_data_out scan_latch_en scan_select set_clk_div slow_clk vccd1
+ vssd1
.ends

* Black-box entry subcircuit for yupferris_bitslam abstract view
.subckt yupferris_bitslam io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for xyz_peppergray_Potato1_top abstract view
.subckt xyz_peppergray_Potato1_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for chase_the_beat abstract view
.subckt chase_the_beat io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_342981109408072274 abstract view
.subckt user_module_342981109408072274 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348255968419643987 abstract view
.subckt user_module_348255968419643987 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347592305412145748 abstract view
.subckt user_module_347592305412145748 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for fraserbc_simon abstract view
.subckt fraserbc_simon io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xuser_module_347688030570545747_21 scanchain_21/module_data_in[0] scanchain_21/module_data_in[1]
+ scanchain_21/module_data_in[2] scanchain_21/module_data_in[3] scanchain_21/module_data_in[4]
+ scanchain_21/module_data_in[5] scanchain_21/module_data_in[6] scanchain_21/module_data_in[7]
+ scanchain_21/module_data_out[0] scanchain_21/module_data_out[1] scanchain_21/module_data_out[2]
+ scanchain_21/module_data_out[3] scanchain_21/module_data_out[4] scanchain_21/module_data_out[5]
+ scanchain_21/module_data_out[6] scanchain_21/module_data_out[7] vccd1 vssd1 user_module_347688030570545747
Xuser_module_339501025136214612_59 scanchain_59/module_data_in[0] scanchain_59/module_data_in[1]
+ scanchain_59/module_data_in[2] scanchain_59/module_data_in[3] scanchain_59/module_data_in[4]
+ scanchain_59/module_data_in[5] scanchain_59/module_data_in[6] scanchain_59/module_data_in[7]
+ scanchain_59/module_data_out[0] scanchain_59/module_data_out[1] scanchain_59/module_data_out[2]
+ scanchain_59/module_data_out[3] scanchain_59/module_data_out[4] scanchain_59/module_data_out[5]
+ scanchain_59/module_data_out[6] scanchain_59/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_397 scanchain_397/clk_in scanchain_398/clk_in scanchain_397/data_in scanchain_398/data_in
+ scanchain_397/latch_enable_in scanchain_398/latch_enable_in scanchain_397/module_data_in[0]
+ scanchain_397/module_data_in[1] scanchain_397/module_data_in[2] scanchain_397/module_data_in[3]
+ scanchain_397/module_data_in[4] scanchain_397/module_data_in[5] scanchain_397/module_data_in[6]
+ scanchain_397/module_data_in[7] scanchain_397/module_data_out[0] scanchain_397/module_data_out[1]
+ scanchain_397/module_data_out[2] scanchain_397/module_data_out[3] scanchain_397/module_data_out[4]
+ scanchain_397/module_data_out[5] scanchain_397/module_data_out[6] scanchain_397/module_data_out[7]
+ scanchain_397/scan_select_in scanchain_398/scan_select_in vccd1 vssd1 scanchain
Xscanchain_386 scanchain_386/clk_in scanchain_387/clk_in scanchain_386/data_in scanchain_387/data_in
+ scanchain_386/latch_enable_in scanchain_387/latch_enable_in scanchain_386/module_data_in[0]
+ scanchain_386/module_data_in[1] scanchain_386/module_data_in[2] scanchain_386/module_data_in[3]
+ scanchain_386/module_data_in[4] scanchain_386/module_data_in[5] scanchain_386/module_data_in[6]
+ scanchain_386/module_data_in[7] scanchain_386/module_data_out[0] scanchain_386/module_data_out[1]
+ scanchain_386/module_data_out[2] scanchain_386/module_data_out[3] scanchain_386/module_data_out[4]
+ scanchain_386/module_data_out[5] scanchain_386/module_data_out[6] scanchain_386/module_data_out[7]
+ scanchain_386/scan_select_in scanchain_387/scan_select_in vccd1 vssd1 scanchain
Xscanchain_364 scanchain_364/clk_in scanchain_365/clk_in scanchain_364/data_in scanchain_365/data_in
+ scanchain_364/latch_enable_in scanchain_365/latch_enable_in scanchain_364/module_data_in[0]
+ scanchain_364/module_data_in[1] scanchain_364/module_data_in[2] scanchain_364/module_data_in[3]
+ scanchain_364/module_data_in[4] scanchain_364/module_data_in[5] scanchain_364/module_data_in[6]
+ scanchain_364/module_data_in[7] scanchain_364/module_data_out[0] scanchain_364/module_data_out[1]
+ scanchain_364/module_data_out[2] scanchain_364/module_data_out[3] scanchain_364/module_data_out[4]
+ scanchain_364/module_data_out[5] scanchain_364/module_data_out[6] scanchain_364/module_data_out[7]
+ scanchain_364/scan_select_in scanchain_365/scan_select_in vccd1 vssd1 scanchain
Xscanchain_375 scanchain_375/clk_in scanchain_376/clk_in scanchain_375/data_in scanchain_376/data_in
+ scanchain_375/latch_enable_in scanchain_376/latch_enable_in scanchain_375/module_data_in[0]
+ scanchain_375/module_data_in[1] scanchain_375/module_data_in[2] scanchain_375/module_data_in[3]
+ scanchain_375/module_data_in[4] scanchain_375/module_data_in[5] scanchain_375/module_data_in[6]
+ scanchain_375/module_data_in[7] scanchain_375/module_data_out[0] scanchain_375/module_data_out[1]
+ scanchain_375/module_data_out[2] scanchain_375/module_data_out[3] scanchain_375/module_data_out[4]
+ scanchain_375/module_data_out[5] scanchain_375/module_data_out[6] scanchain_375/module_data_out[7]
+ scanchain_375/scan_select_in scanchain_376/scan_select_in vccd1 vssd1 scanchain
Xscanchain_353 scanchain_353/clk_in scanchain_354/clk_in scanchain_353/data_in scanchain_354/data_in
+ scanchain_353/latch_enable_in scanchain_354/latch_enable_in scanchain_353/module_data_in[0]
+ scanchain_353/module_data_in[1] scanchain_353/module_data_in[2] scanchain_353/module_data_in[3]
+ scanchain_353/module_data_in[4] scanchain_353/module_data_in[5] scanchain_353/module_data_in[6]
+ scanchain_353/module_data_in[7] scanchain_353/module_data_out[0] scanchain_353/module_data_out[1]
+ scanchain_353/module_data_out[2] scanchain_353/module_data_out[3] scanchain_353/module_data_out[4]
+ scanchain_353/module_data_out[5] scanchain_353/module_data_out[6] scanchain_353/module_data_out[7]
+ scanchain_353/scan_select_in scanchain_354/scan_select_in vccd1 vssd1 scanchain
Xscanchain_342 scanchain_342/clk_in scanchain_343/clk_in scanchain_342/data_in scanchain_343/data_in
+ scanchain_342/latch_enable_in scanchain_343/latch_enable_in scanchain_342/module_data_in[0]
+ scanchain_342/module_data_in[1] scanchain_342/module_data_in[2] scanchain_342/module_data_in[3]
+ scanchain_342/module_data_in[4] scanchain_342/module_data_in[5] scanchain_342/module_data_in[6]
+ scanchain_342/module_data_in[7] scanchain_342/module_data_out[0] scanchain_342/module_data_out[1]
+ scanchain_342/module_data_out[2] scanchain_342/module_data_out[3] scanchain_342/module_data_out[4]
+ scanchain_342/module_data_out[5] scanchain_342/module_data_out[6] scanchain_342/module_data_out[7]
+ scanchain_342/scan_select_in scanchain_343/scan_select_in vccd1 vssd1 scanchain
Xscanchain_331 scanchain_331/clk_in scanchain_332/clk_in scanchain_331/data_in scanchain_332/data_in
+ scanchain_331/latch_enable_in scanchain_332/latch_enable_in scanchain_331/module_data_in[0]
+ scanchain_331/module_data_in[1] scanchain_331/module_data_in[2] scanchain_331/module_data_in[3]
+ scanchain_331/module_data_in[4] scanchain_331/module_data_in[5] scanchain_331/module_data_in[6]
+ scanchain_331/module_data_in[7] scanchain_331/module_data_out[0] scanchain_331/module_data_out[1]
+ scanchain_331/module_data_out[2] scanchain_331/module_data_out[3] scanchain_331/module_data_out[4]
+ scanchain_331/module_data_out[5] scanchain_331/module_data_out[6] scanchain_331/module_data_out[7]
+ scanchain_331/scan_select_in scanchain_332/scan_select_in vccd1 vssd1 scanchain
Xscanchain_320 scanchain_320/clk_in scanchain_321/clk_in scanchain_320/data_in scanchain_321/data_in
+ scanchain_320/latch_enable_in scanchain_321/latch_enable_in scanchain_320/module_data_in[0]
+ scanchain_320/module_data_in[1] scanchain_320/module_data_in[2] scanchain_320/module_data_in[3]
+ scanchain_320/module_data_in[4] scanchain_320/module_data_in[5] scanchain_320/module_data_in[6]
+ scanchain_320/module_data_in[7] scanchain_320/module_data_out[0] scanchain_320/module_data_out[1]
+ scanchain_320/module_data_out[2] scanchain_320/module_data_out[3] scanchain_320/module_data_out[4]
+ scanchain_320/module_data_out[5] scanchain_320/module_data_out[6] scanchain_320/module_data_out[7]
+ scanchain_320/scan_select_in scanchain_321/scan_select_in vccd1 vssd1 scanchain
Xscanchain_19 scanchain_19/clk_in scanchain_20/clk_in scanchain_19/data_in scanchain_20/data_in
+ scanchain_19/latch_enable_in scanchain_20/latch_enable_in scanchain_19/module_data_in[0]
+ scanchain_19/module_data_in[1] scanchain_19/module_data_in[2] scanchain_19/module_data_in[3]
+ scanchain_19/module_data_in[4] scanchain_19/module_data_in[5] scanchain_19/module_data_in[6]
+ scanchain_19/module_data_in[7] scanchain_19/module_data_out[0] scanchain_19/module_data_out[1]
+ scanchain_19/module_data_out[2] scanchain_19/module_data_out[3] scanchain_19/module_data_out[4]
+ scanchain_19/module_data_out[5] scanchain_19/module_data_out[6] scanchain_19/module_data_out[7]
+ scanchain_19/scan_select_in scanchain_20/scan_select_in vccd1 vssd1 scanchain
Xscanchain_150 scanchain_150/clk_in scanchain_151/clk_in scanchain_150/data_in scanchain_151/data_in
+ scanchain_150/latch_enable_in scanchain_151/latch_enable_in scanchain_150/module_data_in[0]
+ scanchain_150/module_data_in[1] scanchain_150/module_data_in[2] scanchain_150/module_data_in[3]
+ scanchain_150/module_data_in[4] scanchain_150/module_data_in[5] scanchain_150/module_data_in[6]
+ scanchain_150/module_data_in[7] scanchain_150/module_data_out[0] scanchain_150/module_data_out[1]
+ scanchain_150/module_data_out[2] scanchain_150/module_data_out[3] scanchain_150/module_data_out[4]
+ scanchain_150/module_data_out[5] scanchain_150/module_data_out[6] scanchain_150/module_data_out[7]
+ scanchain_150/scan_select_in scanchain_151/scan_select_in vccd1 vssd1 scanchain
Xscanchain_161 scanchain_161/clk_in scanchain_162/clk_in scanchain_161/data_in scanchain_162/data_in
+ scanchain_161/latch_enable_in scanchain_162/latch_enable_in scanchain_161/module_data_in[0]
+ scanchain_161/module_data_in[1] scanchain_161/module_data_in[2] scanchain_161/module_data_in[3]
+ scanchain_161/module_data_in[4] scanchain_161/module_data_in[5] scanchain_161/module_data_in[6]
+ scanchain_161/module_data_in[7] scanchain_161/module_data_out[0] scanchain_161/module_data_out[1]
+ scanchain_161/module_data_out[2] scanchain_161/module_data_out[3] scanchain_161/module_data_out[4]
+ scanchain_161/module_data_out[5] scanchain_161/module_data_out[6] scanchain_161/module_data_out[7]
+ scanchain_161/scan_select_in scanchain_162/scan_select_in vccd1 vssd1 scanchain
Xscanchain_194 scanchain_194/clk_in scanchain_195/clk_in scanchain_194/data_in scanchain_195/data_in
+ scanchain_194/latch_enable_in scanchain_195/latch_enable_in scanchain_194/module_data_in[0]
+ scanchain_194/module_data_in[1] scanchain_194/module_data_in[2] scanchain_194/module_data_in[3]
+ scanchain_194/module_data_in[4] scanchain_194/module_data_in[5] scanchain_194/module_data_in[6]
+ scanchain_194/module_data_in[7] scanchain_194/module_data_out[0] scanchain_194/module_data_out[1]
+ scanchain_194/module_data_out[2] scanchain_194/module_data_out[3] scanchain_194/module_data_out[4]
+ scanchain_194/module_data_out[5] scanchain_194/module_data_out[6] scanchain_194/module_data_out[7]
+ scanchain_194/scan_select_in scanchain_195/scan_select_in vccd1 vssd1 scanchain
Xscanchain_183 scanchain_183/clk_in scanchain_184/clk_in scanchain_183/data_in scanchain_184/data_in
+ scanchain_183/latch_enable_in scanchain_184/latch_enable_in scanchain_183/module_data_in[0]
+ scanchain_183/module_data_in[1] scanchain_183/module_data_in[2] scanchain_183/module_data_in[3]
+ scanchain_183/module_data_in[4] scanchain_183/module_data_in[5] scanchain_183/module_data_in[6]
+ scanchain_183/module_data_in[7] scanchain_183/module_data_out[0] scanchain_183/module_data_out[1]
+ scanchain_183/module_data_out[2] scanchain_183/module_data_out[3] scanchain_183/module_data_out[4]
+ scanchain_183/module_data_out[5] scanchain_183/module_data_out[6] scanchain_183/module_data_out[7]
+ scanchain_183/scan_select_in scanchain_184/scan_select_in vccd1 vssd1 scanchain
Xscanchain_172 scanchain_172/clk_in scanchain_173/clk_in scanchain_172/data_in scanchain_173/data_in
+ scanchain_172/latch_enable_in scanchain_173/latch_enable_in scanchain_172/module_data_in[0]
+ scanchain_172/module_data_in[1] scanchain_172/module_data_in[2] scanchain_172/module_data_in[3]
+ scanchain_172/module_data_in[4] scanchain_172/module_data_in[5] scanchain_172/module_data_in[6]
+ scanchain_172/module_data_in[7] scanchain_172/module_data_out[0] scanchain_172/module_data_out[1]
+ scanchain_172/module_data_out[2] scanchain_172/module_data_out[3] scanchain_172/module_data_out[4]
+ scanchain_172/module_data_out[5] scanchain_172/module_data_out[6] scanchain_172/module_data_out[7]
+ scanchain_172/scan_select_in scanchain_173/scan_select_in vccd1 vssd1 scanchain
Xalu_top_7 alu_top_7/io_in[0] alu_top_7/io_in[1] alu_top_7/io_in[2] alu_top_7/io_in[3]
+ alu_top_7/io_in[4] alu_top_7/io_in[5] alu_top_7/io_in[6] alu_top_7/io_in[7] alu_top_7/io_out[0]
+ alu_top_7/io_out[1] alu_top_7/io_out[2] alu_top_7/io_out[3] alu_top_7/io_out[4]
+ alu_top_7/io_out[5] alu_top_7/io_out[6] alu_top_7/io_out[7] vccd1 vssd1 alu_top
Xmigcorre_pwm_5 migcorre_pwm_5/io_in[0] migcorre_pwm_5/io_in[1] migcorre_pwm_5/io_in[2]
+ migcorre_pwm_5/io_in[3] migcorre_pwm_5/io_in[4] migcorre_pwm_5/io_in[5] migcorre_pwm_5/io_in[6]
+ migcorre_pwm_5/io_in[7] migcorre_pwm_5/io_out[0] migcorre_pwm_5/io_out[1] migcorre_pwm_5/io_out[2]
+ migcorre_pwm_5/io_out[3] migcorre_pwm_5/io_out[4] migcorre_pwm_5/io_out[5] migcorre_pwm_5/io_out[6]
+ migcorre_pwm_5/io_out[7] vccd1 vssd1 migcorre_pwm
Xuser_module_339501025136214612_229 scanchain_229/module_data_in[0] scanchain_229/module_data_in[1]
+ scanchain_229/module_data_in[2] scanchain_229/module_data_in[3] scanchain_229/module_data_in[4]
+ scanchain_229/module_data_in[5] scanchain_229/module_data_in[6] scanchain_229/module_data_in[7]
+ scanchain_229/module_data_out[0] scanchain_229/module_data_out[1] scanchain_229/module_data_out[2]
+ scanchain_229/module_data_out[3] scanchain_229/module_data_out[4] scanchain_229/module_data_out[5]
+ scanchain_229/module_data_out[6] scanchain_229/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_207 scanchain_207/module_data_in[0] scanchain_207/module_data_in[1]
+ scanchain_207/module_data_in[2] scanchain_207/module_data_in[3] scanchain_207/module_data_in[4]
+ scanchain_207/module_data_in[5] scanchain_207/module_data_in[6] scanchain_207/module_data_in[7]
+ scanchain_207/module_data_out[0] scanchain_207/module_data_out[1] scanchain_207/module_data_out[2]
+ scanchain_207/module_data_out[3] scanchain_207/module_data_out[4] scanchain_207/module_data_out[5]
+ scanchain_207/module_data_out[6] scanchain_207/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_218 scanchain_218/module_data_in[0] scanchain_218/module_data_in[1]
+ scanchain_218/module_data_in[2] scanchain_218/module_data_in[3] scanchain_218/module_data_in[4]
+ scanchain_218/module_data_in[5] scanchain_218/module_data_in[6] scanchain_218/module_data_in[7]
+ scanchain_218/module_data_out[0] scanchain_218/module_data_out[1] scanchain_218/module_data_out[2]
+ scanchain_218/module_data_out[3] scanchain_218/module_data_out[4] scanchain_218/module_data_out[5]
+ scanchain_218/module_data_out[6] scanchain_218/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_398 scanchain_398/clk_in scanchain_399/clk_in scanchain_398/data_in scanchain_399/data_in
+ scanchain_398/latch_enable_in scanchain_399/latch_enable_in scanchain_398/module_data_in[0]
+ scanchain_398/module_data_in[1] scanchain_398/module_data_in[2] scanchain_398/module_data_in[3]
+ scanchain_398/module_data_in[4] scanchain_398/module_data_in[5] scanchain_398/module_data_in[6]
+ scanchain_398/module_data_in[7] scanchain_398/module_data_out[0] scanchain_398/module_data_out[1]
+ scanchain_398/module_data_out[2] scanchain_398/module_data_out[3] scanchain_398/module_data_out[4]
+ scanchain_398/module_data_out[5] scanchain_398/module_data_out[6] scanchain_398/module_data_out[7]
+ scanchain_398/scan_select_in scanchain_399/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_390 scanchain_390/module_data_in[0] scanchain_390/module_data_in[1]
+ scanchain_390/module_data_in[2] scanchain_390/module_data_in[3] scanchain_390/module_data_in[4]
+ scanchain_390/module_data_in[5] scanchain_390/module_data_in[6] scanchain_390/module_data_in[7]
+ scanchain_390/module_data_out[0] scanchain_390/module_data_out[1] scanchain_390/module_data_out[2]
+ scanchain_390/module_data_out[3] scanchain_390/module_data_out[4] scanchain_390/module_data_out[5]
+ scanchain_390/module_data_out[6] scanchain_390/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_387 scanchain_387/clk_in scanchain_388/clk_in scanchain_387/data_in scanchain_388/data_in
+ scanchain_387/latch_enable_in scanchain_388/latch_enable_in scanchain_387/module_data_in[0]
+ scanchain_387/module_data_in[1] scanchain_387/module_data_in[2] scanchain_387/module_data_in[3]
+ scanchain_387/module_data_in[4] scanchain_387/module_data_in[5] scanchain_387/module_data_in[6]
+ scanchain_387/module_data_in[7] scanchain_387/module_data_out[0] scanchain_387/module_data_out[1]
+ scanchain_387/module_data_out[2] scanchain_387/module_data_out[3] scanchain_387/module_data_out[4]
+ scanchain_387/module_data_out[5] scanchain_387/module_data_out[6] scanchain_387/module_data_out[7]
+ scanchain_387/scan_select_in scanchain_388/scan_select_in vccd1 vssd1 scanchain
Xscanchain_365 scanchain_365/clk_in scanchain_366/clk_in scanchain_365/data_in scanchain_366/data_in
+ scanchain_365/latch_enable_in scanchain_366/latch_enable_in scanchain_365/module_data_in[0]
+ scanchain_365/module_data_in[1] scanchain_365/module_data_in[2] scanchain_365/module_data_in[3]
+ scanchain_365/module_data_in[4] scanchain_365/module_data_in[5] scanchain_365/module_data_in[6]
+ scanchain_365/module_data_in[7] scanchain_365/module_data_out[0] scanchain_365/module_data_out[1]
+ scanchain_365/module_data_out[2] scanchain_365/module_data_out[3] scanchain_365/module_data_out[4]
+ scanchain_365/module_data_out[5] scanchain_365/module_data_out[6] scanchain_365/module_data_out[7]
+ scanchain_365/scan_select_in scanchain_366/scan_select_in vccd1 vssd1 scanchain
Xscanchain_376 scanchain_376/clk_in scanchain_377/clk_in scanchain_376/data_in scanchain_377/data_in
+ scanchain_376/latch_enable_in scanchain_377/latch_enable_in scanchain_376/module_data_in[0]
+ scanchain_376/module_data_in[1] scanchain_376/module_data_in[2] scanchain_376/module_data_in[3]
+ scanchain_376/module_data_in[4] scanchain_376/module_data_in[5] scanchain_376/module_data_in[6]
+ scanchain_376/module_data_in[7] scanchain_376/module_data_out[0] scanchain_376/module_data_out[1]
+ scanchain_376/module_data_out[2] scanchain_376/module_data_out[3] scanchain_376/module_data_out[4]
+ scanchain_376/module_data_out[5] scanchain_376/module_data_out[6] scanchain_376/module_data_out[7]
+ scanchain_376/scan_select_in scanchain_377/scan_select_in vccd1 vssd1 scanchain
Xscanchain_354 scanchain_354/clk_in scanchain_355/clk_in scanchain_354/data_in scanchain_355/data_in
+ scanchain_354/latch_enable_in scanchain_355/latch_enable_in scanchain_354/module_data_in[0]
+ scanchain_354/module_data_in[1] scanchain_354/module_data_in[2] scanchain_354/module_data_in[3]
+ scanchain_354/module_data_in[4] scanchain_354/module_data_in[5] scanchain_354/module_data_in[6]
+ scanchain_354/module_data_in[7] scanchain_354/module_data_out[0] scanchain_354/module_data_out[1]
+ scanchain_354/module_data_out[2] scanchain_354/module_data_out[3] scanchain_354/module_data_out[4]
+ scanchain_354/module_data_out[5] scanchain_354/module_data_out[6] scanchain_354/module_data_out[7]
+ scanchain_354/scan_select_in scanchain_355/scan_select_in vccd1 vssd1 scanchain
Xscanchain_343 scanchain_343/clk_in scanchain_344/clk_in scanchain_343/data_in scanchain_344/data_in
+ scanchain_343/latch_enable_in scanchain_344/latch_enable_in scanchain_343/module_data_in[0]
+ scanchain_343/module_data_in[1] scanchain_343/module_data_in[2] scanchain_343/module_data_in[3]
+ scanchain_343/module_data_in[4] scanchain_343/module_data_in[5] scanchain_343/module_data_in[6]
+ scanchain_343/module_data_in[7] scanchain_343/module_data_out[0] scanchain_343/module_data_out[1]
+ scanchain_343/module_data_out[2] scanchain_343/module_data_out[3] scanchain_343/module_data_out[4]
+ scanchain_343/module_data_out[5] scanchain_343/module_data_out[6] scanchain_343/module_data_out[7]
+ scanchain_343/scan_select_in scanchain_344/scan_select_in vccd1 vssd1 scanchain
Xscanchain_321 scanchain_321/clk_in scanchain_322/clk_in scanchain_321/data_in scanchain_322/data_in
+ scanchain_321/latch_enable_in scanchain_322/latch_enable_in scanchain_321/module_data_in[0]
+ scanchain_321/module_data_in[1] scanchain_321/module_data_in[2] scanchain_321/module_data_in[3]
+ scanchain_321/module_data_in[4] scanchain_321/module_data_in[5] scanchain_321/module_data_in[6]
+ scanchain_321/module_data_in[7] scanchain_321/module_data_out[0] scanchain_321/module_data_out[1]
+ scanchain_321/module_data_out[2] scanchain_321/module_data_out[3] scanchain_321/module_data_out[4]
+ scanchain_321/module_data_out[5] scanchain_321/module_data_out[6] scanchain_321/module_data_out[7]
+ scanchain_321/scan_select_in scanchain_322/scan_select_in vccd1 vssd1 scanchain
Xscanchain_332 scanchain_332/clk_in scanchain_333/clk_in scanchain_332/data_in scanchain_333/data_in
+ scanchain_332/latch_enable_in scanchain_333/latch_enable_in scanchain_332/module_data_in[0]
+ scanchain_332/module_data_in[1] scanchain_332/module_data_in[2] scanchain_332/module_data_in[3]
+ scanchain_332/module_data_in[4] scanchain_332/module_data_in[5] scanchain_332/module_data_in[6]
+ scanchain_332/module_data_in[7] scanchain_332/module_data_out[0] scanchain_332/module_data_out[1]
+ scanchain_332/module_data_out[2] scanchain_332/module_data_out[3] scanchain_332/module_data_out[4]
+ scanchain_332/module_data_out[5] scanchain_332/module_data_out[6] scanchain_332/module_data_out[7]
+ scanchain_332/scan_select_in scanchain_333/scan_select_in vccd1 vssd1 scanchain
Xscanchain_310 scanchain_310/clk_in scanchain_311/clk_in scanchain_310/data_in scanchain_311/data_in
+ scanchain_310/latch_enable_in scanchain_311/latch_enable_in scanchain_310/module_data_in[0]
+ scanchain_310/module_data_in[1] scanchain_310/module_data_in[2] scanchain_310/module_data_in[3]
+ scanchain_310/module_data_in[4] scanchain_310/module_data_in[5] scanchain_310/module_data_in[6]
+ scanchain_310/module_data_in[7] scanchain_310/module_data_out[0] scanchain_310/module_data_out[1]
+ scanchain_310/module_data_out[2] scanchain_310/module_data_out[3] scanchain_310/module_data_out[4]
+ scanchain_310/module_data_out[5] scanchain_310/module_data_out[6] scanchain_310/module_data_out[7]
+ scanchain_310/scan_select_in scanchain_311/scan_select_in vccd1 vssd1 scanchain
Xscanchain_195 scanchain_195/clk_in scanchain_196/clk_in scanchain_195/data_in scanchain_196/data_in
+ scanchain_195/latch_enable_in scanchain_196/latch_enable_in scanchain_195/module_data_in[0]
+ scanchain_195/module_data_in[1] scanchain_195/module_data_in[2] scanchain_195/module_data_in[3]
+ scanchain_195/module_data_in[4] scanchain_195/module_data_in[5] scanchain_195/module_data_in[6]
+ scanchain_195/module_data_in[7] scanchain_195/module_data_out[0] scanchain_195/module_data_out[1]
+ scanchain_195/module_data_out[2] scanchain_195/module_data_out[3] scanchain_195/module_data_out[4]
+ scanchain_195/module_data_out[5] scanchain_195/module_data_out[6] scanchain_195/module_data_out[7]
+ scanchain_195/scan_select_in scanchain_196/scan_select_in vccd1 vssd1 scanchain
Xuser_module_347894637149553236_17 scanchain_17/module_data_in[0] scanchain_17/module_data_in[1]
+ scanchain_17/module_data_in[2] scanchain_17/module_data_in[3] scanchain_17/module_data_in[4]
+ scanchain_17/module_data_in[5] scanchain_17/module_data_in[6] scanchain_17/module_data_in[7]
+ scanchain_17/module_data_out[0] scanchain_17/module_data_out[1] scanchain_17/module_data_out[2]
+ scanchain_17/module_data_out[3] scanchain_17/module_data_out[4] scanchain_17/module_data_out[5]
+ scanchain_17/module_data_out[6] scanchain_17/module_data_out[7] vccd1 vssd1 user_module_347894637149553236
Xscanchain_140 scanchain_140/clk_in scanchain_141/clk_in scanchain_140/data_in scanchain_141/data_in
+ scanchain_140/latch_enable_in scanchain_141/latch_enable_in scanchain_140/module_data_in[0]
+ scanchain_140/module_data_in[1] scanchain_140/module_data_in[2] scanchain_140/module_data_in[3]
+ scanchain_140/module_data_in[4] scanchain_140/module_data_in[5] scanchain_140/module_data_in[6]
+ scanchain_140/module_data_in[7] scanchain_140/module_data_out[0] scanchain_140/module_data_out[1]
+ scanchain_140/module_data_out[2] scanchain_140/module_data_out[3] scanchain_140/module_data_out[4]
+ scanchain_140/module_data_out[5] scanchain_140/module_data_out[6] scanchain_140/module_data_out[7]
+ scanchain_140/scan_select_in scanchain_141/scan_select_in vccd1 vssd1 scanchain
Xscanchain_151 scanchain_151/clk_in scanchain_152/clk_in scanchain_151/data_in scanchain_152/data_in
+ scanchain_151/latch_enable_in scanchain_152/latch_enable_in scanchain_151/module_data_in[0]
+ scanchain_151/module_data_in[1] scanchain_151/module_data_in[2] scanchain_151/module_data_in[3]
+ scanchain_151/module_data_in[4] scanchain_151/module_data_in[5] scanchain_151/module_data_in[6]
+ scanchain_151/module_data_in[7] scanchain_151/module_data_out[0] scanchain_151/module_data_out[1]
+ scanchain_151/module_data_out[2] scanchain_151/module_data_out[3] scanchain_151/module_data_out[4]
+ scanchain_151/module_data_out[5] scanchain_151/module_data_out[6] scanchain_151/module_data_out[7]
+ scanchain_151/scan_select_in scanchain_152/scan_select_in vccd1 vssd1 scanchain
Xscanchain_162 scanchain_162/clk_in scanchain_163/clk_in scanchain_162/data_in scanchain_163/data_in
+ scanchain_162/latch_enable_in scanchain_163/latch_enable_in scanchain_162/module_data_in[0]
+ scanchain_162/module_data_in[1] scanchain_162/module_data_in[2] scanchain_162/module_data_in[3]
+ scanchain_162/module_data_in[4] scanchain_162/module_data_in[5] scanchain_162/module_data_in[6]
+ scanchain_162/module_data_in[7] scanchain_162/module_data_out[0] scanchain_162/module_data_out[1]
+ scanchain_162/module_data_out[2] scanchain_162/module_data_out[3] scanchain_162/module_data_out[4]
+ scanchain_162/module_data_out[5] scanchain_162/module_data_out[6] scanchain_162/module_data_out[7]
+ scanchain_162/scan_select_in scanchain_163/scan_select_in vccd1 vssd1 scanchain
Xscanchain_184 scanchain_184/clk_in scanchain_185/clk_in scanchain_184/data_in scanchain_185/data_in
+ scanchain_184/latch_enable_in scanchain_185/latch_enable_in scanchain_184/module_data_in[0]
+ scanchain_184/module_data_in[1] scanchain_184/module_data_in[2] scanchain_184/module_data_in[3]
+ scanchain_184/module_data_in[4] scanchain_184/module_data_in[5] scanchain_184/module_data_in[6]
+ scanchain_184/module_data_in[7] scanchain_184/module_data_out[0] scanchain_184/module_data_out[1]
+ scanchain_184/module_data_out[2] scanchain_184/module_data_out[3] scanchain_184/module_data_out[4]
+ scanchain_184/module_data_out[5] scanchain_184/module_data_out[6] scanchain_184/module_data_out[7]
+ scanchain_184/scan_select_in scanchain_185/scan_select_in vccd1 vssd1 scanchain
Xscanchain_173 scanchain_173/clk_in scanchain_174/clk_in scanchain_173/data_in scanchain_174/data_in
+ scanchain_173/latch_enable_in scanchain_174/latch_enable_in scanchain_173/module_data_in[0]
+ scanchain_173/module_data_in[1] scanchain_173/module_data_in[2] scanchain_173/module_data_in[3]
+ scanchain_173/module_data_in[4] scanchain_173/module_data_in[5] scanchain_173/module_data_in[6]
+ scanchain_173/module_data_in[7] scanchain_173/module_data_out[0] scanchain_173/module_data_out[1]
+ scanchain_173/module_data_out[2] scanchain_173/module_data_out[3] scanchain_173/module_data_out[4]
+ scanchain_173/module_data_out[5] scanchain_173/module_data_out[6] scanchain_173/module_data_out[7]
+ scanchain_173/scan_select_in scanchain_174/scan_select_in vccd1 vssd1 scanchain
Xazdle_binary_clock_9 scanchain_9/module_data_in[0] scanchain_9/module_data_in[1]
+ scanchain_9/module_data_in[2] scanchain_9/module_data_in[3] scanchain_9/module_data_in[4]
+ scanchain_9/module_data_in[5] scanchain_9/module_data_in[6] scanchain_9/module_data_in[7]
+ scanchain_9/module_data_out[0] scanchain_9/module_data_out[1] scanchain_9/module_data_out[2]
+ scanchain_9/module_data_out[3] scanchain_9/module_data_out[4] scanchain_9/module_data_out[5]
+ scanchain_9/module_data_out[6] scanchain_9/module_data_out[7] vccd1 vssd1 azdle_binary_clock
Xuser_module_339501025136214612_208 scanchain_208/module_data_in[0] scanchain_208/module_data_in[1]
+ scanchain_208/module_data_in[2] scanchain_208/module_data_in[3] scanchain_208/module_data_in[4]
+ scanchain_208/module_data_in[5] scanchain_208/module_data_in[6] scanchain_208/module_data_in[7]
+ scanchain_208/module_data_out[0] scanchain_208/module_data_out[1] scanchain_208/module_data_out[2]
+ scanchain_208/module_data_out[3] scanchain_208/module_data_out[4] scanchain_208/module_data_out[5]
+ scanchain_208/module_data_out[6] scanchain_208/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_219 scanchain_219/module_data_in[0] scanchain_219/module_data_in[1]
+ scanchain_219/module_data_in[2] scanchain_219/module_data_in[3] scanchain_219/module_data_in[4]
+ scanchain_219/module_data_in[5] scanchain_219/module_data_in[6] scanchain_219/module_data_in[7]
+ scanchain_219/module_data_out[0] scanchain_219/module_data_out[1] scanchain_219/module_data_out[2]
+ scanchain_219/module_data_out[3] scanchain_219/module_data_out[4] scanchain_219/module_data_out[5]
+ scanchain_219/module_data_out[6] scanchain_219/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xphasenoisepon_seven_segment_seconds_46 scanchain_46/module_data_in[0] scanchain_46/module_data_in[1]
+ scanchain_46/module_data_in[2] scanchain_46/module_data_in[3] scanchain_46/module_data_in[4]
+ scanchain_46/module_data_in[5] scanchain_46/module_data_in[6] scanchain_46/module_data_in[7]
+ scanchain_46/module_data_out[0] scanchain_46/module_data_out[1] scanchain_46/module_data_out[2]
+ scanchain_46/module_data_out[3] scanchain_46/module_data_out[4] scanchain_46/module_data_out[5]
+ scanchain_46/module_data_out[6] scanchain_46/module_data_out[7] vccd1 vssd1 phasenoisepon_seven_segment_seconds
Xjar_sram_top_11 jar_sram_top_11/io_in[0] jar_sram_top_11/io_in[1] jar_sram_top_11/io_in[2]
+ jar_sram_top_11/io_in[3] jar_sram_top_11/io_in[4] jar_sram_top_11/io_in[5] jar_sram_top_11/io_in[6]
+ jar_sram_top_11/io_in[7] jar_sram_top_11/io_out[0] jar_sram_top_11/io_out[1] jar_sram_top_11/io_out[2]
+ jar_sram_top_11/io_out[3] jar_sram_top_11/io_out[4] jar_sram_top_11/io_out[5] jar_sram_top_11/io_out[6]
+ jar_sram_top_11/io_out[7] vccd1 vssd1 jar_sram_top
Xuser_module_341620484740219475_41 scanchain_41/module_data_in[0] scanchain_41/module_data_in[1]
+ scanchain_41/module_data_in[2] scanchain_41/module_data_in[3] scanchain_41/module_data_in[4]
+ scanchain_41/module_data_in[5] scanchain_41/module_data_in[6] scanchain_41/module_data_in[7]
+ scanchain_41/module_data_out[0] scanchain_41/module_data_out[1] scanchain_41/module_data_out[2]
+ scanchain_41/module_data_out[3] scanchain_41/module_data_out[4] scanchain_41/module_data_out[5]
+ scanchain_41/module_data_out[6] scanchain_41/module_data_out[7] vccd1 vssd1 user_module_341620484740219475
Xscanchain_399 scanchain_399/clk_in scanchain_400/clk_in scanchain_399/data_in scanchain_400/data_in
+ scanchain_399/latch_enable_in scanchain_400/latch_enable_in scanchain_399/module_data_in[0]
+ scanchain_399/module_data_in[1] scanchain_399/module_data_in[2] scanchain_399/module_data_in[3]
+ scanchain_399/module_data_in[4] scanchain_399/module_data_in[5] scanchain_399/module_data_in[6]
+ scanchain_399/module_data_in[7] scanchain_399/module_data_out[0] scanchain_399/module_data_out[1]
+ scanchain_399/module_data_out[2] scanchain_399/module_data_out[3] scanchain_399/module_data_out[4]
+ scanchain_399/module_data_out[5] scanchain_399/module_data_out[6] scanchain_399/module_data_out[7]
+ scanchain_399/scan_select_in scanchain_400/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_391 scanchain_391/module_data_in[0] scanchain_391/module_data_in[1]
+ scanchain_391/module_data_in[2] scanchain_391/module_data_in[3] scanchain_391/module_data_in[4]
+ scanchain_391/module_data_in[5] scanchain_391/module_data_in[6] scanchain_391/module_data_in[7]
+ scanchain_391/module_data_out[0] scanchain_391/module_data_out[1] scanchain_391/module_data_out[2]
+ scanchain_391/module_data_out[3] scanchain_391/module_data_out[4] scanchain_391/module_data_out[5]
+ scanchain_391/module_data_out[6] scanchain_391/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_388 scanchain_388/clk_in scanchain_389/clk_in scanchain_388/data_in scanchain_389/data_in
+ scanchain_388/latch_enable_in scanchain_389/latch_enable_in scanchain_388/module_data_in[0]
+ scanchain_388/module_data_in[1] scanchain_388/module_data_in[2] scanchain_388/module_data_in[3]
+ scanchain_388/module_data_in[4] scanchain_388/module_data_in[5] scanchain_388/module_data_in[6]
+ scanchain_388/module_data_in[7] scanchain_388/module_data_out[0] scanchain_388/module_data_out[1]
+ scanchain_388/module_data_out[2] scanchain_388/module_data_out[3] scanchain_388/module_data_out[4]
+ scanchain_388/module_data_out[5] scanchain_388/module_data_out[6] scanchain_388/module_data_out[7]
+ scanchain_388/scan_select_in scanchain_389/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_380 scanchain_380/module_data_in[0] scanchain_380/module_data_in[1]
+ scanchain_380/module_data_in[2] scanchain_380/module_data_in[3] scanchain_380/module_data_in[4]
+ scanchain_380/module_data_in[5] scanchain_380/module_data_in[6] scanchain_380/module_data_in[7]
+ scanchain_380/module_data_out[0] scanchain_380/module_data_out[1] scanchain_380/module_data_out[2]
+ scanchain_380/module_data_out[3] scanchain_380/module_data_out[4] scanchain_380/module_data_out[5]
+ scanchain_380/module_data_out[6] scanchain_380/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_366 scanchain_366/clk_in scanchain_367/clk_in scanchain_366/data_in scanchain_367/data_in
+ scanchain_366/latch_enable_in scanchain_367/latch_enable_in scanchain_366/module_data_in[0]
+ scanchain_366/module_data_in[1] scanchain_366/module_data_in[2] scanchain_366/module_data_in[3]
+ scanchain_366/module_data_in[4] scanchain_366/module_data_in[5] scanchain_366/module_data_in[6]
+ scanchain_366/module_data_in[7] scanchain_366/module_data_out[0] scanchain_366/module_data_out[1]
+ scanchain_366/module_data_out[2] scanchain_366/module_data_out[3] scanchain_366/module_data_out[4]
+ scanchain_366/module_data_out[5] scanchain_366/module_data_out[6] scanchain_366/module_data_out[7]
+ scanchain_366/scan_select_in scanchain_367/scan_select_in vccd1 vssd1 scanchain
Xscanchain_377 scanchain_377/clk_in scanchain_378/clk_in scanchain_377/data_in scanchain_378/data_in
+ scanchain_377/latch_enable_in scanchain_378/latch_enable_in scanchain_377/module_data_in[0]
+ scanchain_377/module_data_in[1] scanchain_377/module_data_in[2] scanchain_377/module_data_in[3]
+ scanchain_377/module_data_in[4] scanchain_377/module_data_in[5] scanchain_377/module_data_in[6]
+ scanchain_377/module_data_in[7] scanchain_377/module_data_out[0] scanchain_377/module_data_out[1]
+ scanchain_377/module_data_out[2] scanchain_377/module_data_out[3] scanchain_377/module_data_out[4]
+ scanchain_377/module_data_out[5] scanchain_377/module_data_out[6] scanchain_377/module_data_out[7]
+ scanchain_377/scan_select_in scanchain_378/scan_select_in vccd1 vssd1 scanchain
Xscanchain_355 scanchain_355/clk_in scanchain_356/clk_in scanchain_355/data_in scanchain_356/data_in
+ scanchain_355/latch_enable_in scanchain_356/latch_enable_in scanchain_355/module_data_in[0]
+ scanchain_355/module_data_in[1] scanchain_355/module_data_in[2] scanchain_355/module_data_in[3]
+ scanchain_355/module_data_in[4] scanchain_355/module_data_in[5] scanchain_355/module_data_in[6]
+ scanchain_355/module_data_in[7] scanchain_355/module_data_out[0] scanchain_355/module_data_out[1]
+ scanchain_355/module_data_out[2] scanchain_355/module_data_out[3] scanchain_355/module_data_out[4]
+ scanchain_355/module_data_out[5] scanchain_355/module_data_out[6] scanchain_355/module_data_out[7]
+ scanchain_355/scan_select_in scanchain_356/scan_select_in vccd1 vssd1 scanchain
Xscanchain_344 scanchain_344/clk_in scanchain_345/clk_in scanchain_344/data_in scanchain_345/data_in
+ scanchain_344/latch_enable_in scanchain_345/latch_enable_in scanchain_344/module_data_in[0]
+ scanchain_344/module_data_in[1] scanchain_344/module_data_in[2] scanchain_344/module_data_in[3]
+ scanchain_344/module_data_in[4] scanchain_344/module_data_in[5] scanchain_344/module_data_in[6]
+ scanchain_344/module_data_in[7] scanchain_344/module_data_out[0] scanchain_344/module_data_out[1]
+ scanchain_344/module_data_out[2] scanchain_344/module_data_out[3] scanchain_344/module_data_out[4]
+ scanchain_344/module_data_out[5] scanchain_344/module_data_out[6] scanchain_344/module_data_out[7]
+ scanchain_344/scan_select_in scanchain_345/scan_select_in vccd1 vssd1 scanchain
Xscanchain_322 scanchain_322/clk_in scanchain_323/clk_in scanchain_322/data_in scanchain_323/data_in
+ scanchain_322/latch_enable_in scanchain_323/latch_enable_in scanchain_322/module_data_in[0]
+ scanchain_322/module_data_in[1] scanchain_322/module_data_in[2] scanchain_322/module_data_in[3]
+ scanchain_322/module_data_in[4] scanchain_322/module_data_in[5] scanchain_322/module_data_in[6]
+ scanchain_322/module_data_in[7] scanchain_322/module_data_out[0] scanchain_322/module_data_out[1]
+ scanchain_322/module_data_out[2] scanchain_322/module_data_out[3] scanchain_322/module_data_out[4]
+ scanchain_322/module_data_out[5] scanchain_322/module_data_out[6] scanchain_322/module_data_out[7]
+ scanchain_322/scan_select_in scanchain_323/scan_select_in vccd1 vssd1 scanchain
Xscanchain_333 scanchain_333/clk_in scanchain_334/clk_in scanchain_333/data_in scanchain_334/data_in
+ scanchain_333/latch_enable_in scanchain_334/latch_enable_in scanchain_333/module_data_in[0]
+ scanchain_333/module_data_in[1] scanchain_333/module_data_in[2] scanchain_333/module_data_in[3]
+ scanchain_333/module_data_in[4] scanchain_333/module_data_in[5] scanchain_333/module_data_in[6]
+ scanchain_333/module_data_in[7] scanchain_333/module_data_out[0] scanchain_333/module_data_out[1]
+ scanchain_333/module_data_out[2] scanchain_333/module_data_out[3] scanchain_333/module_data_out[4]
+ scanchain_333/module_data_out[5] scanchain_333/module_data_out[6] scanchain_333/module_data_out[7]
+ scanchain_333/scan_select_in scanchain_334/scan_select_in vccd1 vssd1 scanchain
Xscanchain_311 scanchain_311/clk_in scanchain_312/clk_in scanchain_311/data_in scanchain_312/data_in
+ scanchain_311/latch_enable_in scanchain_312/latch_enable_in scanchain_311/module_data_in[0]
+ scanchain_311/module_data_in[1] scanchain_311/module_data_in[2] scanchain_311/module_data_in[3]
+ scanchain_311/module_data_in[4] scanchain_311/module_data_in[5] scanchain_311/module_data_in[6]
+ scanchain_311/module_data_in[7] scanchain_311/module_data_out[0] scanchain_311/module_data_out[1]
+ scanchain_311/module_data_out[2] scanchain_311/module_data_out[3] scanchain_311/module_data_out[4]
+ scanchain_311/module_data_out[5] scanchain_311/module_data_out[6] scanchain_311/module_data_out[7]
+ scanchain_311/scan_select_in scanchain_312/scan_select_in vccd1 vssd1 scanchain
Xscanchain_300 scanchain_300/clk_in scanchain_301/clk_in scanchain_300/data_in scanchain_301/data_in
+ scanchain_300/latch_enable_in scanchain_301/latch_enable_in scanchain_300/module_data_in[0]
+ scanchain_300/module_data_in[1] scanchain_300/module_data_in[2] scanchain_300/module_data_in[3]
+ scanchain_300/module_data_in[4] scanchain_300/module_data_in[5] scanchain_300/module_data_in[6]
+ scanchain_300/module_data_in[7] scanchain_300/module_data_out[0] scanchain_300/module_data_out[1]
+ scanchain_300/module_data_out[2] scanchain_300/module_data_out[3] scanchain_300/module_data_out[4]
+ scanchain_300/module_data_out[5] scanchain_300/module_data_out[6] scanchain_300/module_data_out[7]
+ scanchain_300/scan_select_in scanchain_301/scan_select_in vccd1 vssd1 scanchain
Xscanchain_196 scanchain_196/clk_in scanchain_197/clk_in scanchain_196/data_in scanchain_197/data_in
+ scanchain_196/latch_enable_in scanchain_197/latch_enable_in scanchain_196/module_data_in[0]
+ scanchain_196/module_data_in[1] scanchain_196/module_data_in[2] scanchain_196/module_data_in[3]
+ scanchain_196/module_data_in[4] scanchain_196/module_data_in[5] scanchain_196/module_data_in[6]
+ scanchain_196/module_data_in[7] scanchain_196/module_data_out[0] scanchain_196/module_data_out[1]
+ scanchain_196/module_data_out[2] scanchain_196/module_data_out[3] scanchain_196/module_data_out[4]
+ scanchain_196/module_data_out[5] scanchain_196/module_data_out[6] scanchain_196/module_data_out[7]
+ scanchain_196/scan_select_in scanchain_197/scan_select_in vccd1 vssd1 scanchain
Xscanchain_130 scanchain_130/clk_in scanchain_131/clk_in scanchain_130/data_in scanchain_131/data_in
+ scanchain_130/latch_enable_in scanchain_131/latch_enable_in scanchain_130/module_data_in[0]
+ scanchain_130/module_data_in[1] scanchain_130/module_data_in[2] scanchain_130/module_data_in[3]
+ scanchain_130/module_data_in[4] scanchain_130/module_data_in[5] scanchain_130/module_data_in[6]
+ scanchain_130/module_data_in[7] scanchain_130/module_data_out[0] scanchain_130/module_data_out[1]
+ scanchain_130/module_data_out[2] scanchain_130/module_data_out[3] scanchain_130/module_data_out[4]
+ scanchain_130/module_data_out[5] scanchain_130/module_data_out[6] scanchain_130/module_data_out[7]
+ scanchain_130/scan_select_in scanchain_131/scan_select_in vccd1 vssd1 scanchain
Xscanchain_141 scanchain_141/clk_in scanchain_142/clk_in scanchain_141/data_in scanchain_142/data_in
+ scanchain_141/latch_enable_in scanchain_142/latch_enable_in scanchain_141/module_data_in[0]
+ scanchain_141/module_data_in[1] scanchain_141/module_data_in[2] scanchain_141/module_data_in[3]
+ scanchain_141/module_data_in[4] scanchain_141/module_data_in[5] scanchain_141/module_data_in[6]
+ scanchain_141/module_data_in[7] scanchain_141/module_data_out[0] scanchain_141/module_data_out[1]
+ scanchain_141/module_data_out[2] scanchain_141/module_data_out[3] scanchain_141/module_data_out[4]
+ scanchain_141/module_data_out[5] scanchain_141/module_data_out[6] scanchain_141/module_data_out[7]
+ scanchain_141/scan_select_in scanchain_142/scan_select_in vccd1 vssd1 scanchain
Xscanchain_152 scanchain_152/clk_in scanchain_153/clk_in scanchain_152/data_in scanchain_153/data_in
+ scanchain_152/latch_enable_in scanchain_153/latch_enable_in scanchain_152/module_data_in[0]
+ scanchain_152/module_data_in[1] scanchain_152/module_data_in[2] scanchain_152/module_data_in[3]
+ scanchain_152/module_data_in[4] scanchain_152/module_data_in[5] scanchain_152/module_data_in[6]
+ scanchain_152/module_data_in[7] scanchain_152/module_data_out[0] scanchain_152/module_data_out[1]
+ scanchain_152/module_data_out[2] scanchain_152/module_data_out[3] scanchain_152/module_data_out[4]
+ scanchain_152/module_data_out[5] scanchain_152/module_data_out[6] scanchain_152/module_data_out[7]
+ scanchain_152/scan_select_in scanchain_153/scan_select_in vccd1 vssd1 scanchain
Xscanchain_163 scanchain_163/clk_in scanchain_164/clk_in scanchain_163/data_in scanchain_164/data_in
+ scanchain_163/latch_enable_in scanchain_164/latch_enable_in scanchain_163/module_data_in[0]
+ scanchain_163/module_data_in[1] scanchain_163/module_data_in[2] scanchain_163/module_data_in[3]
+ scanchain_163/module_data_in[4] scanchain_163/module_data_in[5] scanchain_163/module_data_in[6]
+ scanchain_163/module_data_in[7] scanchain_163/module_data_out[0] scanchain_163/module_data_out[1]
+ scanchain_163/module_data_out[2] scanchain_163/module_data_out[3] scanchain_163/module_data_out[4]
+ scanchain_163/module_data_out[5] scanchain_163/module_data_out[6] scanchain_163/module_data_out[7]
+ scanchain_163/scan_select_in scanchain_164/scan_select_in vccd1 vssd1 scanchain
Xscanchain_185 scanchain_185/clk_in scanchain_186/clk_in scanchain_185/data_in scanchain_186/data_in
+ scanchain_185/latch_enable_in scanchain_186/latch_enable_in scanchain_185/module_data_in[0]
+ scanchain_185/module_data_in[1] scanchain_185/module_data_in[2] scanchain_185/module_data_in[3]
+ scanchain_185/module_data_in[4] scanchain_185/module_data_in[5] scanchain_185/module_data_in[6]
+ scanchain_185/module_data_in[7] scanchain_185/module_data_out[0] scanchain_185/module_data_out[1]
+ scanchain_185/module_data_out[2] scanchain_185/module_data_out[3] scanchain_185/module_data_out[4]
+ scanchain_185/module_data_out[5] scanchain_185/module_data_out[6] scanchain_185/module_data_out[7]
+ scanchain_185/scan_select_in scanchain_186/scan_select_in vccd1 vssd1 scanchain
Xscanchain_174 scanchain_174/clk_in scanchain_175/clk_in scanchain_174/data_in scanchain_175/data_in
+ scanchain_174/latch_enable_in scanchain_175/latch_enable_in scanchain_174/module_data_in[0]
+ scanchain_174/module_data_in[1] scanchain_174/module_data_in[2] scanchain_174/module_data_in[3]
+ scanchain_174/module_data_in[4] scanchain_174/module_data_in[5] scanchain_174/module_data_in[6]
+ scanchain_174/module_data_in[7] scanchain_174/module_data_out[0] scanchain_174/module_data_out[1]
+ scanchain_174/module_data_out[2] scanchain_174/module_data_out[3] scanchain_174/module_data_out[4]
+ scanchain_174/module_data_out[5] scanchain_174/module_data_out[6] scanchain_174/module_data_out[7]
+ scanchain_174/scan_select_in scanchain_175/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_209 scanchain_209/module_data_in[0] scanchain_209/module_data_in[1]
+ scanchain_209/module_data_in[2] scanchain_209/module_data_in[3] scanchain_209/module_data_in[4]
+ scanchain_209/module_data_in[5] scanchain_209/module_data_in[6] scanchain_209/module_data_in[7]
+ scanchain_209/module_data_out[0] scanchain_209/module_data_out[1] scanchain_209/module_data_out[2]
+ scanchain_209/module_data_out[3] scanchain_209/module_data_out[4] scanchain_209/module_data_out[5]
+ scanchain_209/module_data_out[6] scanchain_209/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xxor_shift32_evango_52 xor_shift32_evango_52/io_in[0] xor_shift32_evango_52/io_in[1]
+ xor_shift32_evango_52/io_in[2] xor_shift32_evango_52/io_in[3] xor_shift32_evango_52/io_in[4]
+ xor_shift32_evango_52/io_in[5] xor_shift32_evango_52/io_in[6] xor_shift32_evango_52/io_in[7]
+ xor_shift32_evango_52/io_out[0] xor_shift32_evango_52/io_out[1] xor_shift32_evango_52/io_out[2]
+ xor_shift32_evango_52/io_out[3] xor_shift32_evango_52/io_out[4] xor_shift32_evango_52/io_out[5]
+ xor_shift32_evango_52/io_out[6] xor_shift32_evango_52/io_out[7] vccd1 vssd1 xor_shift32_evango
Xuser_module_339501025136214612_392 scanchain_392/module_data_in[0] scanchain_392/module_data_in[1]
+ scanchain_392/module_data_in[2] scanchain_392/module_data_in[3] scanchain_392/module_data_in[4]
+ scanchain_392/module_data_in[5] scanchain_392/module_data_in[6] scanchain_392/module_data_in[7]
+ scanchain_392/module_data_out[0] scanchain_392/module_data_out[1] scanchain_392/module_data_out[2]
+ scanchain_392/module_data_out[3] scanchain_392/module_data_out[4] scanchain_392/module_data_out[5]
+ scanchain_392/module_data_out[6] scanchain_392/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_389 scanchain_389/clk_in scanchain_390/clk_in scanchain_389/data_in scanchain_390/data_in
+ scanchain_389/latch_enable_in scanchain_390/latch_enable_in scanchain_389/module_data_in[0]
+ scanchain_389/module_data_in[1] scanchain_389/module_data_in[2] scanchain_389/module_data_in[3]
+ scanchain_389/module_data_in[4] scanchain_389/module_data_in[5] scanchain_389/module_data_in[6]
+ scanchain_389/module_data_in[7] scanchain_389/module_data_out[0] scanchain_389/module_data_out[1]
+ scanchain_389/module_data_out[2] scanchain_389/module_data_out[3] scanchain_389/module_data_out[4]
+ scanchain_389/module_data_out[5] scanchain_389/module_data_out[6] scanchain_389/module_data_out[7]
+ scanchain_389/scan_select_in scanchain_390/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_381 scanchain_381/module_data_in[0] scanchain_381/module_data_in[1]
+ scanchain_381/module_data_in[2] scanchain_381/module_data_in[3] scanchain_381/module_data_in[4]
+ scanchain_381/module_data_in[5] scanchain_381/module_data_in[6] scanchain_381/module_data_in[7]
+ scanchain_381/module_data_out[0] scanchain_381/module_data_out[1] scanchain_381/module_data_out[2]
+ scanchain_381/module_data_out[3] scanchain_381/module_data_out[4] scanchain_381/module_data_out[5]
+ scanchain_381/module_data_out[6] scanchain_381/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_378 scanchain_378/clk_in scanchain_379/clk_in scanchain_378/data_in scanchain_379/data_in
+ scanchain_378/latch_enable_in scanchain_379/latch_enable_in scanchain_378/module_data_in[0]
+ scanchain_378/module_data_in[1] scanchain_378/module_data_in[2] scanchain_378/module_data_in[3]
+ scanchain_378/module_data_in[4] scanchain_378/module_data_in[5] scanchain_378/module_data_in[6]
+ scanchain_378/module_data_in[7] scanchain_378/module_data_out[0] scanchain_378/module_data_out[1]
+ scanchain_378/module_data_out[2] scanchain_378/module_data_out[3] scanchain_378/module_data_out[4]
+ scanchain_378/module_data_out[5] scanchain_378/module_data_out[6] scanchain_378/module_data_out[7]
+ scanchain_378/scan_select_in scanchain_379/scan_select_in vccd1 vssd1 scanchain
Xscanchain_367 scanchain_367/clk_in scanchain_368/clk_in scanchain_367/data_in scanchain_368/data_in
+ scanchain_367/latch_enable_in scanchain_368/latch_enable_in scanchain_367/module_data_in[0]
+ scanchain_367/module_data_in[1] scanchain_367/module_data_in[2] scanchain_367/module_data_in[3]
+ scanchain_367/module_data_in[4] scanchain_367/module_data_in[5] scanchain_367/module_data_in[6]
+ scanchain_367/module_data_in[7] scanchain_367/module_data_out[0] scanchain_367/module_data_out[1]
+ scanchain_367/module_data_out[2] scanchain_367/module_data_out[3] scanchain_367/module_data_out[4]
+ scanchain_367/module_data_out[5] scanchain_367/module_data_out[6] scanchain_367/module_data_out[7]
+ scanchain_367/scan_select_in scanchain_368/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_370 scanchain_370/module_data_in[0] scanchain_370/module_data_in[1]
+ scanchain_370/module_data_in[2] scanchain_370/module_data_in[3] scanchain_370/module_data_in[4]
+ scanchain_370/module_data_in[5] scanchain_370/module_data_in[6] scanchain_370/module_data_in[7]
+ scanchain_370/module_data_out[0] scanchain_370/module_data_out[1] scanchain_370/module_data_out[2]
+ scanchain_370/module_data_out[3] scanchain_370/module_data_out[4] scanchain_370/module_data_out[5]
+ scanchain_370/module_data_out[6] scanchain_370/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_356 scanchain_356/clk_in scanchain_357/clk_in scanchain_356/data_in scanchain_357/data_in
+ scanchain_356/latch_enable_in scanchain_357/latch_enable_in scanchain_356/module_data_in[0]
+ scanchain_356/module_data_in[1] scanchain_356/module_data_in[2] scanchain_356/module_data_in[3]
+ scanchain_356/module_data_in[4] scanchain_356/module_data_in[5] scanchain_356/module_data_in[6]
+ scanchain_356/module_data_in[7] scanchain_356/module_data_out[0] scanchain_356/module_data_out[1]
+ scanchain_356/module_data_out[2] scanchain_356/module_data_out[3] scanchain_356/module_data_out[4]
+ scanchain_356/module_data_out[5] scanchain_356/module_data_out[6] scanchain_356/module_data_out[7]
+ scanchain_356/scan_select_in scanchain_357/scan_select_in vccd1 vssd1 scanchain
Xscanchain_345 scanchain_345/clk_in scanchain_346/clk_in scanchain_345/data_in scanchain_346/data_in
+ scanchain_345/latch_enable_in scanchain_346/latch_enable_in scanchain_345/module_data_in[0]
+ scanchain_345/module_data_in[1] scanchain_345/module_data_in[2] scanchain_345/module_data_in[3]
+ scanchain_345/module_data_in[4] scanchain_345/module_data_in[5] scanchain_345/module_data_in[6]
+ scanchain_345/module_data_in[7] scanchain_345/module_data_out[0] scanchain_345/module_data_out[1]
+ scanchain_345/module_data_out[2] scanchain_345/module_data_out[3] scanchain_345/module_data_out[4]
+ scanchain_345/module_data_out[5] scanchain_345/module_data_out[6] scanchain_345/module_data_out[7]
+ scanchain_345/scan_select_in scanchain_346/scan_select_in vccd1 vssd1 scanchain
Xscanchain_323 scanchain_323/clk_in scanchain_324/clk_in scanchain_323/data_in scanchain_324/data_in
+ scanchain_323/latch_enable_in scanchain_324/latch_enable_in scanchain_323/module_data_in[0]
+ scanchain_323/module_data_in[1] scanchain_323/module_data_in[2] scanchain_323/module_data_in[3]
+ scanchain_323/module_data_in[4] scanchain_323/module_data_in[5] scanchain_323/module_data_in[6]
+ scanchain_323/module_data_in[7] scanchain_323/module_data_out[0] scanchain_323/module_data_out[1]
+ scanchain_323/module_data_out[2] scanchain_323/module_data_out[3] scanchain_323/module_data_out[4]
+ scanchain_323/module_data_out[5] scanchain_323/module_data_out[6] scanchain_323/module_data_out[7]
+ scanchain_323/scan_select_in scanchain_324/scan_select_in vccd1 vssd1 scanchain
Xscanchain_334 scanchain_334/clk_in scanchain_335/clk_in scanchain_334/data_in scanchain_335/data_in
+ scanchain_334/latch_enable_in scanchain_335/latch_enable_in scanchain_334/module_data_in[0]
+ scanchain_334/module_data_in[1] scanchain_334/module_data_in[2] scanchain_334/module_data_in[3]
+ scanchain_334/module_data_in[4] scanchain_334/module_data_in[5] scanchain_334/module_data_in[6]
+ scanchain_334/module_data_in[7] scanchain_334/module_data_out[0] scanchain_334/module_data_out[1]
+ scanchain_334/module_data_out[2] scanchain_334/module_data_out[3] scanchain_334/module_data_out[4]
+ scanchain_334/module_data_out[5] scanchain_334/module_data_out[6] scanchain_334/module_data_out[7]
+ scanchain_334/scan_select_in scanchain_335/scan_select_in vccd1 vssd1 scanchain
Xscanchain_312 scanchain_312/clk_in scanchain_313/clk_in scanchain_312/data_in scanchain_313/data_in
+ scanchain_312/latch_enable_in scanchain_313/latch_enable_in scanchain_312/module_data_in[0]
+ scanchain_312/module_data_in[1] scanchain_312/module_data_in[2] scanchain_312/module_data_in[3]
+ scanchain_312/module_data_in[4] scanchain_312/module_data_in[5] scanchain_312/module_data_in[6]
+ scanchain_312/module_data_in[7] scanchain_312/module_data_out[0] scanchain_312/module_data_out[1]
+ scanchain_312/module_data_out[2] scanchain_312/module_data_out[3] scanchain_312/module_data_out[4]
+ scanchain_312/module_data_out[5] scanchain_312/module_data_out[6] scanchain_312/module_data_out[7]
+ scanchain_312/scan_select_in scanchain_313/scan_select_in vccd1 vssd1 scanchain
Xscanchain_301 scanchain_301/clk_in scanchain_302/clk_in scanchain_301/data_in scanchain_302/data_in
+ scanchain_301/latch_enable_in scanchain_302/latch_enable_in scanchain_301/module_data_in[0]
+ scanchain_301/module_data_in[1] scanchain_301/module_data_in[2] scanchain_301/module_data_in[3]
+ scanchain_301/module_data_in[4] scanchain_301/module_data_in[5] scanchain_301/module_data_in[6]
+ scanchain_301/module_data_in[7] scanchain_301/module_data_out[0] scanchain_301/module_data_out[1]
+ scanchain_301/module_data_out[2] scanchain_301/module_data_out[3] scanchain_301/module_data_out[4]
+ scanchain_301/module_data_out[5] scanchain_301/module_data_out[6] scanchain_301/module_data_out[7]
+ scanchain_301/scan_select_in scanchain_302/scan_select_in vccd1 vssd1 scanchain
Xrc5_top_43 rc5_top_43/io_in[0] rc5_top_43/io_in[1] rc5_top_43/io_in[2] rc5_top_43/io_in[3]
+ rc5_top_43/io_in[4] rc5_top_43/io_in[5] rc5_top_43/io_in[6] rc5_top_43/io_in[7]
+ rc5_top_43/io_out[0] rc5_top_43/io_out[1] rc5_top_43/io_out[2] rc5_top_43/io_out[3]
+ rc5_top_43/io_out[4] rc5_top_43/io_out[5] rc5_top_43/io_out[6] rc5_top_43/io_out[7]
+ vccd1 vssd1 rc5_top
Xscanchain_197 scanchain_197/clk_in scanchain_198/clk_in scanchain_197/data_in scanchain_198/data_in
+ scanchain_197/latch_enable_in scanchain_198/latch_enable_in scanchain_197/module_data_in[0]
+ scanchain_197/module_data_in[1] scanchain_197/module_data_in[2] scanchain_197/module_data_in[3]
+ scanchain_197/module_data_in[4] scanchain_197/module_data_in[5] scanchain_197/module_data_in[6]
+ scanchain_197/module_data_in[7] scanchain_197/module_data_out[0] scanchain_197/module_data_out[1]
+ scanchain_197/module_data_out[2] scanchain_197/module_data_out[3] scanchain_197/module_data_out[4]
+ scanchain_197/module_data_out[5] scanchain_197/module_data_out[6] scanchain_197/module_data_out[7]
+ scanchain_197/scan_select_in scanchain_198/scan_select_in vccd1 vssd1 scanchain
Xscanchain_120 scanchain_120/clk_in scanchain_121/clk_in scanchain_120/data_in scanchain_121/data_in
+ scanchain_120/latch_enable_in scanchain_121/latch_enable_in scanchain_120/module_data_in[0]
+ scanchain_120/module_data_in[1] scanchain_120/module_data_in[2] scanchain_120/module_data_in[3]
+ scanchain_120/module_data_in[4] scanchain_120/module_data_in[5] scanchain_120/module_data_in[6]
+ scanchain_120/module_data_in[7] scanchain_120/module_data_out[0] scanchain_120/module_data_out[1]
+ scanchain_120/module_data_out[2] scanchain_120/module_data_out[3] scanchain_120/module_data_out[4]
+ scanchain_120/module_data_out[5] scanchain_120/module_data_out[6] scanchain_120/module_data_out[7]
+ scanchain_120/scan_select_in scanchain_121/scan_select_in vccd1 vssd1 scanchain
Xscanchain_142 scanchain_142/clk_in scanchain_143/clk_in scanchain_142/data_in scanchain_143/data_in
+ scanchain_142/latch_enable_in scanchain_143/latch_enable_in scanchain_142/module_data_in[0]
+ scanchain_142/module_data_in[1] scanchain_142/module_data_in[2] scanchain_142/module_data_in[3]
+ scanchain_142/module_data_in[4] scanchain_142/module_data_in[5] scanchain_142/module_data_in[6]
+ scanchain_142/module_data_in[7] scanchain_142/module_data_out[0] scanchain_142/module_data_out[1]
+ scanchain_142/module_data_out[2] scanchain_142/module_data_out[3] scanchain_142/module_data_out[4]
+ scanchain_142/module_data_out[5] scanchain_142/module_data_out[6] scanchain_142/module_data_out[7]
+ scanchain_142/scan_select_in scanchain_143/scan_select_in vccd1 vssd1 scanchain
Xscanchain_131 scanchain_131/clk_in scanchain_132/clk_in scanchain_131/data_in scanchain_132/data_in
+ scanchain_131/latch_enable_in scanchain_132/latch_enable_in scanchain_131/module_data_in[0]
+ scanchain_131/module_data_in[1] scanchain_131/module_data_in[2] scanchain_131/module_data_in[3]
+ scanchain_131/module_data_in[4] scanchain_131/module_data_in[5] scanchain_131/module_data_in[6]
+ scanchain_131/module_data_in[7] scanchain_131/module_data_out[0] scanchain_131/module_data_out[1]
+ scanchain_131/module_data_out[2] scanchain_131/module_data_out[3] scanchain_131/module_data_out[4]
+ scanchain_131/module_data_out[5] scanchain_131/module_data_out[6] scanchain_131/module_data_out[7]
+ scanchain_131/scan_select_in scanchain_132/scan_select_in vccd1 vssd1 scanchain
Xscanchain_153 scanchain_153/clk_in scanchain_154/clk_in scanchain_153/data_in scanchain_154/data_in
+ scanchain_153/latch_enable_in scanchain_154/latch_enable_in scanchain_153/module_data_in[0]
+ scanchain_153/module_data_in[1] scanchain_153/module_data_in[2] scanchain_153/module_data_in[3]
+ scanchain_153/module_data_in[4] scanchain_153/module_data_in[5] scanchain_153/module_data_in[6]
+ scanchain_153/module_data_in[7] scanchain_153/module_data_out[0] scanchain_153/module_data_out[1]
+ scanchain_153/module_data_out[2] scanchain_153/module_data_out[3] scanchain_153/module_data_out[4]
+ scanchain_153/module_data_out[5] scanchain_153/module_data_out[6] scanchain_153/module_data_out[7]
+ scanchain_153/scan_select_in scanchain_154/scan_select_in vccd1 vssd1 scanchain
Xscanchain_164 scanchain_164/clk_in scanchain_165/clk_in scanchain_164/data_in scanchain_165/data_in
+ scanchain_164/latch_enable_in scanchain_165/latch_enable_in scanchain_164/module_data_in[0]
+ scanchain_164/module_data_in[1] scanchain_164/module_data_in[2] scanchain_164/module_data_in[3]
+ scanchain_164/module_data_in[4] scanchain_164/module_data_in[5] scanchain_164/module_data_in[6]
+ scanchain_164/module_data_in[7] scanchain_164/module_data_out[0] scanchain_164/module_data_out[1]
+ scanchain_164/module_data_out[2] scanchain_164/module_data_out[3] scanchain_164/module_data_out[4]
+ scanchain_164/module_data_out[5] scanchain_164/module_data_out[6] scanchain_164/module_data_out[7]
+ scanchain_164/scan_select_in scanchain_165/scan_select_in vccd1 vssd1 scanchain
Xscanchain_186 scanchain_186/clk_in scanchain_187/clk_in scanchain_186/data_in scanchain_187/data_in
+ scanchain_186/latch_enable_in scanchain_187/latch_enable_in scanchain_186/module_data_in[0]
+ scanchain_186/module_data_in[1] scanchain_186/module_data_in[2] scanchain_186/module_data_in[3]
+ scanchain_186/module_data_in[4] scanchain_186/module_data_in[5] scanchain_186/module_data_in[6]
+ scanchain_186/module_data_in[7] scanchain_186/module_data_out[0] scanchain_186/module_data_out[1]
+ scanchain_186/module_data_out[2] scanchain_186/module_data_out[3] scanchain_186/module_data_out[4]
+ scanchain_186/module_data_out[5] scanchain_186/module_data_out[6] scanchain_186/module_data_out[7]
+ scanchain_186/scan_select_in scanchain_187/scan_select_in vccd1 vssd1 scanchain
Xscanchain_175 scanchain_175/clk_in scanchain_176/clk_in scanchain_175/data_in scanchain_176/data_in
+ scanchain_175/latch_enable_in scanchain_176/latch_enable_in scanchain_175/module_data_in[0]
+ scanchain_175/module_data_in[1] scanchain_175/module_data_in[2] scanchain_175/module_data_in[3]
+ scanchain_175/module_data_in[4] scanchain_175/module_data_in[5] scanchain_175/module_data_in[6]
+ scanchain_175/module_data_in[7] scanchain_175/module_data_out[0] scanchain_175/module_data_out[1]
+ scanchain_175/module_data_out[2] scanchain_175/module_data_out[3] scanchain_175/module_data_out[4]
+ scanchain_175/module_data_out[5] scanchain_175/module_data_out[6] scanchain_175/module_data_out[7]
+ scanchain_175/scan_select_in scanchain_176/scan_select_in vccd1 vssd1 scanchain
Xtt2_tholin_multiplier_49 scanchain_49/module_data_in[0] scanchain_49/module_data_in[1]
+ scanchain_49/module_data_in[2] scanchain_49/module_data_in[3] scanchain_49/module_data_in[4]
+ scanchain_49/module_data_in[5] scanchain_49/module_data_in[6] scanchain_49/module_data_in[7]
+ scanchain_49/module_data_out[0] scanchain_49/module_data_out[1] scanchain_49/module_data_out[2]
+ scanchain_49/module_data_out[3] scanchain_49/module_data_out[4] scanchain_49/module_data_out[5]
+ scanchain_49/module_data_out[6] scanchain_49/module_data_out[7] vccd1 vssd1 tt2_tholin_multiplier
Xuser_module_346916357828248146_18 scanchain_18/module_data_in[0] scanchain_18/module_data_in[1]
+ scanchain_18/module_data_in[2] scanchain_18/module_data_in[3] scanchain_18/module_data_in[4]
+ scanchain_18/module_data_in[5] scanchain_18/module_data_in[6] scanchain_18/module_data_in[7]
+ scanchain_18/module_data_out[0] scanchain_18/module_data_out[1] scanchain_18/module_data_out[2]
+ scanchain_18/module_data_out[3] scanchain_18/module_data_out[4] scanchain_18/module_data_out[5]
+ scanchain_18/module_data_out[6] scanchain_18/module_data_out[7] vccd1 vssd1 user_module_346916357828248146
Xuser_module_339501025136214612_393 scanchain_393/module_data_in[0] scanchain_393/module_data_in[1]
+ scanchain_393/module_data_in[2] scanchain_393/module_data_in[3] scanchain_393/module_data_in[4]
+ scanchain_393/module_data_in[5] scanchain_393/module_data_in[6] scanchain_393/module_data_in[7]
+ scanchain_393/module_data_out[0] scanchain_393/module_data_out[1] scanchain_393/module_data_out[2]
+ scanchain_393/module_data_out[3] scanchain_393/module_data_out[4] scanchain_393/module_data_out[5]
+ scanchain_393/module_data_out[6] scanchain_393/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_382 scanchain_382/module_data_in[0] scanchain_382/module_data_in[1]
+ scanchain_382/module_data_in[2] scanchain_382/module_data_in[3] scanchain_382/module_data_in[4]
+ scanchain_382/module_data_in[5] scanchain_382/module_data_in[6] scanchain_382/module_data_in[7]
+ scanchain_382/module_data_out[0] scanchain_382/module_data_out[1] scanchain_382/module_data_out[2]
+ scanchain_382/module_data_out[3] scanchain_382/module_data_out[4] scanchain_382/module_data_out[5]
+ scanchain_382/module_data_out[6] scanchain_382/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_360 scanchain_360/module_data_in[0] scanchain_360/module_data_in[1]
+ scanchain_360/module_data_in[2] scanchain_360/module_data_in[3] scanchain_360/module_data_in[4]
+ scanchain_360/module_data_in[5] scanchain_360/module_data_in[6] scanchain_360/module_data_in[7]
+ scanchain_360/module_data_out[0] scanchain_360/module_data_out[1] scanchain_360/module_data_out[2]
+ scanchain_360/module_data_out[3] scanchain_360/module_data_out[4] scanchain_360/module_data_out[5]
+ scanchain_360/module_data_out[6] scanchain_360/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_371 scanchain_371/module_data_in[0] scanchain_371/module_data_in[1]
+ scanchain_371/module_data_in[2] scanchain_371/module_data_in[3] scanchain_371/module_data_in[4]
+ scanchain_371/module_data_in[5] scanchain_371/module_data_in[6] scanchain_371/module_data_in[7]
+ scanchain_371/module_data_out[0] scanchain_371/module_data_out[1] scanchain_371/module_data_out[2]
+ scanchain_371/module_data_out[3] scanchain_371/module_data_out[4] scanchain_371/module_data_out[5]
+ scanchain_371/module_data_out[6] scanchain_371/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_379 scanchain_379/clk_in scanchain_380/clk_in scanchain_379/data_in scanchain_380/data_in
+ scanchain_379/latch_enable_in scanchain_380/latch_enable_in scanchain_379/module_data_in[0]
+ scanchain_379/module_data_in[1] scanchain_379/module_data_in[2] scanchain_379/module_data_in[3]
+ scanchain_379/module_data_in[4] scanchain_379/module_data_in[5] scanchain_379/module_data_in[6]
+ scanchain_379/module_data_in[7] scanchain_379/module_data_out[0] scanchain_379/module_data_out[1]
+ scanchain_379/module_data_out[2] scanchain_379/module_data_out[3] scanchain_379/module_data_out[4]
+ scanchain_379/module_data_out[5] scanchain_379/module_data_out[6] scanchain_379/module_data_out[7]
+ scanchain_379/scan_select_in scanchain_380/scan_select_in vccd1 vssd1 scanchain
Xscanchain_368 scanchain_368/clk_in scanchain_369/clk_in scanchain_368/data_in scanchain_369/data_in
+ scanchain_368/latch_enable_in scanchain_369/latch_enable_in scanchain_368/module_data_in[0]
+ scanchain_368/module_data_in[1] scanchain_368/module_data_in[2] scanchain_368/module_data_in[3]
+ scanchain_368/module_data_in[4] scanchain_368/module_data_in[5] scanchain_368/module_data_in[6]
+ scanchain_368/module_data_in[7] scanchain_368/module_data_out[0] scanchain_368/module_data_out[1]
+ scanchain_368/module_data_out[2] scanchain_368/module_data_out[3] scanchain_368/module_data_out[4]
+ scanchain_368/module_data_out[5] scanchain_368/module_data_out[6] scanchain_368/module_data_out[7]
+ scanchain_368/scan_select_in scanchain_369/scan_select_in vccd1 vssd1 scanchain
Xscanchain_357 scanchain_357/clk_in scanchain_358/clk_in scanchain_357/data_in scanchain_358/data_in
+ scanchain_357/latch_enable_in scanchain_358/latch_enable_in scanchain_357/module_data_in[0]
+ scanchain_357/module_data_in[1] scanchain_357/module_data_in[2] scanchain_357/module_data_in[3]
+ scanchain_357/module_data_in[4] scanchain_357/module_data_in[5] scanchain_357/module_data_in[6]
+ scanchain_357/module_data_in[7] scanchain_357/module_data_out[0] scanchain_357/module_data_out[1]
+ scanchain_357/module_data_out[2] scanchain_357/module_data_out[3] scanchain_357/module_data_out[4]
+ scanchain_357/module_data_out[5] scanchain_357/module_data_out[6] scanchain_357/module_data_out[7]
+ scanchain_357/scan_select_in scanchain_358/scan_select_in vccd1 vssd1 scanchain
Xscanchain_346 scanchain_346/clk_in scanchain_347/clk_in scanchain_346/data_in scanchain_347/data_in
+ scanchain_346/latch_enable_in scanchain_347/latch_enable_in scanchain_346/module_data_in[0]
+ scanchain_346/module_data_in[1] scanchain_346/module_data_in[2] scanchain_346/module_data_in[3]
+ scanchain_346/module_data_in[4] scanchain_346/module_data_in[5] scanchain_346/module_data_in[6]
+ scanchain_346/module_data_in[7] scanchain_346/module_data_out[0] scanchain_346/module_data_out[1]
+ scanchain_346/module_data_out[2] scanchain_346/module_data_out[3] scanchain_346/module_data_out[4]
+ scanchain_346/module_data_out[5] scanchain_346/module_data_out[6] scanchain_346/module_data_out[7]
+ scanchain_346/scan_select_in scanchain_347/scan_select_in vccd1 vssd1 scanchain
Xscanchain_324 scanchain_324/clk_in scanchain_325/clk_in scanchain_324/data_in scanchain_325/data_in
+ scanchain_324/latch_enable_in scanchain_325/latch_enable_in scanchain_324/module_data_in[0]
+ scanchain_324/module_data_in[1] scanchain_324/module_data_in[2] scanchain_324/module_data_in[3]
+ scanchain_324/module_data_in[4] scanchain_324/module_data_in[5] scanchain_324/module_data_in[6]
+ scanchain_324/module_data_in[7] scanchain_324/module_data_out[0] scanchain_324/module_data_out[1]
+ scanchain_324/module_data_out[2] scanchain_324/module_data_out[3] scanchain_324/module_data_out[4]
+ scanchain_324/module_data_out[5] scanchain_324/module_data_out[6] scanchain_324/module_data_out[7]
+ scanchain_324/scan_select_in scanchain_325/scan_select_in vccd1 vssd1 scanchain
Xscanchain_335 scanchain_335/clk_in scanchain_336/clk_in scanchain_335/data_in scanchain_336/data_in
+ scanchain_335/latch_enable_in scanchain_336/latch_enable_in scanchain_335/module_data_in[0]
+ scanchain_335/module_data_in[1] scanchain_335/module_data_in[2] scanchain_335/module_data_in[3]
+ scanchain_335/module_data_in[4] scanchain_335/module_data_in[5] scanchain_335/module_data_in[6]
+ scanchain_335/module_data_in[7] scanchain_335/module_data_out[0] scanchain_335/module_data_out[1]
+ scanchain_335/module_data_out[2] scanchain_335/module_data_out[3] scanchain_335/module_data_out[4]
+ scanchain_335/module_data_out[5] scanchain_335/module_data_out[6] scanchain_335/module_data_out[7]
+ scanchain_335/scan_select_in scanchain_336/scan_select_in vccd1 vssd1 scanchain
Xscanchain_313 scanchain_313/clk_in scanchain_314/clk_in scanchain_313/data_in scanchain_314/data_in
+ scanchain_313/latch_enable_in scanchain_314/latch_enable_in scanchain_313/module_data_in[0]
+ scanchain_313/module_data_in[1] scanchain_313/module_data_in[2] scanchain_313/module_data_in[3]
+ scanchain_313/module_data_in[4] scanchain_313/module_data_in[5] scanchain_313/module_data_in[6]
+ scanchain_313/module_data_in[7] scanchain_313/module_data_out[0] scanchain_313/module_data_out[1]
+ scanchain_313/module_data_out[2] scanchain_313/module_data_out[3] scanchain_313/module_data_out[4]
+ scanchain_313/module_data_out[5] scanchain_313/module_data_out[6] scanchain_313/module_data_out[7]
+ scanchain_313/scan_select_in scanchain_314/scan_select_in vccd1 vssd1 scanchain
Xscanchain_302 scanchain_302/clk_in scanchain_303/clk_in scanchain_302/data_in scanchain_303/data_in
+ scanchain_302/latch_enable_in scanchain_303/latch_enable_in scanchain_302/module_data_in[0]
+ scanchain_302/module_data_in[1] scanchain_302/module_data_in[2] scanchain_302/module_data_in[3]
+ scanchain_302/module_data_in[4] scanchain_302/module_data_in[5] scanchain_302/module_data_in[6]
+ scanchain_302/module_data_in[7] scanchain_302/module_data_out[0] scanchain_302/module_data_out[1]
+ scanchain_302/module_data_out[2] scanchain_302/module_data_out[3] scanchain_302/module_data_out[4]
+ scanchain_302/module_data_out[5] scanchain_302/module_data_out[6] scanchain_302/module_data_out[7]
+ scanchain_302/scan_select_in scanchain_303/scan_select_in vccd1 vssd1 scanchain
Xscanchain_198 scanchain_198/clk_in scanchain_199/clk_in scanchain_198/data_in scanchain_199/data_in
+ scanchain_198/latch_enable_in scanchain_199/latch_enable_in scanchain_198/module_data_in[0]
+ scanchain_198/module_data_in[1] scanchain_198/module_data_in[2] scanchain_198/module_data_in[3]
+ scanchain_198/module_data_in[4] scanchain_198/module_data_in[5] scanchain_198/module_data_in[6]
+ scanchain_198/module_data_in[7] scanchain_198/module_data_out[0] scanchain_198/module_data_out[1]
+ scanchain_198/module_data_out[2] scanchain_198/module_data_out[3] scanchain_198/module_data_out[4]
+ scanchain_198/module_data_out[5] scanchain_198/module_data_out[6] scanchain_198/module_data_out[7]
+ scanchain_198/scan_select_in scanchain_199/scan_select_in vccd1 vssd1 scanchain
Xscanchain_110 scanchain_110/clk_in scanchain_111/clk_in scanchain_110/data_in scanchain_111/data_in
+ scanchain_110/latch_enable_in scanchain_111/latch_enable_in scanchain_110/module_data_in[0]
+ scanchain_110/module_data_in[1] scanchain_110/module_data_in[2] scanchain_110/module_data_in[3]
+ scanchain_110/module_data_in[4] scanchain_110/module_data_in[5] scanchain_110/module_data_in[6]
+ scanchain_110/module_data_in[7] scanchain_110/module_data_out[0] scanchain_110/module_data_out[1]
+ scanchain_110/module_data_out[2] scanchain_110/module_data_out[3] scanchain_110/module_data_out[4]
+ scanchain_110/module_data_out[5] scanchain_110/module_data_out[6] scanchain_110/module_data_out[7]
+ scanchain_110/scan_select_in scanchain_111/scan_select_in vccd1 vssd1 scanchain
Xscanchain_121 scanchain_121/clk_in scanchain_122/clk_in scanchain_121/data_in scanchain_122/data_in
+ scanchain_121/latch_enable_in scanchain_122/latch_enable_in scanchain_121/module_data_in[0]
+ scanchain_121/module_data_in[1] scanchain_121/module_data_in[2] scanchain_121/module_data_in[3]
+ scanchain_121/module_data_in[4] scanchain_121/module_data_in[5] scanchain_121/module_data_in[6]
+ scanchain_121/module_data_in[7] scanchain_121/module_data_out[0] scanchain_121/module_data_out[1]
+ scanchain_121/module_data_out[2] scanchain_121/module_data_out[3] scanchain_121/module_data_out[4]
+ scanchain_121/module_data_out[5] scanchain_121/module_data_out[6] scanchain_121/module_data_out[7]
+ scanchain_121/scan_select_in scanchain_122/scan_select_in vccd1 vssd1 scanchain
Xscanchain_143 scanchain_143/clk_in scanchain_144/clk_in scanchain_143/data_in scanchain_144/data_in
+ scanchain_143/latch_enable_in scanchain_144/latch_enable_in scanchain_143/module_data_in[0]
+ scanchain_143/module_data_in[1] scanchain_143/module_data_in[2] scanchain_143/module_data_in[3]
+ scanchain_143/module_data_in[4] scanchain_143/module_data_in[5] scanchain_143/module_data_in[6]
+ scanchain_143/module_data_in[7] scanchain_143/module_data_out[0] scanchain_143/module_data_out[1]
+ scanchain_143/module_data_out[2] scanchain_143/module_data_out[3] scanchain_143/module_data_out[4]
+ scanchain_143/module_data_out[5] scanchain_143/module_data_out[6] scanchain_143/module_data_out[7]
+ scanchain_143/scan_select_in scanchain_144/scan_select_in vccd1 vssd1 scanchain
Xscanchain_132 scanchain_132/clk_in scanchain_133/clk_in scanchain_132/data_in scanchain_133/data_in
+ scanchain_132/latch_enable_in scanchain_133/latch_enable_in scanchain_132/module_data_in[0]
+ scanchain_132/module_data_in[1] scanchain_132/module_data_in[2] scanchain_132/module_data_in[3]
+ scanchain_132/module_data_in[4] scanchain_132/module_data_in[5] scanchain_132/module_data_in[6]
+ scanchain_132/module_data_in[7] scanchain_132/module_data_out[0] scanchain_132/module_data_out[1]
+ scanchain_132/module_data_out[2] scanchain_132/module_data_out[3] scanchain_132/module_data_out[4]
+ scanchain_132/module_data_out[5] scanchain_132/module_data_out[6] scanchain_132/module_data_out[7]
+ scanchain_132/scan_select_in scanchain_133/scan_select_in vccd1 vssd1 scanchain
Xscanchain_154 scanchain_154/clk_in scanchain_155/clk_in scanchain_154/data_in scanchain_155/data_in
+ scanchain_154/latch_enable_in scanchain_155/latch_enable_in scanchain_154/module_data_in[0]
+ scanchain_154/module_data_in[1] scanchain_154/module_data_in[2] scanchain_154/module_data_in[3]
+ scanchain_154/module_data_in[4] scanchain_154/module_data_in[5] scanchain_154/module_data_in[6]
+ scanchain_154/module_data_in[7] scanchain_154/module_data_out[0] scanchain_154/module_data_out[1]
+ scanchain_154/module_data_out[2] scanchain_154/module_data_out[3] scanchain_154/module_data_out[4]
+ scanchain_154/module_data_out[5] scanchain_154/module_data_out[6] scanchain_154/module_data_out[7]
+ scanchain_154/scan_select_in scanchain_155/scan_select_in vccd1 vssd1 scanchain
Xscanchain_165 scanchain_165/clk_in scanchain_166/clk_in scanchain_165/data_in scanchain_166/data_in
+ scanchain_165/latch_enable_in scanchain_166/latch_enable_in scanchain_165/module_data_in[0]
+ scanchain_165/module_data_in[1] scanchain_165/module_data_in[2] scanchain_165/module_data_in[3]
+ scanchain_165/module_data_in[4] scanchain_165/module_data_in[5] scanchain_165/module_data_in[6]
+ scanchain_165/module_data_in[7] scanchain_165/module_data_out[0] scanchain_165/module_data_out[1]
+ scanchain_165/module_data_out[2] scanchain_165/module_data_out[3] scanchain_165/module_data_out[4]
+ scanchain_165/module_data_out[5] scanchain_165/module_data_out[6] scanchain_165/module_data_out[7]
+ scanchain_165/scan_select_in scanchain_166/scan_select_in vccd1 vssd1 scanchain
Xscanchain_187 scanchain_187/clk_in scanchain_188/clk_in scanchain_187/data_in scanchain_188/data_in
+ scanchain_187/latch_enable_in scanchain_188/latch_enable_in scanchain_187/module_data_in[0]
+ scanchain_187/module_data_in[1] scanchain_187/module_data_in[2] scanchain_187/module_data_in[3]
+ scanchain_187/module_data_in[4] scanchain_187/module_data_in[5] scanchain_187/module_data_in[6]
+ scanchain_187/module_data_in[7] scanchain_187/module_data_out[0] scanchain_187/module_data_out[1]
+ scanchain_187/module_data_out[2] scanchain_187/module_data_out[3] scanchain_187/module_data_out[4]
+ scanchain_187/module_data_out[5] scanchain_187/module_data_out[6] scanchain_187/module_data_out[7]
+ scanchain_187/scan_select_in scanchain_188/scan_select_in vccd1 vssd1 scanchain
Xscanchain_176 scanchain_176/clk_in scanchain_177/clk_in scanchain_176/data_in scanchain_177/data_in
+ scanchain_176/latch_enable_in scanchain_177/latch_enable_in scanchain_176/module_data_in[0]
+ scanchain_176/module_data_in[1] scanchain_176/module_data_in[2] scanchain_176/module_data_in[3]
+ scanchain_176/module_data_in[4] scanchain_176/module_data_in[5] scanchain_176/module_data_in[6]
+ scanchain_176/module_data_in[7] scanchain_176/module_data_out[0] scanchain_176/module_data_out[1]
+ scanchain_176/module_data_out[2] scanchain_176/module_data_out[3] scanchain_176/module_data_out[4]
+ scanchain_176/module_data_out[5] scanchain_176/module_data_out[6] scanchain_176/module_data_out[7]
+ scanchain_176/scan_select_in scanchain_177/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_190 scanchain_190/module_data_in[0] scanchain_190/module_data_in[1]
+ scanchain_190/module_data_in[2] scanchain_190/module_data_in[3] scanchain_190/module_data_in[4]
+ scanchain_190/module_data_in[5] scanchain_190/module_data_in[6] scanchain_190/module_data_in[7]
+ scanchain_190/module_data_out[0] scanchain_190/module_data_out[1] scanchain_190/module_data_out[2]
+ scanchain_190/module_data_out[3] scanchain_190/module_data_out[4] scanchain_190/module_data_out[5]
+ scanchain_190/module_data_out[6] scanchain_190/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xchrisruk_matrix_3 chrisruk_matrix_3/io_in[0] chrisruk_matrix_3/io_in[1] chrisruk_matrix_3/io_in[2]
+ chrisruk_matrix_3/io_in[3] chrisruk_matrix_3/io_in[4] chrisruk_matrix_3/io_in[5]
+ chrisruk_matrix_3/io_in[6] chrisruk_matrix_3/io_in[7] chrisruk_matrix_3/io_out[0]
+ chrisruk_matrix_3/io_out[1] chrisruk_matrix_3/io_out[2] chrisruk_matrix_3/io_out[3]
+ chrisruk_matrix_3/io_out[4] chrisruk_matrix_3/io_out[5] chrisruk_matrix_3/io_out[6]
+ chrisruk_matrix_3/io_out[7] vccd1 vssd1 chrisruk_matrix
Xuser_module_339501025136214612_394 scanchain_394/module_data_in[0] scanchain_394/module_data_in[1]
+ scanchain_394/module_data_in[2] scanchain_394/module_data_in[3] scanchain_394/module_data_in[4]
+ scanchain_394/module_data_in[5] scanchain_394/module_data_in[6] scanchain_394/module_data_in[7]
+ scanchain_394/module_data_out[0] scanchain_394/module_data_out[1] scanchain_394/module_data_out[2]
+ scanchain_394/module_data_out[3] scanchain_394/module_data_out[4] scanchain_394/module_data_out[5]
+ scanchain_394/module_data_out[6] scanchain_394/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_383 scanchain_383/module_data_in[0] scanchain_383/module_data_in[1]
+ scanchain_383/module_data_in[2] scanchain_383/module_data_in[3] scanchain_383/module_data_in[4]
+ scanchain_383/module_data_in[5] scanchain_383/module_data_in[6] scanchain_383/module_data_in[7]
+ scanchain_383/module_data_out[0] scanchain_383/module_data_out[1] scanchain_383/module_data_out[2]
+ scanchain_383/module_data_out[3] scanchain_383/module_data_out[4] scanchain_383/module_data_out[5]
+ scanchain_383/module_data_out[6] scanchain_383/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_361 scanchain_361/module_data_in[0] scanchain_361/module_data_in[1]
+ scanchain_361/module_data_in[2] scanchain_361/module_data_in[3] scanchain_361/module_data_in[4]
+ scanchain_361/module_data_in[5] scanchain_361/module_data_in[6] scanchain_361/module_data_in[7]
+ scanchain_361/module_data_out[0] scanchain_361/module_data_out[1] scanchain_361/module_data_out[2]
+ scanchain_361/module_data_out[3] scanchain_361/module_data_out[4] scanchain_361/module_data_out[5]
+ scanchain_361/module_data_out[6] scanchain_361/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_372 scanchain_372/module_data_in[0] scanchain_372/module_data_in[1]
+ scanchain_372/module_data_in[2] scanchain_372/module_data_in[3] scanchain_372/module_data_in[4]
+ scanchain_372/module_data_in[5] scanchain_372/module_data_in[6] scanchain_372/module_data_in[7]
+ scanchain_372/module_data_out[0] scanchain_372/module_data_out[1] scanchain_372/module_data_out[2]
+ scanchain_372/module_data_out[3] scanchain_372/module_data_out[4] scanchain_372/module_data_out[5]
+ scanchain_372/module_data_out[6] scanchain_372/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_350 scanchain_350/module_data_in[0] scanchain_350/module_data_in[1]
+ scanchain_350/module_data_in[2] scanchain_350/module_data_in[3] scanchain_350/module_data_in[4]
+ scanchain_350/module_data_in[5] scanchain_350/module_data_in[6] scanchain_350/module_data_in[7]
+ scanchain_350/module_data_out[0] scanchain_350/module_data_out[1] scanchain_350/module_data_out[2]
+ scanchain_350/module_data_out[3] scanchain_350/module_data_out[4] scanchain_350/module_data_out[5]
+ scanchain_350/module_data_out[6] scanchain_350/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_369 scanchain_369/clk_in scanchain_370/clk_in scanchain_369/data_in scanchain_370/data_in
+ scanchain_369/latch_enable_in scanchain_370/latch_enable_in scanchain_369/module_data_in[0]
+ scanchain_369/module_data_in[1] scanchain_369/module_data_in[2] scanchain_369/module_data_in[3]
+ scanchain_369/module_data_in[4] scanchain_369/module_data_in[5] scanchain_369/module_data_in[6]
+ scanchain_369/module_data_in[7] scanchain_369/module_data_out[0] scanchain_369/module_data_out[1]
+ scanchain_369/module_data_out[2] scanchain_369/module_data_out[3] scanchain_369/module_data_out[4]
+ scanchain_369/module_data_out[5] scanchain_369/module_data_out[6] scanchain_369/module_data_out[7]
+ scanchain_369/scan_select_in scanchain_370/scan_select_in vccd1 vssd1 scanchain
Xscanchain_358 scanchain_358/clk_in scanchain_359/clk_in scanchain_358/data_in scanchain_359/data_in
+ scanchain_358/latch_enable_in scanchain_359/latch_enable_in scanchain_358/module_data_in[0]
+ scanchain_358/module_data_in[1] scanchain_358/module_data_in[2] scanchain_358/module_data_in[3]
+ scanchain_358/module_data_in[4] scanchain_358/module_data_in[5] scanchain_358/module_data_in[6]
+ scanchain_358/module_data_in[7] scanchain_358/module_data_out[0] scanchain_358/module_data_out[1]
+ scanchain_358/module_data_out[2] scanchain_358/module_data_out[3] scanchain_358/module_data_out[4]
+ scanchain_358/module_data_out[5] scanchain_358/module_data_out[6] scanchain_358/module_data_out[7]
+ scanchain_358/scan_select_in scanchain_359/scan_select_in vccd1 vssd1 scanchain
Xscanchain_347 scanchain_347/clk_in scanchain_348/clk_in scanchain_347/data_in scanchain_348/data_in
+ scanchain_347/latch_enable_in scanchain_348/latch_enable_in scanchain_347/module_data_in[0]
+ scanchain_347/module_data_in[1] scanchain_347/module_data_in[2] scanchain_347/module_data_in[3]
+ scanchain_347/module_data_in[4] scanchain_347/module_data_in[5] scanchain_347/module_data_in[6]
+ scanchain_347/module_data_in[7] scanchain_347/module_data_out[0] scanchain_347/module_data_out[1]
+ scanchain_347/module_data_out[2] scanchain_347/module_data_out[3] scanchain_347/module_data_out[4]
+ scanchain_347/module_data_out[5] scanchain_347/module_data_out[6] scanchain_347/module_data_out[7]
+ scanchain_347/scan_select_in scanchain_348/scan_select_in vccd1 vssd1 scanchain
Xscanchain_325 scanchain_325/clk_in scanchain_326/clk_in scanchain_325/data_in scanchain_326/data_in
+ scanchain_325/latch_enable_in scanchain_326/latch_enable_in scanchain_325/module_data_in[0]
+ scanchain_325/module_data_in[1] scanchain_325/module_data_in[2] scanchain_325/module_data_in[3]
+ scanchain_325/module_data_in[4] scanchain_325/module_data_in[5] scanchain_325/module_data_in[6]
+ scanchain_325/module_data_in[7] scanchain_325/module_data_out[0] scanchain_325/module_data_out[1]
+ scanchain_325/module_data_out[2] scanchain_325/module_data_out[3] scanchain_325/module_data_out[4]
+ scanchain_325/module_data_out[5] scanchain_325/module_data_out[6] scanchain_325/module_data_out[7]
+ scanchain_325/scan_select_in scanchain_326/scan_select_in vccd1 vssd1 scanchain
Xscanchain_336 scanchain_336/clk_in scanchain_337/clk_in scanchain_336/data_in scanchain_337/data_in
+ scanchain_336/latch_enable_in scanchain_337/latch_enable_in scanchain_336/module_data_in[0]
+ scanchain_336/module_data_in[1] scanchain_336/module_data_in[2] scanchain_336/module_data_in[3]
+ scanchain_336/module_data_in[4] scanchain_336/module_data_in[5] scanchain_336/module_data_in[6]
+ scanchain_336/module_data_in[7] scanchain_336/module_data_out[0] scanchain_336/module_data_out[1]
+ scanchain_336/module_data_out[2] scanchain_336/module_data_out[3] scanchain_336/module_data_out[4]
+ scanchain_336/module_data_out[5] scanchain_336/module_data_out[6] scanchain_336/module_data_out[7]
+ scanchain_336/scan_select_in scanchain_337/scan_select_in vccd1 vssd1 scanchain
Xscanchain_314 scanchain_314/clk_in scanchain_315/clk_in scanchain_314/data_in scanchain_315/data_in
+ scanchain_314/latch_enable_in scanchain_315/latch_enable_in scanchain_314/module_data_in[0]
+ scanchain_314/module_data_in[1] scanchain_314/module_data_in[2] scanchain_314/module_data_in[3]
+ scanchain_314/module_data_in[4] scanchain_314/module_data_in[5] scanchain_314/module_data_in[6]
+ scanchain_314/module_data_in[7] scanchain_314/module_data_out[0] scanchain_314/module_data_out[1]
+ scanchain_314/module_data_out[2] scanchain_314/module_data_out[3] scanchain_314/module_data_out[4]
+ scanchain_314/module_data_out[5] scanchain_314/module_data_out[6] scanchain_314/module_data_out[7]
+ scanchain_314/scan_select_in scanchain_315/scan_select_in vccd1 vssd1 scanchain
Xscanchain_303 scanchain_303/clk_in scanchain_304/clk_in scanchain_303/data_in scanchain_304/data_in
+ scanchain_303/latch_enable_in scanchain_304/latch_enable_in scanchain_303/module_data_in[0]
+ scanchain_303/module_data_in[1] scanchain_303/module_data_in[2] scanchain_303/module_data_in[3]
+ scanchain_303/module_data_in[4] scanchain_303/module_data_in[5] scanchain_303/module_data_in[6]
+ scanchain_303/module_data_in[7] scanchain_303/module_data_out[0] scanchain_303/module_data_out[1]
+ scanchain_303/module_data_out[2] scanchain_303/module_data_out[3] scanchain_303/module_data_out[4]
+ scanchain_303/module_data_out[5] scanchain_303/module_data_out[6] scanchain_303/module_data_out[7]
+ scanchain_303/scan_select_in scanchain_304/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_191 scanchain_191/module_data_in[0] scanchain_191/module_data_in[1]
+ scanchain_191/module_data_in[2] scanchain_191/module_data_in[3] scanchain_191/module_data_in[4]
+ scanchain_191/module_data_in[5] scanchain_191/module_data_in[6] scanchain_191/module_data_in[7]
+ scanchain_191/module_data_out[0] scanchain_191/module_data_out[1] scanchain_191/module_data_out[2]
+ scanchain_191/module_data_out[3] scanchain_191/module_data_out[4] scanchain_191/module_data_out[5]
+ scanchain_191/module_data_out[6] scanchain_191/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_111 scanchain_111/clk_in scanchain_112/clk_in scanchain_111/data_in scanchain_112/data_in
+ scanchain_111/latch_enable_in scanchain_112/latch_enable_in scanchain_111/module_data_in[0]
+ scanchain_111/module_data_in[1] scanchain_111/module_data_in[2] scanchain_111/module_data_in[3]
+ scanchain_111/module_data_in[4] scanchain_111/module_data_in[5] scanchain_111/module_data_in[6]
+ scanchain_111/module_data_in[7] scanchain_111/module_data_out[0] scanchain_111/module_data_out[1]
+ scanchain_111/module_data_out[2] scanchain_111/module_data_out[3] scanchain_111/module_data_out[4]
+ scanchain_111/module_data_out[5] scanchain_111/module_data_out[6] scanchain_111/module_data_out[7]
+ scanchain_111/scan_select_in scanchain_112/scan_select_in vccd1 vssd1 scanchain
Xscanchain_100 scanchain_99/clk_out scanchain_101/clk_in scanchain_99/data_out scanchain_101/data_in
+ scanchain_99/latch_enable_out scanchain_101/latch_enable_in scanchain_100/module_data_in[0]
+ scanchain_100/module_data_in[1] scanchain_100/module_data_in[2] scanchain_100/module_data_in[3]
+ scanchain_100/module_data_in[4] scanchain_100/module_data_in[5] scanchain_100/module_data_in[6]
+ scanchain_100/module_data_in[7] scanchain_100/module_data_out[0] scanchain_100/module_data_out[1]
+ scanchain_100/module_data_out[2] scanchain_100/module_data_out[3] scanchain_100/module_data_out[4]
+ scanchain_100/module_data_out[5] scanchain_100/module_data_out[6] scanchain_100/module_data_out[7]
+ scanchain_99/scan_select_out scanchain_101/scan_select_in vccd1 vssd1 scanchain
Xscanchain_122 scanchain_122/clk_in scanchain_123/clk_in scanchain_122/data_in scanchain_123/data_in
+ scanchain_122/latch_enable_in scanchain_123/latch_enable_in scanchain_122/module_data_in[0]
+ scanchain_122/module_data_in[1] scanchain_122/module_data_in[2] scanchain_122/module_data_in[3]
+ scanchain_122/module_data_in[4] scanchain_122/module_data_in[5] scanchain_122/module_data_in[6]
+ scanchain_122/module_data_in[7] scanchain_122/module_data_out[0] scanchain_122/module_data_out[1]
+ scanchain_122/module_data_out[2] scanchain_122/module_data_out[3] scanchain_122/module_data_out[4]
+ scanchain_122/module_data_out[5] scanchain_122/module_data_out[6] scanchain_122/module_data_out[7]
+ scanchain_122/scan_select_in scanchain_123/scan_select_in vccd1 vssd1 scanchain
Xscanchain_144 scanchain_144/clk_in scanchain_145/clk_in scanchain_144/data_in scanchain_145/data_in
+ scanchain_144/latch_enable_in scanchain_145/latch_enable_in scanchain_144/module_data_in[0]
+ scanchain_144/module_data_in[1] scanchain_144/module_data_in[2] scanchain_144/module_data_in[3]
+ scanchain_144/module_data_in[4] scanchain_144/module_data_in[5] scanchain_144/module_data_in[6]
+ scanchain_144/module_data_in[7] scanchain_144/module_data_out[0] scanchain_144/module_data_out[1]
+ scanchain_144/module_data_out[2] scanchain_144/module_data_out[3] scanchain_144/module_data_out[4]
+ scanchain_144/module_data_out[5] scanchain_144/module_data_out[6] scanchain_144/module_data_out[7]
+ scanchain_144/scan_select_in scanchain_145/scan_select_in vccd1 vssd1 scanchain
Xscanchain_133 scanchain_133/clk_in scanchain_134/clk_in scanchain_133/data_in scanchain_134/data_in
+ scanchain_133/latch_enable_in scanchain_134/latch_enable_in scanchain_133/module_data_in[0]
+ scanchain_133/module_data_in[1] scanchain_133/module_data_in[2] scanchain_133/module_data_in[3]
+ scanchain_133/module_data_in[4] scanchain_133/module_data_in[5] scanchain_133/module_data_in[6]
+ scanchain_133/module_data_in[7] scanchain_133/module_data_out[0] scanchain_133/module_data_out[1]
+ scanchain_133/module_data_out[2] scanchain_133/module_data_out[3] scanchain_133/module_data_out[4]
+ scanchain_133/module_data_out[5] scanchain_133/module_data_out[6] scanchain_133/module_data_out[7]
+ scanchain_133/scan_select_in scanchain_134/scan_select_in vccd1 vssd1 scanchain
Xscanchain_155 scanchain_155/clk_in scanchain_156/clk_in scanchain_155/data_in scanchain_156/data_in
+ scanchain_155/latch_enable_in scanchain_156/latch_enable_in scanchain_155/module_data_in[0]
+ scanchain_155/module_data_in[1] scanchain_155/module_data_in[2] scanchain_155/module_data_in[3]
+ scanchain_155/module_data_in[4] scanchain_155/module_data_in[5] scanchain_155/module_data_in[6]
+ scanchain_155/module_data_in[7] scanchain_155/module_data_out[0] scanchain_155/module_data_out[1]
+ scanchain_155/module_data_out[2] scanchain_155/module_data_out[3] scanchain_155/module_data_out[4]
+ scanchain_155/module_data_out[5] scanchain_155/module_data_out[6] scanchain_155/module_data_out[7]
+ scanchain_155/scan_select_in scanchain_156/scan_select_in vccd1 vssd1 scanchain
Xscanchain_166 scanchain_166/clk_in scanchain_167/clk_in scanchain_166/data_in scanchain_167/data_in
+ scanchain_166/latch_enable_in scanchain_167/latch_enable_in scanchain_166/module_data_in[0]
+ scanchain_166/module_data_in[1] scanchain_166/module_data_in[2] scanchain_166/module_data_in[3]
+ scanchain_166/module_data_in[4] scanchain_166/module_data_in[5] scanchain_166/module_data_in[6]
+ scanchain_166/module_data_in[7] scanchain_166/module_data_out[0] scanchain_166/module_data_out[1]
+ scanchain_166/module_data_out[2] scanchain_166/module_data_out[3] scanchain_166/module_data_out[4]
+ scanchain_166/module_data_out[5] scanchain_166/module_data_out[6] scanchain_166/module_data_out[7]
+ scanchain_166/scan_select_in scanchain_167/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_180 scanchain_180/module_data_in[0] scanchain_180/module_data_in[1]
+ scanchain_180/module_data_in[2] scanchain_180/module_data_in[3] scanchain_180/module_data_in[4]
+ scanchain_180/module_data_in[5] scanchain_180/module_data_in[6] scanchain_180/module_data_in[7]
+ scanchain_180/module_data_out[0] scanchain_180/module_data_out[1] scanchain_180/module_data_out[2]
+ scanchain_180/module_data_out[3] scanchain_180/module_data_out[4] scanchain_180/module_data_out[5]
+ scanchain_180/module_data_out[6] scanchain_180/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_199 scanchain_199/clk_in scanchain_200/clk_in scanchain_199/data_in scanchain_200/data_in
+ scanchain_199/latch_enable_in scanchain_200/latch_enable_in scanchain_199/module_data_in[0]
+ scanchain_199/module_data_in[1] scanchain_199/module_data_in[2] scanchain_199/module_data_in[3]
+ scanchain_199/module_data_in[4] scanchain_199/module_data_in[5] scanchain_199/module_data_in[6]
+ scanchain_199/module_data_in[7] scanchain_199/module_data_out[0] scanchain_199/module_data_out[1]
+ scanchain_199/module_data_out[2] scanchain_199/module_data_out[3] scanchain_199/module_data_out[4]
+ scanchain_199/module_data_out[5] scanchain_199/module_data_out[6] scanchain_199/module_data_out[7]
+ scanchain_199/scan_select_in scanchain_200/scan_select_in vccd1 vssd1 scanchain
Xyubex_egg_timer_29 yubex_egg_timer_29/io_in[0] yubex_egg_timer_29/io_in[1] yubex_egg_timer_29/io_in[2]
+ yubex_egg_timer_29/io_in[3] yubex_egg_timer_29/io_in[4] yubex_egg_timer_29/io_in[5]
+ yubex_egg_timer_29/io_in[6] yubex_egg_timer_29/io_in[7] yubex_egg_timer_29/io_out[0]
+ yubex_egg_timer_29/io_out[1] yubex_egg_timer_29/io_out[2] yubex_egg_timer_29/io_out[3]
+ yubex_egg_timer_29/io_out[4] yubex_egg_timer_29/io_out[5] yubex_egg_timer_29/io_out[6]
+ yubex_egg_timer_29/io_out[7] vccd1 vssd1 yubex_egg_timer
Xuser_module_347619669052490324_56 scanchain_56/module_data_in[0] scanchain_56/module_data_in[1]
+ scanchain_56/module_data_in[2] scanchain_56/module_data_in[3] scanchain_56/module_data_in[4]
+ scanchain_56/module_data_in[5] scanchain_56/module_data_in[6] scanchain_56/module_data_in[7]
+ scanchain_56/module_data_out[0] scanchain_56/module_data_out[1] scanchain_56/module_data_out[2]
+ scanchain_56/module_data_out[3] scanchain_56/module_data_out[4] scanchain_56/module_data_out[5]
+ scanchain_56/module_data_out[6] scanchain_56/module_data_out[7] vccd1 vssd1 user_module_347619669052490324
Xscanchain_177 scanchain_177/clk_in scanchain_178/clk_in scanchain_177/data_in scanchain_178/data_in
+ scanchain_177/latch_enable_in scanchain_178/latch_enable_in scanchain_177/module_data_in[0]
+ scanchain_177/module_data_in[1] scanchain_177/module_data_in[2] scanchain_177/module_data_in[3]
+ scanchain_177/module_data_in[4] scanchain_177/module_data_in[5] scanchain_177/module_data_in[6]
+ scanchain_177/module_data_in[7] scanchain_177/module_data_out[0] scanchain_177/module_data_out[1]
+ scanchain_177/module_data_out[2] scanchain_177/module_data_out[3] scanchain_177/module_data_out[4]
+ scanchain_177/module_data_out[5] scanchain_177/module_data_out[6] scanchain_177/module_data_out[7]
+ scanchain_177/scan_select_in scanchain_178/scan_select_in vccd1 vssd1 scanchain
Xscanchain_188 scanchain_188/clk_in scanchain_189/clk_in scanchain_188/data_in scanchain_189/data_in
+ scanchain_188/latch_enable_in scanchain_189/latch_enable_in scanchain_188/module_data_in[0]
+ scanchain_188/module_data_in[1] scanchain_188/module_data_in[2] scanchain_188/module_data_in[3]
+ scanchain_188/module_data_in[4] scanchain_188/module_data_in[5] scanchain_188/module_data_in[6]
+ scanchain_188/module_data_in[7] scanchain_188/module_data_out[0] scanchain_188/module_data_out[1]
+ scanchain_188/module_data_out[2] scanchain_188/module_data_out[3] scanchain_188/module_data_out[4]
+ scanchain_188/module_data_out[5] scanchain_188/module_data_out[6] scanchain_188/module_data_out[7]
+ scanchain_188/scan_select_in scanchain_189/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_395 scanchain_395/module_data_in[0] scanchain_395/module_data_in[1]
+ scanchain_395/module_data_in[2] scanchain_395/module_data_in[3] scanchain_395/module_data_in[4]
+ scanchain_395/module_data_in[5] scanchain_395/module_data_in[6] scanchain_395/module_data_in[7]
+ scanchain_395/module_data_out[0] scanchain_395/module_data_out[1] scanchain_395/module_data_out[2]
+ scanchain_395/module_data_out[3] scanchain_395/module_data_out[4] scanchain_395/module_data_out[5]
+ scanchain_395/module_data_out[6] scanchain_395/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_384 scanchain_384/module_data_in[0] scanchain_384/module_data_in[1]
+ scanchain_384/module_data_in[2] scanchain_384/module_data_in[3] scanchain_384/module_data_in[4]
+ scanchain_384/module_data_in[5] scanchain_384/module_data_in[6] scanchain_384/module_data_in[7]
+ scanchain_384/module_data_out[0] scanchain_384/module_data_out[1] scanchain_384/module_data_out[2]
+ scanchain_384/module_data_out[3] scanchain_384/module_data_out[4] scanchain_384/module_data_out[5]
+ scanchain_384/module_data_out[6] scanchain_384/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_359 scanchain_359/clk_in scanchain_360/clk_in scanchain_359/data_in scanchain_360/data_in
+ scanchain_359/latch_enable_in scanchain_360/latch_enable_in scanchain_359/module_data_in[0]
+ scanchain_359/module_data_in[1] scanchain_359/module_data_in[2] scanchain_359/module_data_in[3]
+ scanchain_359/module_data_in[4] scanchain_359/module_data_in[5] scanchain_359/module_data_in[6]
+ scanchain_359/module_data_in[7] scanchain_359/module_data_out[0] scanchain_359/module_data_out[1]
+ scanchain_359/module_data_out[2] scanchain_359/module_data_out[3] scanchain_359/module_data_out[4]
+ scanchain_359/module_data_out[5] scanchain_359/module_data_out[6] scanchain_359/module_data_out[7]
+ scanchain_359/scan_select_in scanchain_360/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_362 scanchain_362/module_data_in[0] scanchain_362/module_data_in[1]
+ scanchain_362/module_data_in[2] scanchain_362/module_data_in[3] scanchain_362/module_data_in[4]
+ scanchain_362/module_data_in[5] scanchain_362/module_data_in[6] scanchain_362/module_data_in[7]
+ scanchain_362/module_data_out[0] scanchain_362/module_data_out[1] scanchain_362/module_data_out[2]
+ scanchain_362/module_data_out[3] scanchain_362/module_data_out[4] scanchain_362/module_data_out[5]
+ scanchain_362/module_data_out[6] scanchain_362/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_373 scanchain_373/module_data_in[0] scanchain_373/module_data_in[1]
+ scanchain_373/module_data_in[2] scanchain_373/module_data_in[3] scanchain_373/module_data_in[4]
+ scanchain_373/module_data_in[5] scanchain_373/module_data_in[6] scanchain_373/module_data_in[7]
+ scanchain_373/module_data_out[0] scanchain_373/module_data_out[1] scanchain_373/module_data_out[2]
+ scanchain_373/module_data_out[3] scanchain_373/module_data_out[4] scanchain_373/module_data_out[5]
+ scanchain_373/module_data_out[6] scanchain_373/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_351 scanchain_351/module_data_in[0] scanchain_351/module_data_in[1]
+ scanchain_351/module_data_in[2] scanchain_351/module_data_in[3] scanchain_351/module_data_in[4]
+ scanchain_351/module_data_in[5] scanchain_351/module_data_in[6] scanchain_351/module_data_in[7]
+ scanchain_351/module_data_out[0] scanchain_351/module_data_out[1] scanchain_351/module_data_out[2]
+ scanchain_351/module_data_out[3] scanchain_351/module_data_out[4] scanchain_351/module_data_out[5]
+ scanchain_351/module_data_out[6] scanchain_351/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_348 scanchain_348/clk_in scanchain_349/clk_in scanchain_348/data_in scanchain_349/data_in
+ scanchain_348/latch_enable_in scanchain_349/latch_enable_in scanchain_348/module_data_in[0]
+ scanchain_348/module_data_in[1] scanchain_348/module_data_in[2] scanchain_348/module_data_in[3]
+ scanchain_348/module_data_in[4] scanchain_348/module_data_in[5] scanchain_348/module_data_in[6]
+ scanchain_348/module_data_in[7] scanchain_348/module_data_out[0] scanchain_348/module_data_out[1]
+ scanchain_348/module_data_out[2] scanchain_348/module_data_out[3] scanchain_348/module_data_out[4]
+ scanchain_348/module_data_out[5] scanchain_348/module_data_out[6] scanchain_348/module_data_out[7]
+ scanchain_348/scan_select_in scanchain_349/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_340 scanchain_340/module_data_in[0] scanchain_340/module_data_in[1]
+ scanchain_340/module_data_in[2] scanchain_340/module_data_in[3] scanchain_340/module_data_in[4]
+ scanchain_340/module_data_in[5] scanchain_340/module_data_in[6] scanchain_340/module_data_in[7]
+ scanchain_340/module_data_out[0] scanchain_340/module_data_out[1] scanchain_340/module_data_out[2]
+ scanchain_340/module_data_out[3] scanchain_340/module_data_out[4] scanchain_340/module_data_out[5]
+ scanchain_340/module_data_out[6] scanchain_340/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_326 scanchain_326/clk_in scanchain_327/clk_in scanchain_326/data_in scanchain_327/data_in
+ scanchain_326/latch_enable_in scanchain_327/latch_enable_in scanchain_326/module_data_in[0]
+ scanchain_326/module_data_in[1] scanchain_326/module_data_in[2] scanchain_326/module_data_in[3]
+ scanchain_326/module_data_in[4] scanchain_326/module_data_in[5] scanchain_326/module_data_in[6]
+ scanchain_326/module_data_in[7] scanchain_326/module_data_out[0] scanchain_326/module_data_out[1]
+ scanchain_326/module_data_out[2] scanchain_326/module_data_out[3] scanchain_326/module_data_out[4]
+ scanchain_326/module_data_out[5] scanchain_326/module_data_out[6] scanchain_326/module_data_out[7]
+ scanchain_326/scan_select_in scanchain_327/scan_select_in vccd1 vssd1 scanchain
Xscanchain_337 scanchain_337/clk_in scanchain_338/clk_in scanchain_337/data_in scanchain_338/data_in
+ scanchain_337/latch_enable_in scanchain_338/latch_enable_in scanchain_337/module_data_in[0]
+ scanchain_337/module_data_in[1] scanchain_337/module_data_in[2] scanchain_337/module_data_in[3]
+ scanchain_337/module_data_in[4] scanchain_337/module_data_in[5] scanchain_337/module_data_in[6]
+ scanchain_337/module_data_in[7] scanchain_337/module_data_out[0] scanchain_337/module_data_out[1]
+ scanchain_337/module_data_out[2] scanchain_337/module_data_out[3] scanchain_337/module_data_out[4]
+ scanchain_337/module_data_out[5] scanchain_337/module_data_out[6] scanchain_337/module_data_out[7]
+ scanchain_337/scan_select_in scanchain_338/scan_select_in vccd1 vssd1 scanchain
Xscanchain_315 scanchain_315/clk_in scanchain_316/clk_in scanchain_315/data_in scanchain_316/data_in
+ scanchain_315/latch_enable_in scanchain_316/latch_enable_in scanchain_315/module_data_in[0]
+ scanchain_315/module_data_in[1] scanchain_315/module_data_in[2] scanchain_315/module_data_in[3]
+ scanchain_315/module_data_in[4] scanchain_315/module_data_in[5] scanchain_315/module_data_in[6]
+ scanchain_315/module_data_in[7] scanchain_315/module_data_out[0] scanchain_315/module_data_out[1]
+ scanchain_315/module_data_out[2] scanchain_315/module_data_out[3] scanchain_315/module_data_out[4]
+ scanchain_315/module_data_out[5] scanchain_315/module_data_out[6] scanchain_315/module_data_out[7]
+ scanchain_315/scan_select_in scanchain_316/scan_select_in vccd1 vssd1 scanchain
Xscanchain_304 scanchain_304/clk_in scanchain_305/clk_in scanchain_304/data_in scanchain_305/data_in
+ scanchain_304/latch_enable_in scanchain_305/latch_enable_in scanchain_304/module_data_in[0]
+ scanchain_304/module_data_in[1] scanchain_304/module_data_in[2] scanchain_304/module_data_in[3]
+ scanchain_304/module_data_in[4] scanchain_304/module_data_in[5] scanchain_304/module_data_in[6]
+ scanchain_304/module_data_in[7] scanchain_304/module_data_out[0] scanchain_304/module_data_out[1]
+ scanchain_304/module_data_out[2] scanchain_304/module_data_out[3] scanchain_304/module_data_out[4]
+ scanchain_304/module_data_out[5] scanchain_304/module_data_out[6] scanchain_304/module_data_out[7]
+ scanchain_304/scan_select_in scanchain_305/scan_select_in vccd1 vssd1 scanchain
Xuser_module_348121131386929746_28 scanchain_28/module_data_in[0] scanchain_28/module_data_in[1]
+ scanchain_28/module_data_in[2] scanchain_28/module_data_in[3] scanchain_28/module_data_in[4]
+ scanchain_28/module_data_in[5] scanchain_28/module_data_in[6] scanchain_28/module_data_in[7]
+ scanchain_28/module_data_out[0] scanchain_28/module_data_out[1] scanchain_28/module_data_out[2]
+ scanchain_28/module_data_out[3] scanchain_28/module_data_out[4] scanchain_28/module_data_out[5]
+ scanchain_28/module_data_out[6] scanchain_28/module_data_out[7] vccd1 vssd1 user_module_348121131386929746
Xuser_module_339501025136214612_192 scanchain_192/module_data_in[0] scanchain_192/module_data_in[1]
+ scanchain_192/module_data_in[2] scanchain_192/module_data_in[3] scanchain_192/module_data_in[4]
+ scanchain_192/module_data_in[5] scanchain_192/module_data_in[6] scanchain_192/module_data_in[7]
+ scanchain_192/module_data_out[0] scanchain_192/module_data_out[1] scanchain_192/module_data_out[2]
+ scanchain_192/module_data_out[3] scanchain_192/module_data_out[4] scanchain_192/module_data_out[5]
+ scanchain_192/module_data_out[6] scanchain_192/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_181 scanchain_181/module_data_in[0] scanchain_181/module_data_in[1]
+ scanchain_181/module_data_in[2] scanchain_181/module_data_in[3] scanchain_181/module_data_in[4]
+ scanchain_181/module_data_in[5] scanchain_181/module_data_in[6] scanchain_181/module_data_in[7]
+ scanchain_181/module_data_out[0] scanchain_181/module_data_out[1] scanchain_181/module_data_out[2]
+ scanchain_181/module_data_out[3] scanchain_181/module_data_out[4] scanchain_181/module_data_out[5]
+ scanchain_181/module_data_out[6] scanchain_181/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_170 scanchain_170/module_data_in[0] scanchain_170/module_data_in[1]
+ scanchain_170/module_data_in[2] scanchain_170/module_data_in[3] scanchain_170/module_data_in[4]
+ scanchain_170/module_data_in[5] scanchain_170/module_data_in[6] scanchain_170/module_data_in[7]
+ scanchain_170/module_data_out[0] scanchain_170/module_data_out[1] scanchain_170/module_data_out[2]
+ scanchain_170/module_data_out[3] scanchain_170/module_data_out[4] scanchain_170/module_data_out[5]
+ scanchain_170/module_data_out[6] scanchain_170/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_101 scanchain_101/clk_in scanchain_102/clk_in scanchain_101/data_in scanchain_102/data_in
+ scanchain_101/latch_enable_in scanchain_102/latch_enable_in scanchain_101/module_data_in[0]
+ scanchain_101/module_data_in[1] scanchain_101/module_data_in[2] scanchain_101/module_data_in[3]
+ scanchain_101/module_data_in[4] scanchain_101/module_data_in[5] scanchain_101/module_data_in[6]
+ scanchain_101/module_data_in[7] scanchain_101/module_data_out[0] scanchain_101/module_data_out[1]
+ scanchain_101/module_data_out[2] scanchain_101/module_data_out[3] scanchain_101/module_data_out[4]
+ scanchain_101/module_data_out[5] scanchain_101/module_data_out[6] scanchain_101/module_data_out[7]
+ scanchain_101/scan_select_in scanchain_102/scan_select_in vccd1 vssd1 scanchain
Xscanchain_112 scanchain_112/clk_in scanchain_113/clk_in scanchain_112/data_in scanchain_113/data_in
+ scanchain_112/latch_enable_in scanchain_113/latch_enable_in scanchain_112/module_data_in[0]
+ scanchain_112/module_data_in[1] scanchain_112/module_data_in[2] scanchain_112/module_data_in[3]
+ scanchain_112/module_data_in[4] scanchain_112/module_data_in[5] scanchain_112/module_data_in[6]
+ scanchain_112/module_data_in[7] scanchain_112/module_data_out[0] scanchain_112/module_data_out[1]
+ scanchain_112/module_data_out[2] scanchain_112/module_data_out[3] scanchain_112/module_data_out[4]
+ scanchain_112/module_data_out[5] scanchain_112/module_data_out[6] scanchain_112/module_data_out[7]
+ scanchain_112/scan_select_in scanchain_113/scan_select_in vccd1 vssd1 scanchain
Xscanchain_123 scanchain_123/clk_in scanchain_124/clk_in scanchain_123/data_in scanchain_124/data_in
+ scanchain_123/latch_enable_in scanchain_124/latch_enable_in scanchain_123/module_data_in[0]
+ scanchain_123/module_data_in[1] scanchain_123/module_data_in[2] scanchain_123/module_data_in[3]
+ scanchain_123/module_data_in[4] scanchain_123/module_data_in[5] scanchain_123/module_data_in[6]
+ scanchain_123/module_data_in[7] scanchain_123/module_data_out[0] scanchain_123/module_data_out[1]
+ scanchain_123/module_data_out[2] scanchain_123/module_data_out[3] scanchain_123/module_data_out[4]
+ scanchain_123/module_data_out[5] scanchain_123/module_data_out[6] scanchain_123/module_data_out[7]
+ scanchain_123/scan_select_in scanchain_124/scan_select_in vccd1 vssd1 scanchain
Xscanchain_145 scanchain_145/clk_in scanchain_146/clk_in scanchain_145/data_in scanchain_146/data_in
+ scanchain_145/latch_enable_in scanchain_146/latch_enable_in scanchain_145/module_data_in[0]
+ scanchain_145/module_data_in[1] scanchain_145/module_data_in[2] scanchain_145/module_data_in[3]
+ scanchain_145/module_data_in[4] scanchain_145/module_data_in[5] scanchain_145/module_data_in[6]
+ scanchain_145/module_data_in[7] scanchain_145/module_data_out[0] scanchain_145/module_data_out[1]
+ scanchain_145/module_data_out[2] scanchain_145/module_data_out[3] scanchain_145/module_data_out[4]
+ scanchain_145/module_data_out[5] scanchain_145/module_data_out[6] scanchain_145/module_data_out[7]
+ scanchain_145/scan_select_in scanchain_146/scan_select_in vccd1 vssd1 scanchain
Xscanchain_134 scanchain_134/clk_in scanchain_135/clk_in scanchain_134/data_in scanchain_135/data_in
+ scanchain_134/latch_enable_in scanchain_135/latch_enable_in scanchain_134/module_data_in[0]
+ scanchain_134/module_data_in[1] scanchain_134/module_data_in[2] scanchain_134/module_data_in[3]
+ scanchain_134/module_data_in[4] scanchain_134/module_data_in[5] scanchain_134/module_data_in[6]
+ scanchain_134/module_data_in[7] scanchain_134/module_data_out[0] scanchain_134/module_data_out[1]
+ scanchain_134/module_data_out[2] scanchain_134/module_data_out[3] scanchain_134/module_data_out[4]
+ scanchain_134/module_data_out[5] scanchain_134/module_data_out[6] scanchain_134/module_data_out[7]
+ scanchain_134/scan_select_in scanchain_135/scan_select_in vccd1 vssd1 scanchain
Xscanchain_156 scanchain_156/clk_in scanchain_157/clk_in scanchain_156/data_in scanchain_157/data_in
+ scanchain_156/latch_enable_in scanchain_157/latch_enable_in scanchain_156/module_data_in[0]
+ scanchain_156/module_data_in[1] scanchain_156/module_data_in[2] scanchain_156/module_data_in[3]
+ scanchain_156/module_data_in[4] scanchain_156/module_data_in[5] scanchain_156/module_data_in[6]
+ scanchain_156/module_data_in[7] scanchain_156/module_data_out[0] scanchain_156/module_data_out[1]
+ scanchain_156/module_data_out[2] scanchain_156/module_data_out[3] scanchain_156/module_data_out[4]
+ scanchain_156/module_data_out[5] scanchain_156/module_data_out[6] scanchain_156/module_data_out[7]
+ scanchain_156/scan_select_in scanchain_157/scan_select_in vccd1 vssd1 scanchain
Xscanchain_167 scanchain_167/clk_in scanchain_168/clk_in scanchain_167/data_in scanchain_168/data_in
+ scanchain_167/latch_enable_in scanchain_168/latch_enable_in scanchain_167/module_data_in[0]
+ scanchain_167/module_data_in[1] scanchain_167/module_data_in[2] scanchain_167/module_data_in[3]
+ scanchain_167/module_data_in[4] scanchain_167/module_data_in[5] scanchain_167/module_data_in[6]
+ scanchain_167/module_data_in[7] scanchain_167/module_data_out[0] scanchain_167/module_data_out[1]
+ scanchain_167/module_data_out[2] scanchain_167/module_data_out[3] scanchain_167/module_data_out[4]
+ scanchain_167/module_data_out[5] scanchain_167/module_data_out[6] scanchain_167/module_data_out[7]
+ scanchain_167/scan_select_in scanchain_168/scan_select_in vccd1 vssd1 scanchain
Xscanchain_178 scanchain_178/clk_in scanchain_179/clk_in scanchain_178/data_in scanchain_179/data_in
+ scanchain_178/latch_enable_in scanchain_179/latch_enable_in scanchain_178/module_data_in[0]
+ scanchain_178/module_data_in[1] scanchain_178/module_data_in[2] scanchain_178/module_data_in[3]
+ scanchain_178/module_data_in[4] scanchain_178/module_data_in[5] scanchain_178/module_data_in[6]
+ scanchain_178/module_data_in[7] scanchain_178/module_data_out[0] scanchain_178/module_data_out[1]
+ scanchain_178/module_data_out[2] scanchain_178/module_data_out[3] scanchain_178/module_data_out[4]
+ scanchain_178/module_data_out[5] scanchain_178/module_data_out[6] scanchain_178/module_data_out[7]
+ scanchain_178/scan_select_in scanchain_179/scan_select_in vccd1 vssd1 scanchain
Xscanchain_189 scanchain_189/clk_in scanchain_190/clk_in scanchain_189/data_in scanchain_190/data_in
+ scanchain_189/latch_enable_in scanchain_190/latch_enable_in scanchain_189/module_data_in[0]
+ scanchain_189/module_data_in[1] scanchain_189/module_data_in[2] scanchain_189/module_data_in[3]
+ scanchain_189/module_data_in[4] scanchain_189/module_data_in[5] scanchain_189/module_data_in[6]
+ scanchain_189/module_data_in[7] scanchain_189/module_data_out[0] scanchain_189/module_data_out[1]
+ scanchain_189/module_data_out[2] scanchain_189/module_data_out[3] scanchain_189/module_data_out[4]
+ scanchain_189/module_data_out[5] scanchain_189/module_data_out[6] scanchain_189/module_data_out[7]
+ scanchain_189/scan_select_in scanchain_190/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_396 scanchain_396/module_data_in[0] scanchain_396/module_data_in[1]
+ scanchain_396/module_data_in[2] scanchain_396/module_data_in[3] scanchain_396/module_data_in[4]
+ scanchain_396/module_data_in[5] scanchain_396/module_data_in[6] scanchain_396/module_data_in[7]
+ scanchain_396/module_data_out[0] scanchain_396/module_data_out[1] scanchain_396/module_data_out[2]
+ scanchain_396/module_data_out[3] scanchain_396/module_data_out[4] scanchain_396/module_data_out[5]
+ scanchain_396/module_data_out[6] scanchain_396/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_385 scanchain_385/module_data_in[0] scanchain_385/module_data_in[1]
+ scanchain_385/module_data_in[2] scanchain_385/module_data_in[3] scanchain_385/module_data_in[4]
+ scanchain_385/module_data_in[5] scanchain_385/module_data_in[6] scanchain_385/module_data_in[7]
+ scanchain_385/module_data_out[0] scanchain_385/module_data_out[1] scanchain_385/module_data_out[2]
+ scanchain_385/module_data_out[3] scanchain_385/module_data_out[4] scanchain_385/module_data_out[5]
+ scanchain_385/module_data_out[6] scanchain_385/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_363 scanchain_363/module_data_in[0] scanchain_363/module_data_in[1]
+ scanchain_363/module_data_in[2] scanchain_363/module_data_in[3] scanchain_363/module_data_in[4]
+ scanchain_363/module_data_in[5] scanchain_363/module_data_in[6] scanchain_363/module_data_in[7]
+ scanchain_363/module_data_out[0] scanchain_363/module_data_out[1] scanchain_363/module_data_out[2]
+ scanchain_363/module_data_out[3] scanchain_363/module_data_out[4] scanchain_363/module_data_out[5]
+ scanchain_363/module_data_out[6] scanchain_363/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_374 scanchain_374/module_data_in[0] scanchain_374/module_data_in[1]
+ scanchain_374/module_data_in[2] scanchain_374/module_data_in[3] scanchain_374/module_data_in[4]
+ scanchain_374/module_data_in[5] scanchain_374/module_data_in[6] scanchain_374/module_data_in[7]
+ scanchain_374/module_data_out[0] scanchain_374/module_data_out[1] scanchain_374/module_data_out[2]
+ scanchain_374/module_data_out[3] scanchain_374/module_data_out[4] scanchain_374/module_data_out[5]
+ scanchain_374/module_data_out[6] scanchain_374/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_352 scanchain_352/module_data_in[0] scanchain_352/module_data_in[1]
+ scanchain_352/module_data_in[2] scanchain_352/module_data_in[3] scanchain_352/module_data_in[4]
+ scanchain_352/module_data_in[5] scanchain_352/module_data_in[6] scanchain_352/module_data_in[7]
+ scanchain_352/module_data_out[0] scanchain_352/module_data_out[1] scanchain_352/module_data_out[2]
+ scanchain_352/module_data_out[3] scanchain_352/module_data_out[4] scanchain_352/module_data_out[5]
+ scanchain_352/module_data_out[6] scanchain_352/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_349 scanchain_349/clk_in scanchain_350/clk_in scanchain_349/data_in scanchain_350/data_in
+ scanchain_349/latch_enable_in scanchain_350/latch_enable_in scanchain_349/module_data_in[0]
+ scanchain_349/module_data_in[1] scanchain_349/module_data_in[2] scanchain_349/module_data_in[3]
+ scanchain_349/module_data_in[4] scanchain_349/module_data_in[5] scanchain_349/module_data_in[6]
+ scanchain_349/module_data_in[7] scanchain_349/module_data_out[0] scanchain_349/module_data_out[1]
+ scanchain_349/module_data_out[2] scanchain_349/module_data_out[3] scanchain_349/module_data_out[4]
+ scanchain_349/module_data_out[5] scanchain_349/module_data_out[6] scanchain_349/module_data_out[7]
+ scanchain_349/scan_select_in scanchain_350/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_341 scanchain_341/module_data_in[0] scanchain_341/module_data_in[1]
+ scanchain_341/module_data_in[2] scanchain_341/module_data_in[3] scanchain_341/module_data_in[4]
+ scanchain_341/module_data_in[5] scanchain_341/module_data_in[6] scanchain_341/module_data_in[7]
+ scanchain_341/module_data_out[0] scanchain_341/module_data_out[1] scanchain_341/module_data_out[2]
+ scanchain_341/module_data_out[3] scanchain_341/module_data_out[4] scanchain_341/module_data_out[5]
+ scanchain_341/module_data_out[6] scanchain_341/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_327 scanchain_327/clk_in scanchain_328/clk_in scanchain_327/data_in scanchain_328/data_in
+ scanchain_327/latch_enable_in scanchain_328/latch_enable_in scanchain_327/module_data_in[0]
+ scanchain_327/module_data_in[1] scanchain_327/module_data_in[2] scanchain_327/module_data_in[3]
+ scanchain_327/module_data_in[4] scanchain_327/module_data_in[5] scanchain_327/module_data_in[6]
+ scanchain_327/module_data_in[7] scanchain_327/module_data_out[0] scanchain_327/module_data_out[1]
+ scanchain_327/module_data_out[2] scanchain_327/module_data_out[3] scanchain_327/module_data_out[4]
+ scanchain_327/module_data_out[5] scanchain_327/module_data_out[6] scanchain_327/module_data_out[7]
+ scanchain_327/scan_select_in scanchain_328/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_330 scanchain_330/module_data_in[0] scanchain_330/module_data_in[1]
+ scanchain_330/module_data_in[2] scanchain_330/module_data_in[3] scanchain_330/module_data_in[4]
+ scanchain_330/module_data_in[5] scanchain_330/module_data_in[6] scanchain_330/module_data_in[7]
+ scanchain_330/module_data_out[0] scanchain_330/module_data_out[1] scanchain_330/module_data_out[2]
+ scanchain_330/module_data_out[3] scanchain_330/module_data_out[4] scanchain_330/module_data_out[5]
+ scanchain_330/module_data_out[6] scanchain_330/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_338 scanchain_338/clk_in scanchain_339/clk_in scanchain_338/data_in scanchain_339/data_in
+ scanchain_338/latch_enable_in scanchain_339/latch_enable_in scanchain_338/module_data_in[0]
+ scanchain_338/module_data_in[1] scanchain_338/module_data_in[2] scanchain_338/module_data_in[3]
+ scanchain_338/module_data_in[4] scanchain_338/module_data_in[5] scanchain_338/module_data_in[6]
+ scanchain_338/module_data_in[7] scanchain_338/module_data_out[0] scanchain_338/module_data_out[1]
+ scanchain_338/module_data_out[2] scanchain_338/module_data_out[3] scanchain_338/module_data_out[4]
+ scanchain_338/module_data_out[5] scanchain_338/module_data_out[6] scanchain_338/module_data_out[7]
+ scanchain_338/scan_select_in scanchain_339/scan_select_in vccd1 vssd1 scanchain
Xscanchain_316 scanchain_316/clk_in scanchain_317/clk_in scanchain_316/data_in scanchain_317/data_in
+ scanchain_316/latch_enable_in scanchain_317/latch_enable_in scanchain_316/module_data_in[0]
+ scanchain_316/module_data_in[1] scanchain_316/module_data_in[2] scanchain_316/module_data_in[3]
+ scanchain_316/module_data_in[4] scanchain_316/module_data_in[5] scanchain_316/module_data_in[6]
+ scanchain_316/module_data_in[7] scanchain_316/module_data_out[0] scanchain_316/module_data_out[1]
+ scanchain_316/module_data_out[2] scanchain_316/module_data_out[3] scanchain_316/module_data_out[4]
+ scanchain_316/module_data_out[5] scanchain_316/module_data_out[6] scanchain_316/module_data_out[7]
+ scanchain_316/scan_select_in scanchain_317/scan_select_in vccd1 vssd1 scanchain
Xscanchain_305 scanchain_305/clk_in scanchain_306/clk_in scanchain_305/data_in scanchain_306/data_in
+ scanchain_305/latch_enable_in scanchain_306/latch_enable_in scanchain_305/module_data_in[0]
+ scanchain_305/module_data_in[1] scanchain_305/module_data_in[2] scanchain_305/module_data_in[3]
+ scanchain_305/module_data_in[4] scanchain_305/module_data_in[5] scanchain_305/module_data_in[6]
+ scanchain_305/module_data_in[7] scanchain_305/module_data_out[0] scanchain_305/module_data_out[1]
+ scanchain_305/module_data_out[2] scanchain_305/module_data_out[3] scanchain_305/module_data_out[4]
+ scanchain_305/module_data_out[5] scanchain_305/module_data_out[6] scanchain_305/module_data_out[7]
+ scanchain_305/scan_select_in scanchain_306/scan_select_in vccd1 vssd1 scanchain
Xtt2_tholin_multiplexed_counter_50 scanchain_50/module_data_in[0] scanchain_50/module_data_in[1]
+ scanchain_50/module_data_in[2] scanchain_50/module_data_in[3] scanchain_50/module_data_in[4]
+ scanchain_50/module_data_in[5] scanchain_50/module_data_in[6] scanchain_50/module_data_in[7]
+ scanchain_50/module_data_out[0] scanchain_50/module_data_out[1] scanchain_50/module_data_out[2]
+ scanchain_50/module_data_out[3] scanchain_50/module_data_out[4] scanchain_50/module_data_out[5]
+ scanchain_50/module_data_out[6] scanchain_50/module_data_out[7] vccd1 vssd1 tt2_tholin_multiplexed_counter
Xuser_module_339501025136214612_193 scanchain_193/module_data_in[0] scanchain_193/module_data_in[1]
+ scanchain_193/module_data_in[2] scanchain_193/module_data_in[3] scanchain_193/module_data_in[4]
+ scanchain_193/module_data_in[5] scanchain_193/module_data_in[6] scanchain_193/module_data_in[7]
+ scanchain_193/module_data_out[0] scanchain_193/module_data_out[1] scanchain_193/module_data_out[2]
+ scanchain_193/module_data_out[3] scanchain_193/module_data_out[4] scanchain_193/module_data_out[5]
+ scanchain_193/module_data_out[6] scanchain_193/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_160 scanchain_160/module_data_in[0] scanchain_160/module_data_in[1]
+ scanchain_160/module_data_in[2] scanchain_160/module_data_in[3] scanchain_160/module_data_in[4]
+ scanchain_160/module_data_in[5] scanchain_160/module_data_in[6] scanchain_160/module_data_in[7]
+ scanchain_160/module_data_out[0] scanchain_160/module_data_out[1] scanchain_160/module_data_out[2]
+ scanchain_160/module_data_out[3] scanchain_160/module_data_out[4] scanchain_160/module_data_out[5]
+ scanchain_160/module_data_out[6] scanchain_160/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_182 scanchain_182/module_data_in[0] scanchain_182/module_data_in[1]
+ scanchain_182/module_data_in[2] scanchain_182/module_data_in[3] scanchain_182/module_data_in[4]
+ scanchain_182/module_data_in[5] scanchain_182/module_data_in[6] scanchain_182/module_data_in[7]
+ scanchain_182/module_data_out[0] scanchain_182/module_data_out[1] scanchain_182/module_data_out[2]
+ scanchain_182/module_data_out[3] scanchain_182/module_data_out[4] scanchain_182/module_data_out[5]
+ scanchain_182/module_data_out[6] scanchain_182/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_171 scanchain_171/module_data_in[0] scanchain_171/module_data_in[1]
+ scanchain_171/module_data_in[2] scanchain_171/module_data_in[3] scanchain_171/module_data_in[4]
+ scanchain_171/module_data_in[5] scanchain_171/module_data_in[6] scanchain_171/module_data_in[7]
+ scanchain_171/module_data_out[0] scanchain_171/module_data_out[1] scanchain_171/module_data_out[2]
+ scanchain_171/module_data_out[3] scanchain_171/module_data_out[4] scanchain_171/module_data_out[5]
+ scanchain_171/module_data_out[6] scanchain_171/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_102 scanchain_102/clk_in scanchain_103/clk_in scanchain_102/data_in scanchain_103/data_in
+ scanchain_102/latch_enable_in scanchain_103/latch_enable_in scanchain_102/module_data_in[0]
+ scanchain_102/module_data_in[1] scanchain_102/module_data_in[2] scanchain_102/module_data_in[3]
+ scanchain_102/module_data_in[4] scanchain_102/module_data_in[5] scanchain_102/module_data_in[6]
+ scanchain_102/module_data_in[7] scanchain_102/module_data_out[0] scanchain_102/module_data_out[1]
+ scanchain_102/module_data_out[2] scanchain_102/module_data_out[3] scanchain_102/module_data_out[4]
+ scanchain_102/module_data_out[5] scanchain_102/module_data_out[6] scanchain_102/module_data_out[7]
+ scanchain_102/scan_select_in scanchain_103/scan_select_in vccd1 vssd1 scanchain
Xscanchain_113 scanchain_113/clk_in scanchain_114/clk_in scanchain_113/data_in scanchain_114/data_in
+ scanchain_113/latch_enable_in scanchain_114/latch_enable_in scanchain_113/module_data_in[0]
+ scanchain_113/module_data_in[1] scanchain_113/module_data_in[2] scanchain_113/module_data_in[3]
+ scanchain_113/module_data_in[4] scanchain_113/module_data_in[5] scanchain_113/module_data_in[6]
+ scanchain_113/module_data_in[7] scanchain_113/module_data_out[0] scanchain_113/module_data_out[1]
+ scanchain_113/module_data_out[2] scanchain_113/module_data_out[3] scanchain_113/module_data_out[4]
+ scanchain_113/module_data_out[5] scanchain_113/module_data_out[6] scanchain_113/module_data_out[7]
+ scanchain_113/scan_select_in scanchain_114/scan_select_in vccd1 vssd1 scanchain
Xscanchain_124 scanchain_124/clk_in scanchain_125/clk_in scanchain_124/data_in scanchain_125/data_in
+ scanchain_124/latch_enable_in scanchain_125/latch_enable_in scanchain_124/module_data_in[0]
+ scanchain_124/module_data_in[1] scanchain_124/module_data_in[2] scanchain_124/module_data_in[3]
+ scanchain_124/module_data_in[4] scanchain_124/module_data_in[5] scanchain_124/module_data_in[6]
+ scanchain_124/module_data_in[7] scanchain_124/module_data_out[0] scanchain_124/module_data_out[1]
+ scanchain_124/module_data_out[2] scanchain_124/module_data_out[3] scanchain_124/module_data_out[4]
+ scanchain_124/module_data_out[5] scanchain_124/module_data_out[6] scanchain_124/module_data_out[7]
+ scanchain_124/scan_select_in scanchain_125/scan_select_in vccd1 vssd1 scanchain
Xscanchain_146 scanchain_146/clk_in scanchain_147/clk_in scanchain_146/data_in scanchain_147/data_in
+ scanchain_146/latch_enable_in scanchain_147/latch_enable_in scanchain_146/module_data_in[0]
+ scanchain_146/module_data_in[1] scanchain_146/module_data_in[2] scanchain_146/module_data_in[3]
+ scanchain_146/module_data_in[4] scanchain_146/module_data_in[5] scanchain_146/module_data_in[6]
+ scanchain_146/module_data_in[7] scanchain_146/module_data_out[0] scanchain_146/module_data_out[1]
+ scanchain_146/module_data_out[2] scanchain_146/module_data_out[3] scanchain_146/module_data_out[4]
+ scanchain_146/module_data_out[5] scanchain_146/module_data_out[6] scanchain_146/module_data_out[7]
+ scanchain_146/scan_select_in scanchain_147/scan_select_in vccd1 vssd1 scanchain
Xscanchain_135 scanchain_135/clk_in scanchain_136/clk_in scanchain_135/data_in scanchain_136/data_in
+ scanchain_135/latch_enable_in scanchain_136/latch_enable_in scanchain_135/module_data_in[0]
+ scanchain_135/module_data_in[1] scanchain_135/module_data_in[2] scanchain_135/module_data_in[3]
+ scanchain_135/module_data_in[4] scanchain_135/module_data_in[5] scanchain_135/module_data_in[6]
+ scanchain_135/module_data_in[7] scanchain_135/module_data_out[0] scanchain_135/module_data_out[1]
+ scanchain_135/module_data_out[2] scanchain_135/module_data_out[3] scanchain_135/module_data_out[4]
+ scanchain_135/module_data_out[5] scanchain_135/module_data_out[6] scanchain_135/module_data_out[7]
+ scanchain_135/scan_select_in scanchain_136/scan_select_in vccd1 vssd1 scanchain
Xscanchain_157 scanchain_157/clk_in scanchain_158/clk_in scanchain_157/data_in scanchain_158/data_in
+ scanchain_157/latch_enable_in scanchain_158/latch_enable_in scanchain_157/module_data_in[0]
+ scanchain_157/module_data_in[1] scanchain_157/module_data_in[2] scanchain_157/module_data_in[3]
+ scanchain_157/module_data_in[4] scanchain_157/module_data_in[5] scanchain_157/module_data_in[6]
+ scanchain_157/module_data_in[7] scanchain_157/module_data_out[0] scanchain_157/module_data_out[1]
+ scanchain_157/module_data_out[2] scanchain_157/module_data_out[3] scanchain_157/module_data_out[4]
+ scanchain_157/module_data_out[5] scanchain_157/module_data_out[6] scanchain_157/module_data_out[7]
+ scanchain_157/scan_select_in scanchain_158/scan_select_in vccd1 vssd1 scanchain
Xscanchain_168 scanchain_168/clk_in scanchain_169/clk_in scanchain_168/data_in scanchain_169/data_in
+ scanchain_168/latch_enable_in scanchain_169/latch_enable_in scanchain_168/module_data_in[0]
+ scanchain_168/module_data_in[1] scanchain_168/module_data_in[2] scanchain_168/module_data_in[3]
+ scanchain_168/module_data_in[4] scanchain_168/module_data_in[5] scanchain_168/module_data_in[6]
+ scanchain_168/module_data_in[7] scanchain_168/module_data_out[0] scanchain_168/module_data_out[1]
+ scanchain_168/module_data_out[2] scanchain_168/module_data_out[3] scanchain_168/module_data_out[4]
+ scanchain_168/module_data_out[5] scanchain_168/module_data_out[6] scanchain_168/module_data_out[7]
+ scanchain_168/scan_select_in scanchain_169/scan_select_in vccd1 vssd1 scanchain
Xscanchain_179 scanchain_179/clk_in scanchain_180/clk_in scanchain_179/data_in scanchain_180/data_in
+ scanchain_179/latch_enable_in scanchain_180/latch_enable_in scanchain_179/module_data_in[0]
+ scanchain_179/module_data_in[1] scanchain_179/module_data_in[2] scanchain_179/module_data_in[3]
+ scanchain_179/module_data_in[4] scanchain_179/module_data_in[5] scanchain_179/module_data_in[6]
+ scanchain_179/module_data_in[7] scanchain_179/module_data_out[0] scanchain_179/module_data_out[1]
+ scanchain_179/module_data_out[2] scanchain_179/module_data_out[3] scanchain_179/module_data_out[4]
+ scanchain_179/module_data_out[5] scanchain_179/module_data_out[6] scanchain_179/module_data_out[7]
+ scanchain_179/scan_select_in scanchain_180/scan_select_in vccd1 vssd1 scanchain
Xjleightcap_top_54 jleightcap_top_54/io_in[0] jleightcap_top_54/io_in[1] jleightcap_top_54/io_in[2]
+ jleightcap_top_54/io_in[3] jleightcap_top_54/io_in[4] jleightcap_top_54/io_in[5]
+ jleightcap_top_54/io_in[6] jleightcap_top_54/io_in[7] jleightcap_top_54/io_out[0]
+ jleightcap_top_54/io_out[1] jleightcap_top_54/io_out[2] jleightcap_top_54/io_out[3]
+ jleightcap_top_54/io_out[4] jleightcap_top_54/io_out[5] jleightcap_top_54/io_out[6]
+ jleightcap_top_54/io_out[7] vccd1 vssd1 jleightcap_top
Xuser_module_339501025136214612_0 scanchain_0/module_data_in[0] scanchain_0/module_data_in[1]
+ scanchain_0/module_data_in[2] scanchain_0/module_data_in[3] scanchain_0/module_data_in[4]
+ scanchain_0/module_data_in[5] scanchain_0/module_data_in[6] scanchain_0/module_data_in[7]
+ scanchain_0/module_data_out[0] scanchain_0/module_data_out[1] scanchain_0/module_data_out[2]
+ scanchain_0/module_data_out[3] scanchain_0/module_data_out[4] scanchain_0/module_data_out[5]
+ scanchain_0/module_data_out[6] scanchain_0/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_397 scanchain_397/module_data_in[0] scanchain_397/module_data_in[1]
+ scanchain_397/module_data_in[2] scanchain_397/module_data_in[3] scanchain_397/module_data_in[4]
+ scanchain_397/module_data_in[5] scanchain_397/module_data_in[6] scanchain_397/module_data_in[7]
+ scanchain_397/module_data_out[0] scanchain_397/module_data_out[1] scanchain_397/module_data_out[2]
+ scanchain_397/module_data_out[3] scanchain_397/module_data_out[4] scanchain_397/module_data_out[5]
+ scanchain_397/module_data_out[6] scanchain_397/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_386 scanchain_386/module_data_in[0] scanchain_386/module_data_in[1]
+ scanchain_386/module_data_in[2] scanchain_386/module_data_in[3] scanchain_386/module_data_in[4]
+ scanchain_386/module_data_in[5] scanchain_386/module_data_in[6] scanchain_386/module_data_in[7]
+ scanchain_386/module_data_out[0] scanchain_386/module_data_out[1] scanchain_386/module_data_out[2]
+ scanchain_386/module_data_out[3] scanchain_386/module_data_out[4] scanchain_386/module_data_out[5]
+ scanchain_386/module_data_out[6] scanchain_386/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_364 scanchain_364/module_data_in[0] scanchain_364/module_data_in[1]
+ scanchain_364/module_data_in[2] scanchain_364/module_data_in[3] scanchain_364/module_data_in[4]
+ scanchain_364/module_data_in[5] scanchain_364/module_data_in[6] scanchain_364/module_data_in[7]
+ scanchain_364/module_data_out[0] scanchain_364/module_data_out[1] scanchain_364/module_data_out[2]
+ scanchain_364/module_data_out[3] scanchain_364/module_data_out[4] scanchain_364/module_data_out[5]
+ scanchain_364/module_data_out[6] scanchain_364/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_375 scanchain_375/module_data_in[0] scanchain_375/module_data_in[1]
+ scanchain_375/module_data_in[2] scanchain_375/module_data_in[3] scanchain_375/module_data_in[4]
+ scanchain_375/module_data_in[5] scanchain_375/module_data_in[6] scanchain_375/module_data_in[7]
+ scanchain_375/module_data_out[0] scanchain_375/module_data_out[1] scanchain_375/module_data_out[2]
+ scanchain_375/module_data_out[3] scanchain_375/module_data_out[4] scanchain_375/module_data_out[5]
+ scanchain_375/module_data_out[6] scanchain_375/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_353 scanchain_353/module_data_in[0] scanchain_353/module_data_in[1]
+ scanchain_353/module_data_in[2] scanchain_353/module_data_in[3] scanchain_353/module_data_in[4]
+ scanchain_353/module_data_in[5] scanchain_353/module_data_in[6] scanchain_353/module_data_in[7]
+ scanchain_353/module_data_out[0] scanchain_353/module_data_out[1] scanchain_353/module_data_out[2]
+ scanchain_353/module_data_out[3] scanchain_353/module_data_out[4] scanchain_353/module_data_out[5]
+ scanchain_353/module_data_out[6] scanchain_353/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_342 scanchain_342/module_data_in[0] scanchain_342/module_data_in[1]
+ scanchain_342/module_data_in[2] scanchain_342/module_data_in[3] scanchain_342/module_data_in[4]
+ scanchain_342/module_data_in[5] scanchain_342/module_data_in[6] scanchain_342/module_data_in[7]
+ scanchain_342/module_data_out[0] scanchain_342/module_data_out[1] scanchain_342/module_data_out[2]
+ scanchain_342/module_data_out[3] scanchain_342/module_data_out[4] scanchain_342/module_data_out[5]
+ scanchain_342/module_data_out[6] scanchain_342/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_328 scanchain_328/clk_in scanchain_329/clk_in scanchain_328/data_in scanchain_329/data_in
+ scanchain_328/latch_enable_in scanchain_329/latch_enable_in scanchain_328/module_data_in[0]
+ scanchain_328/module_data_in[1] scanchain_328/module_data_in[2] scanchain_328/module_data_in[3]
+ scanchain_328/module_data_in[4] scanchain_328/module_data_in[5] scanchain_328/module_data_in[6]
+ scanchain_328/module_data_in[7] scanchain_328/module_data_out[0] scanchain_328/module_data_out[1]
+ scanchain_328/module_data_out[2] scanchain_328/module_data_out[3] scanchain_328/module_data_out[4]
+ scanchain_328/module_data_out[5] scanchain_328/module_data_out[6] scanchain_328/module_data_out[7]
+ scanchain_328/scan_select_in scanchain_329/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_331 scanchain_331/module_data_in[0] scanchain_331/module_data_in[1]
+ scanchain_331/module_data_in[2] scanchain_331/module_data_in[3] scanchain_331/module_data_in[4]
+ scanchain_331/module_data_in[5] scanchain_331/module_data_in[6] scanchain_331/module_data_in[7]
+ scanchain_331/module_data_out[0] scanchain_331/module_data_out[1] scanchain_331/module_data_out[2]
+ scanchain_331/module_data_out[3] scanchain_331/module_data_out[4] scanchain_331/module_data_out[5]
+ scanchain_331/module_data_out[6] scanchain_331/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_339 scanchain_339/clk_in scanchain_340/clk_in scanchain_339/data_in scanchain_340/data_in
+ scanchain_339/latch_enable_in scanchain_340/latch_enable_in scanchain_339/module_data_in[0]
+ scanchain_339/module_data_in[1] scanchain_339/module_data_in[2] scanchain_339/module_data_in[3]
+ scanchain_339/module_data_in[4] scanchain_339/module_data_in[5] scanchain_339/module_data_in[6]
+ scanchain_339/module_data_in[7] scanchain_339/module_data_out[0] scanchain_339/module_data_out[1]
+ scanchain_339/module_data_out[2] scanchain_339/module_data_out[3] scanchain_339/module_data_out[4]
+ scanchain_339/module_data_out[5] scanchain_339/module_data_out[6] scanchain_339/module_data_out[7]
+ scanchain_339/scan_select_in scanchain_340/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_320 scanchain_320/module_data_in[0] scanchain_320/module_data_in[1]
+ scanchain_320/module_data_in[2] scanchain_320/module_data_in[3] scanchain_320/module_data_in[4]
+ scanchain_320/module_data_in[5] scanchain_320/module_data_in[6] scanchain_320/module_data_in[7]
+ scanchain_320/module_data_out[0] scanchain_320/module_data_out[1] scanchain_320/module_data_out[2]
+ scanchain_320/module_data_out[3] scanchain_320/module_data_out[4] scanchain_320/module_data_out[5]
+ scanchain_320/module_data_out[6] scanchain_320/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_317 scanchain_317/clk_in scanchain_318/clk_in scanchain_317/data_in scanchain_318/data_in
+ scanchain_317/latch_enable_in scanchain_318/latch_enable_in scanchain_317/module_data_in[0]
+ scanchain_317/module_data_in[1] scanchain_317/module_data_in[2] scanchain_317/module_data_in[3]
+ scanchain_317/module_data_in[4] scanchain_317/module_data_in[5] scanchain_317/module_data_in[6]
+ scanchain_317/module_data_in[7] scanchain_317/module_data_out[0] scanchain_317/module_data_out[1]
+ scanchain_317/module_data_out[2] scanchain_317/module_data_out[3] scanchain_317/module_data_out[4]
+ scanchain_317/module_data_out[5] scanchain_317/module_data_out[6] scanchain_317/module_data_out[7]
+ scanchain_317/scan_select_in scanchain_318/scan_select_in vccd1 vssd1 scanchain
Xscanchain_306 scanchain_306/clk_in scanchain_307/clk_in scanchain_306/data_in scanchain_307/data_in
+ scanchain_306/latch_enable_in scanchain_307/latch_enable_in scanchain_306/module_data_in[0]
+ scanchain_306/module_data_in[1] scanchain_306/module_data_in[2] scanchain_306/module_data_in[3]
+ scanchain_306/module_data_in[4] scanchain_306/module_data_in[5] scanchain_306/module_data_in[6]
+ scanchain_306/module_data_in[7] scanchain_306/module_data_out[0] scanchain_306/module_data_out[1]
+ scanchain_306/module_data_out[2] scanchain_306/module_data_out[3] scanchain_306/module_data_out[4]
+ scanchain_306/module_data_out[5] scanchain_306/module_data_out[6] scanchain_306/module_data_out[7]
+ scanchain_306/scan_select_in scanchain_307/scan_select_in vccd1 vssd1 scanchain
Xuser_module_348195845106041428_27 scanchain_27/module_data_in[0] scanchain_27/module_data_in[1]
+ scanchain_27/module_data_in[2] scanchain_27/module_data_in[3] scanchain_27/module_data_in[4]
+ scanchain_27/module_data_in[5] scanchain_27/module_data_in[6] scanchain_27/module_data_in[7]
+ scanchain_27/module_data_out[0] scanchain_27/module_data_out[1] scanchain_27/module_data_out[2]
+ scanchain_27/module_data_out[3] scanchain_27/module_data_out[4] scanchain_27/module_data_out[5]
+ scanchain_27/module_data_out[6] scanchain_27/module_data_out[7] vccd1 vssd1 user_module_348195845106041428
Xuser_module_339501025136214612_194 scanchain_194/module_data_in[0] scanchain_194/module_data_in[1]
+ scanchain_194/module_data_in[2] scanchain_194/module_data_in[3] scanchain_194/module_data_in[4]
+ scanchain_194/module_data_in[5] scanchain_194/module_data_in[6] scanchain_194/module_data_in[7]
+ scanchain_194/module_data_out[0] scanchain_194/module_data_out[1] scanchain_194/module_data_out[2]
+ scanchain_194/module_data_out[3] scanchain_194/module_data_out[4] scanchain_194/module_data_out[5]
+ scanchain_194/module_data_out[6] scanchain_194/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_103 scanchain_103/clk_in scanchain_104/clk_in scanchain_103/data_in scanchain_104/data_in
+ scanchain_103/latch_enable_in scanchain_104/latch_enable_in scanchain_103/module_data_in[0]
+ scanchain_103/module_data_in[1] scanchain_103/module_data_in[2] scanchain_103/module_data_in[3]
+ scanchain_103/module_data_in[4] scanchain_103/module_data_in[5] scanchain_103/module_data_in[6]
+ scanchain_103/module_data_in[7] scanchain_103/module_data_out[0] scanchain_103/module_data_out[1]
+ scanchain_103/module_data_out[2] scanchain_103/module_data_out[3] scanchain_103/module_data_out[4]
+ scanchain_103/module_data_out[5] scanchain_103/module_data_out[6] scanchain_103/module_data_out[7]
+ scanchain_103/scan_select_in scanchain_104/scan_select_in vccd1 vssd1 scanchain
Xscanchain_114 scanchain_114/clk_in scanchain_115/clk_in scanchain_114/data_in scanchain_115/data_in
+ scanchain_114/latch_enable_in scanchain_115/latch_enable_in scanchain_114/module_data_in[0]
+ scanchain_114/module_data_in[1] scanchain_114/module_data_in[2] scanchain_114/module_data_in[3]
+ scanchain_114/module_data_in[4] scanchain_114/module_data_in[5] scanchain_114/module_data_in[6]
+ scanchain_114/module_data_in[7] scanchain_114/module_data_out[0] scanchain_114/module_data_out[1]
+ scanchain_114/module_data_out[2] scanchain_114/module_data_out[3] scanchain_114/module_data_out[4]
+ scanchain_114/module_data_out[5] scanchain_114/module_data_out[6] scanchain_114/module_data_out[7]
+ scanchain_114/scan_select_in scanchain_115/scan_select_in vccd1 vssd1 scanchain
Xscanchain_125 scanchain_125/clk_in scanchain_126/clk_in scanchain_125/data_in scanchain_126/data_in
+ scanchain_125/latch_enable_in scanchain_126/latch_enable_in scanchain_125/module_data_in[0]
+ scanchain_125/module_data_in[1] scanchain_125/module_data_in[2] scanchain_125/module_data_in[3]
+ scanchain_125/module_data_in[4] scanchain_125/module_data_in[5] scanchain_125/module_data_in[6]
+ scanchain_125/module_data_in[7] scanchain_125/module_data_out[0] scanchain_125/module_data_out[1]
+ scanchain_125/module_data_out[2] scanchain_125/module_data_out[3] scanchain_125/module_data_out[4]
+ scanchain_125/module_data_out[5] scanchain_125/module_data_out[6] scanchain_125/module_data_out[7]
+ scanchain_125/scan_select_in scanchain_126/scan_select_in vccd1 vssd1 scanchain
Xscanchain_147 scanchain_147/clk_in scanchain_148/clk_in scanchain_147/data_in scanchain_148/data_in
+ scanchain_147/latch_enable_in scanchain_148/latch_enable_in scanchain_147/module_data_in[0]
+ scanchain_147/module_data_in[1] scanchain_147/module_data_in[2] scanchain_147/module_data_in[3]
+ scanchain_147/module_data_in[4] scanchain_147/module_data_in[5] scanchain_147/module_data_in[6]
+ scanchain_147/module_data_in[7] scanchain_147/module_data_out[0] scanchain_147/module_data_out[1]
+ scanchain_147/module_data_out[2] scanchain_147/module_data_out[3] scanchain_147/module_data_out[4]
+ scanchain_147/module_data_out[5] scanchain_147/module_data_out[6] scanchain_147/module_data_out[7]
+ scanchain_147/scan_select_in scanchain_148/scan_select_in vccd1 vssd1 scanchain
Xscanchain_136 scanchain_136/clk_in scanchain_137/clk_in scanchain_136/data_in scanchain_137/data_in
+ scanchain_136/latch_enable_in scanchain_137/latch_enable_in scanchain_136/module_data_in[0]
+ scanchain_136/module_data_in[1] scanchain_136/module_data_in[2] scanchain_136/module_data_in[3]
+ scanchain_136/module_data_in[4] scanchain_136/module_data_in[5] scanchain_136/module_data_in[6]
+ scanchain_136/module_data_in[7] scanchain_136/module_data_out[0] scanchain_136/module_data_out[1]
+ scanchain_136/module_data_out[2] scanchain_136/module_data_out[3] scanchain_136/module_data_out[4]
+ scanchain_136/module_data_out[5] scanchain_136/module_data_out[6] scanchain_136/module_data_out[7]
+ scanchain_136/scan_select_in scanchain_137/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_150 scanchain_150/module_data_in[0] scanchain_150/module_data_in[1]
+ scanchain_150/module_data_in[2] scanchain_150/module_data_in[3] scanchain_150/module_data_in[4]
+ scanchain_150/module_data_in[5] scanchain_150/module_data_in[6] scanchain_150/module_data_in[7]
+ scanchain_150/module_data_out[0] scanchain_150/module_data_out[1] scanchain_150/module_data_out[2]
+ scanchain_150/module_data_out[3] scanchain_150/module_data_out[4] scanchain_150/module_data_out[5]
+ scanchain_150/module_data_out[6] scanchain_150/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_158 scanchain_158/clk_in scanchain_159/clk_in scanchain_158/data_in scanchain_159/data_in
+ scanchain_158/latch_enable_in scanchain_159/latch_enable_in scanchain_158/module_data_in[0]
+ scanchain_158/module_data_in[1] scanchain_158/module_data_in[2] scanchain_158/module_data_in[3]
+ scanchain_158/module_data_in[4] scanchain_158/module_data_in[5] scanchain_158/module_data_in[6]
+ scanchain_158/module_data_in[7] scanchain_158/module_data_out[0] scanchain_158/module_data_out[1]
+ scanchain_158/module_data_out[2] scanchain_158/module_data_out[3] scanchain_158/module_data_out[4]
+ scanchain_158/module_data_out[5] scanchain_158/module_data_out[6] scanchain_158/module_data_out[7]
+ scanchain_158/scan_select_in scanchain_159/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_161 scanchain_161/module_data_in[0] scanchain_161/module_data_in[1]
+ scanchain_161/module_data_in[2] scanchain_161/module_data_in[3] scanchain_161/module_data_in[4]
+ scanchain_161/module_data_in[5] scanchain_161/module_data_in[6] scanchain_161/module_data_in[7]
+ scanchain_161/module_data_out[0] scanchain_161/module_data_out[1] scanchain_161/module_data_out[2]
+ scanchain_161/module_data_out[3] scanchain_161/module_data_out[4] scanchain_161/module_data_out[5]
+ scanchain_161/module_data_out[6] scanchain_161/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_183 scanchain_183/module_data_in[0] scanchain_183/module_data_in[1]
+ scanchain_183/module_data_in[2] scanchain_183/module_data_in[3] scanchain_183/module_data_in[4]
+ scanchain_183/module_data_in[5] scanchain_183/module_data_in[6] scanchain_183/module_data_in[7]
+ scanchain_183/module_data_out[0] scanchain_183/module_data_out[1] scanchain_183/module_data_out[2]
+ scanchain_183/module_data_out[3] scanchain_183/module_data_out[4] scanchain_183/module_data_out[5]
+ scanchain_183/module_data_out[6] scanchain_183/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_172 scanchain_172/module_data_in[0] scanchain_172/module_data_in[1]
+ scanchain_172/module_data_in[2] scanchain_172/module_data_in[3] scanchain_172/module_data_in[4]
+ scanchain_172/module_data_in[5] scanchain_172/module_data_in[6] scanchain_172/module_data_in[7]
+ scanchain_172/module_data_out[0] scanchain_172/module_data_out[1] scanchain_172/module_data_out[2]
+ scanchain_172/module_data_out[3] scanchain_172/module_data_out[4] scanchain_172/module_data_out[5]
+ scanchain_172/module_data_out[6] scanchain_172/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_169 scanchain_169/clk_in scanchain_170/clk_in scanchain_169/data_in scanchain_170/data_in
+ scanchain_169/latch_enable_in scanchain_170/latch_enable_in scanchain_169/module_data_in[0]
+ scanchain_169/module_data_in[1] scanchain_169/module_data_in[2] scanchain_169/module_data_in[3]
+ scanchain_169/module_data_in[4] scanchain_169/module_data_in[5] scanchain_169/module_data_in[6]
+ scanchain_169/module_data_in[7] scanchain_169/module_data_out[0] scanchain_169/module_data_out[1]
+ scanchain_169/module_data_out[2] scanchain_169/module_data_out[3] scanchain_169/module_data_out[4]
+ scanchain_169/module_data_out[5] scanchain_169/module_data_out[6] scanchain_169/module_data_out[7]
+ scanchain_169/scan_select_in scanchain_170/scan_select_in vccd1 vssd1 scanchain
Xxor_shift32_quantamhd_51 scanchain_51/module_data_in[0] scanchain_51/module_data_in[1]
+ scanchain_51/module_data_in[2] scanchain_51/module_data_in[3] scanchain_51/module_data_in[4]
+ scanchain_51/module_data_in[5] scanchain_51/module_data_in[6] scanchain_51/module_data_in[7]
+ scanchain_51/module_data_out[0] scanchain_51/module_data_out[1] scanchain_51/module_data_out[2]
+ scanchain_51/module_data_out[3] scanchain_51/module_data_out[4] scanchain_51/module_data_out[5]
+ scanchain_51/module_data_out[6] scanchain_51/module_data_out[7] vccd1 vssd1 xor_shift32_quantamhd
Xmbikovitsky_top_33 mbikovitsky_top_33/io_in[0] mbikovitsky_top_33/io_in[1] mbikovitsky_top_33/io_in[2]
+ mbikovitsky_top_33/io_in[3] mbikovitsky_top_33/io_in[4] mbikovitsky_top_33/io_in[5]
+ mbikovitsky_top_33/io_in[6] mbikovitsky_top_33/io_in[7] mbikovitsky_top_33/io_out[0]
+ mbikovitsky_top_33/io_out[1] mbikovitsky_top_33/io_out[2] mbikovitsky_top_33/io_out[3]
+ mbikovitsky_top_33/io_out[4] mbikovitsky_top_33/io_out[5] mbikovitsky_top_33/io_out[6]
+ mbikovitsky_top_33/io_out[7] vccd1 vssd1 mbikovitsky_top
Xmeriac_tt02_play_tune_45 scanchain_45/module_data_in[0] scanchain_45/module_data_in[1]
+ scanchain_45/module_data_in[2] scanchain_45/module_data_in[3] scanchain_45/module_data_in[4]
+ scanchain_45/module_data_in[5] scanchain_45/module_data_in[6] scanchain_45/module_data_in[7]
+ scanchain_45/module_data_out[0] scanchain_45/module_data_out[1] scanchain_45/module_data_out[2]
+ scanchain_45/module_data_out[3] scanchain_45/module_data_out[4] scanchain_45/module_data_out[5]
+ scanchain_45/module_data_out[6] scanchain_45/module_data_out[7] vccd1 vssd1 meriac_tt02_play_tune
Xuser_module_339501025136214612_398 scanchain_398/module_data_in[0] scanchain_398/module_data_in[1]
+ scanchain_398/module_data_in[2] scanchain_398/module_data_in[3] scanchain_398/module_data_in[4]
+ scanchain_398/module_data_in[5] scanchain_398/module_data_in[6] scanchain_398/module_data_in[7]
+ scanchain_398/module_data_out[0] scanchain_398/module_data_out[1] scanchain_398/module_data_out[2]
+ scanchain_398/module_data_out[3] scanchain_398/module_data_out[4] scanchain_398/module_data_out[5]
+ scanchain_398/module_data_out[6] scanchain_398/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_387 scanchain_387/module_data_in[0] scanchain_387/module_data_in[1]
+ scanchain_387/module_data_in[2] scanchain_387/module_data_in[3] scanchain_387/module_data_in[4]
+ scanchain_387/module_data_in[5] scanchain_387/module_data_in[6] scanchain_387/module_data_in[7]
+ scanchain_387/module_data_out[0] scanchain_387/module_data_out[1] scanchain_387/module_data_out[2]
+ scanchain_387/module_data_out[3] scanchain_387/module_data_out[4] scanchain_387/module_data_out[5]
+ scanchain_387/module_data_out[6] scanchain_387/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_365 scanchain_365/module_data_in[0] scanchain_365/module_data_in[1]
+ scanchain_365/module_data_in[2] scanchain_365/module_data_in[3] scanchain_365/module_data_in[4]
+ scanchain_365/module_data_in[5] scanchain_365/module_data_in[6] scanchain_365/module_data_in[7]
+ scanchain_365/module_data_out[0] scanchain_365/module_data_out[1] scanchain_365/module_data_out[2]
+ scanchain_365/module_data_out[3] scanchain_365/module_data_out[4] scanchain_365/module_data_out[5]
+ scanchain_365/module_data_out[6] scanchain_365/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_376 scanchain_376/module_data_in[0] scanchain_376/module_data_in[1]
+ scanchain_376/module_data_in[2] scanchain_376/module_data_in[3] scanchain_376/module_data_in[4]
+ scanchain_376/module_data_in[5] scanchain_376/module_data_in[6] scanchain_376/module_data_in[7]
+ scanchain_376/module_data_out[0] scanchain_376/module_data_out[1] scanchain_376/module_data_out[2]
+ scanchain_376/module_data_out[3] scanchain_376/module_data_out[4] scanchain_376/module_data_out[5]
+ scanchain_376/module_data_out[6] scanchain_376/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_354 scanchain_354/module_data_in[0] scanchain_354/module_data_in[1]
+ scanchain_354/module_data_in[2] scanchain_354/module_data_in[3] scanchain_354/module_data_in[4]
+ scanchain_354/module_data_in[5] scanchain_354/module_data_in[6] scanchain_354/module_data_in[7]
+ scanchain_354/module_data_out[0] scanchain_354/module_data_out[1] scanchain_354/module_data_out[2]
+ scanchain_354/module_data_out[3] scanchain_354/module_data_out[4] scanchain_354/module_data_out[5]
+ scanchain_354/module_data_out[6] scanchain_354/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_343 scanchain_343/module_data_in[0] scanchain_343/module_data_in[1]
+ scanchain_343/module_data_in[2] scanchain_343/module_data_in[3] scanchain_343/module_data_in[4]
+ scanchain_343/module_data_in[5] scanchain_343/module_data_in[6] scanchain_343/module_data_in[7]
+ scanchain_343/module_data_out[0] scanchain_343/module_data_out[1] scanchain_343/module_data_out[2]
+ scanchain_343/module_data_out[3] scanchain_343/module_data_out[4] scanchain_343/module_data_out[5]
+ scanchain_343/module_data_out[6] scanchain_343/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_321 scanchain_321/module_data_in[0] scanchain_321/module_data_in[1]
+ scanchain_321/module_data_in[2] scanchain_321/module_data_in[3] scanchain_321/module_data_in[4]
+ scanchain_321/module_data_in[5] scanchain_321/module_data_in[6] scanchain_321/module_data_in[7]
+ scanchain_321/module_data_out[0] scanchain_321/module_data_out[1] scanchain_321/module_data_out[2]
+ scanchain_321/module_data_out[3] scanchain_321/module_data_out[4] scanchain_321/module_data_out[5]
+ scanchain_321/module_data_out[6] scanchain_321/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_332 scanchain_332/module_data_in[0] scanchain_332/module_data_in[1]
+ scanchain_332/module_data_in[2] scanchain_332/module_data_in[3] scanchain_332/module_data_in[4]
+ scanchain_332/module_data_in[5] scanchain_332/module_data_in[6] scanchain_332/module_data_in[7]
+ scanchain_332/module_data_out[0] scanchain_332/module_data_out[1] scanchain_332/module_data_out[2]
+ scanchain_332/module_data_out[3] scanchain_332/module_data_out[4] scanchain_332/module_data_out[5]
+ scanchain_332/module_data_out[6] scanchain_332/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_310 scanchain_310/module_data_in[0] scanchain_310/module_data_in[1]
+ scanchain_310/module_data_in[2] scanchain_310/module_data_in[3] scanchain_310/module_data_in[4]
+ scanchain_310/module_data_in[5] scanchain_310/module_data_in[6] scanchain_310/module_data_in[7]
+ scanchain_310/module_data_out[0] scanchain_310/module_data_out[1] scanchain_310/module_data_out[2]
+ scanchain_310/module_data_out[3] scanchain_310/module_data_out[4] scanchain_310/module_data_out[5]
+ scanchain_310/module_data_out[6] scanchain_310/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_307 scanchain_307/clk_in scanchain_308/clk_in scanchain_307/data_in scanchain_308/data_in
+ scanchain_307/latch_enable_in scanchain_308/latch_enable_in scanchain_307/module_data_in[0]
+ scanchain_307/module_data_in[1] scanchain_307/module_data_in[2] scanchain_307/module_data_in[3]
+ scanchain_307/module_data_in[4] scanchain_307/module_data_in[5] scanchain_307/module_data_in[6]
+ scanchain_307/module_data_in[7] scanchain_307/module_data_out[0] scanchain_307/module_data_out[1]
+ scanchain_307/module_data_out[2] scanchain_307/module_data_out[3] scanchain_307/module_data_out[4]
+ scanchain_307/module_data_out[5] scanchain_307/module_data_out[6] scanchain_307/module_data_out[7]
+ scanchain_307/scan_select_in scanchain_308/scan_select_in vccd1 vssd1 scanchain
Xscanchain_329 scanchain_329/clk_in scanchain_330/clk_in scanchain_329/data_in scanchain_330/data_in
+ scanchain_329/latch_enable_in scanchain_330/latch_enable_in scanchain_329/module_data_in[0]
+ scanchain_329/module_data_in[1] scanchain_329/module_data_in[2] scanchain_329/module_data_in[3]
+ scanchain_329/module_data_in[4] scanchain_329/module_data_in[5] scanchain_329/module_data_in[6]
+ scanchain_329/module_data_in[7] scanchain_329/module_data_out[0] scanchain_329/module_data_out[1]
+ scanchain_329/module_data_out[2] scanchain_329/module_data_out[3] scanchain_329/module_data_out[4]
+ scanchain_329/module_data_out[5] scanchain_329/module_data_out[6] scanchain_329/module_data_out[7]
+ scanchain_329/scan_select_in scanchain_330/scan_select_in vccd1 vssd1 scanchain
Xscanchain_318 scanchain_318/clk_in scanchain_319/clk_in scanchain_318/data_in scanchain_319/data_in
+ scanchain_318/latch_enable_in scanchain_319/latch_enable_in scanchain_318/module_data_in[0]
+ scanchain_318/module_data_in[1] scanchain_318/module_data_in[2] scanchain_318/module_data_in[3]
+ scanchain_318/module_data_in[4] scanchain_318/module_data_in[5] scanchain_318/module_data_in[6]
+ scanchain_318/module_data_in[7] scanchain_318/module_data_out[0] scanchain_318/module_data_out[1]
+ scanchain_318/module_data_out[2] scanchain_318/module_data_out[3] scanchain_318/module_data_out[4]
+ scanchain_318/module_data_out[5] scanchain_318/module_data_out[6] scanchain_318/module_data_out[7]
+ scanchain_318/scan_select_in scanchain_319/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_195 scanchain_195/module_data_in[0] scanchain_195/module_data_in[1]
+ scanchain_195/module_data_in[2] scanchain_195/module_data_in[3] scanchain_195/module_data_in[4]
+ scanchain_195/module_data_in[5] scanchain_195/module_data_in[6] scanchain_195/module_data_in[7]
+ scanchain_195/module_data_out[0] scanchain_195/module_data_out[1] scanchain_195/module_data_out[2]
+ scanchain_195/module_data_out[3] scanchain_195/module_data_out[4] scanchain_195/module_data_out[5]
+ scanchain_195/module_data_out[6] scanchain_195/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_104 scanchain_104/clk_in scanchain_105/clk_in scanchain_104/data_in scanchain_105/data_in
+ scanchain_104/latch_enable_in scanchain_105/latch_enable_in scanchain_104/module_data_in[0]
+ scanchain_104/module_data_in[1] scanchain_104/module_data_in[2] scanchain_104/module_data_in[3]
+ scanchain_104/module_data_in[4] scanchain_104/module_data_in[5] scanchain_104/module_data_in[6]
+ scanchain_104/module_data_in[7] scanchain_104/module_data_out[0] scanchain_104/module_data_out[1]
+ scanchain_104/module_data_out[2] scanchain_104/module_data_out[3] scanchain_104/module_data_out[4]
+ scanchain_104/module_data_out[5] scanchain_104/module_data_out[6] scanchain_104/module_data_out[7]
+ scanchain_104/scan_select_in scanchain_105/scan_select_in vccd1 vssd1 scanchain
Xscanchain_115 scanchain_115/clk_in scanchain_116/clk_in scanchain_115/data_in scanchain_116/data_in
+ scanchain_115/latch_enable_in scanchain_116/latch_enable_in scanchain_115/module_data_in[0]
+ scanchain_115/module_data_in[1] scanchain_115/module_data_in[2] scanchain_115/module_data_in[3]
+ scanchain_115/module_data_in[4] scanchain_115/module_data_in[5] scanchain_115/module_data_in[6]
+ scanchain_115/module_data_in[7] scanchain_115/module_data_out[0] scanchain_115/module_data_out[1]
+ scanchain_115/module_data_out[2] scanchain_115/module_data_out[3] scanchain_115/module_data_out[4]
+ scanchain_115/module_data_out[5] scanchain_115/module_data_out[6] scanchain_115/module_data_out[7]
+ scanchain_115/scan_select_in scanchain_116/scan_select_in vccd1 vssd1 scanchain
Xscanchain_126 scanchain_126/clk_in scanchain_127/clk_in scanchain_126/data_in scanchain_127/data_in
+ scanchain_126/latch_enable_in scanchain_127/latch_enable_in scanchain_126/module_data_in[0]
+ scanchain_126/module_data_in[1] scanchain_126/module_data_in[2] scanchain_126/module_data_in[3]
+ scanchain_126/module_data_in[4] scanchain_126/module_data_in[5] scanchain_126/module_data_in[6]
+ scanchain_126/module_data_in[7] scanchain_126/module_data_out[0] scanchain_126/module_data_out[1]
+ scanchain_126/module_data_out[2] scanchain_126/module_data_out[3] scanchain_126/module_data_out[4]
+ scanchain_126/module_data_out[5] scanchain_126/module_data_out[6] scanchain_126/module_data_out[7]
+ scanchain_126/scan_select_in scanchain_127/scan_select_in vccd1 vssd1 scanchain
Xscanchain_148 scanchain_148/clk_in scanchain_149/clk_in scanchain_148/data_in scanchain_149/data_in
+ scanchain_148/latch_enable_in scanchain_149/latch_enable_in scanchain_148/module_data_in[0]
+ scanchain_148/module_data_in[1] scanchain_148/module_data_in[2] scanchain_148/module_data_in[3]
+ scanchain_148/module_data_in[4] scanchain_148/module_data_in[5] scanchain_148/module_data_in[6]
+ scanchain_148/module_data_in[7] scanchain_148/module_data_out[0] scanchain_148/module_data_out[1]
+ scanchain_148/module_data_out[2] scanchain_148/module_data_out[3] scanchain_148/module_data_out[4]
+ scanchain_148/module_data_out[5] scanchain_148/module_data_out[6] scanchain_148/module_data_out[7]
+ scanchain_148/scan_select_in scanchain_149/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_140 scanchain_140/module_data_in[0] scanchain_140/module_data_in[1]
+ scanchain_140/module_data_in[2] scanchain_140/module_data_in[3] scanchain_140/module_data_in[4]
+ scanchain_140/module_data_in[5] scanchain_140/module_data_in[6] scanchain_140/module_data_in[7]
+ scanchain_140/module_data_out[0] scanchain_140/module_data_out[1] scanchain_140/module_data_out[2]
+ scanchain_140/module_data_out[3] scanchain_140/module_data_out[4] scanchain_140/module_data_out[5]
+ scanchain_140/module_data_out[6] scanchain_140/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_137 scanchain_137/clk_in scanchain_138/clk_in scanchain_137/data_in scanchain_138/data_in
+ scanchain_137/latch_enable_in scanchain_138/latch_enable_in scanchain_137/module_data_in[0]
+ scanchain_137/module_data_in[1] scanchain_137/module_data_in[2] scanchain_137/module_data_in[3]
+ scanchain_137/module_data_in[4] scanchain_137/module_data_in[5] scanchain_137/module_data_in[6]
+ scanchain_137/module_data_in[7] scanchain_137/module_data_out[0] scanchain_137/module_data_out[1]
+ scanchain_137/module_data_out[2] scanchain_137/module_data_out[3] scanchain_137/module_data_out[4]
+ scanchain_137/module_data_out[5] scanchain_137/module_data_out[6] scanchain_137/module_data_out[7]
+ scanchain_137/scan_select_in scanchain_138/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_151 scanchain_151/module_data_in[0] scanchain_151/module_data_in[1]
+ scanchain_151/module_data_in[2] scanchain_151/module_data_in[3] scanchain_151/module_data_in[4]
+ scanchain_151/module_data_in[5] scanchain_151/module_data_in[6] scanchain_151/module_data_in[7]
+ scanchain_151/module_data_out[0] scanchain_151/module_data_out[1] scanchain_151/module_data_out[2]
+ scanchain_151/module_data_out[3] scanchain_151/module_data_out[4] scanchain_151/module_data_out[5]
+ scanchain_151/module_data_out[6] scanchain_151/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_159 scanchain_159/clk_in scanchain_160/clk_in scanchain_159/data_in scanchain_160/data_in
+ scanchain_159/latch_enable_in scanchain_160/latch_enable_in scanchain_159/module_data_in[0]
+ scanchain_159/module_data_in[1] scanchain_159/module_data_in[2] scanchain_159/module_data_in[3]
+ scanchain_159/module_data_in[4] scanchain_159/module_data_in[5] scanchain_159/module_data_in[6]
+ scanchain_159/module_data_in[7] scanchain_159/module_data_out[0] scanchain_159/module_data_out[1]
+ scanchain_159/module_data_out[2] scanchain_159/module_data_out[3] scanchain_159/module_data_out[4]
+ scanchain_159/module_data_out[5] scanchain_159/module_data_out[6] scanchain_159/module_data_out[7]
+ scanchain_159/scan_select_in scanchain_160/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_162 scanchain_162/module_data_in[0] scanchain_162/module_data_in[1]
+ scanchain_162/module_data_in[2] scanchain_162/module_data_in[3] scanchain_162/module_data_in[4]
+ scanchain_162/module_data_in[5] scanchain_162/module_data_in[6] scanchain_162/module_data_in[7]
+ scanchain_162/module_data_out[0] scanchain_162/module_data_out[1] scanchain_162/module_data_out[2]
+ scanchain_162/module_data_out[3] scanchain_162/module_data_out[4] scanchain_162/module_data_out[5]
+ scanchain_162/module_data_out[6] scanchain_162/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_184 scanchain_184/module_data_in[0] scanchain_184/module_data_in[1]
+ scanchain_184/module_data_in[2] scanchain_184/module_data_in[3] scanchain_184/module_data_in[4]
+ scanchain_184/module_data_in[5] scanchain_184/module_data_in[6] scanchain_184/module_data_in[7]
+ scanchain_184/module_data_out[0] scanchain_184/module_data_out[1] scanchain_184/module_data_out[2]
+ scanchain_184/module_data_out[3] scanchain_184/module_data_out[4] scanchain_184/module_data_out[5]
+ scanchain_184/module_data_out[6] scanchain_184/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_173 scanchain_173/module_data_in[0] scanchain_173/module_data_in[1]
+ scanchain_173/module_data_in[2] scanchain_173/module_data_in[3] scanchain_173/module_data_in[4]
+ scanchain_173/module_data_in[5] scanchain_173/module_data_in[6] scanchain_173/module_data_in[7]
+ scanchain_173/module_data_out[0] scanchain_173/module_data_out[1] scanchain_173/module_data_out[2]
+ scanchain_173/module_data_out[3] scanchain_173/module_data_out[4] scanchain_173/module_data_out[5]
+ scanchain_173/module_data_out[6] scanchain_173/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_347690870424732244_12 scanchain_12/module_data_in[0] scanchain_12/module_data_in[1]
+ scanchain_12/module_data_in[2] scanchain_12/module_data_in[3] scanchain_12/module_data_in[4]
+ scanchain_12/module_data_in[5] scanchain_12/module_data_in[6] scanchain_12/module_data_in[7]
+ scanchain_12/module_data_out[0] scanchain_12/module_data_out[1] scanchain_12/module_data_out[2]
+ scanchain_12/module_data_out[3] scanchain_12/module_data_out[4] scanchain_12/module_data_out[5]
+ scanchain_12/module_data_out[6] scanchain_12/module_data_out[7] vccd1 vssd1 user_module_347690870424732244
Xuser_module_339501025136214612_399 scanchain_399/module_data_in[0] scanchain_399/module_data_in[1]
+ scanchain_399/module_data_in[2] scanchain_399/module_data_in[3] scanchain_399/module_data_in[4]
+ scanchain_399/module_data_in[5] scanchain_399/module_data_in[6] scanchain_399/module_data_in[7]
+ scanchain_399/module_data_out[0] scanchain_399/module_data_out[1] scanchain_399/module_data_out[2]
+ scanchain_399/module_data_out[3] scanchain_399/module_data_out[4] scanchain_399/module_data_out[5]
+ scanchain_399/module_data_out[6] scanchain_399/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_388 scanchain_388/module_data_in[0] scanchain_388/module_data_in[1]
+ scanchain_388/module_data_in[2] scanchain_388/module_data_in[3] scanchain_388/module_data_in[4]
+ scanchain_388/module_data_in[5] scanchain_388/module_data_in[6] scanchain_388/module_data_in[7]
+ scanchain_388/module_data_out[0] scanchain_388/module_data_out[1] scanchain_388/module_data_out[2]
+ scanchain_388/module_data_out[3] scanchain_388/module_data_out[4] scanchain_388/module_data_out[5]
+ scanchain_388/module_data_out[6] scanchain_388/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_366 scanchain_366/module_data_in[0] scanchain_366/module_data_in[1]
+ scanchain_366/module_data_in[2] scanchain_366/module_data_in[3] scanchain_366/module_data_in[4]
+ scanchain_366/module_data_in[5] scanchain_366/module_data_in[6] scanchain_366/module_data_in[7]
+ scanchain_366/module_data_out[0] scanchain_366/module_data_out[1] scanchain_366/module_data_out[2]
+ scanchain_366/module_data_out[3] scanchain_366/module_data_out[4] scanchain_366/module_data_out[5]
+ scanchain_366/module_data_out[6] scanchain_366/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_377 scanchain_377/module_data_in[0] scanchain_377/module_data_in[1]
+ scanchain_377/module_data_in[2] scanchain_377/module_data_in[3] scanchain_377/module_data_in[4]
+ scanchain_377/module_data_in[5] scanchain_377/module_data_in[6] scanchain_377/module_data_in[7]
+ scanchain_377/module_data_out[0] scanchain_377/module_data_out[1] scanchain_377/module_data_out[2]
+ scanchain_377/module_data_out[3] scanchain_377/module_data_out[4] scanchain_377/module_data_out[5]
+ scanchain_377/module_data_out[6] scanchain_377/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_355 scanchain_355/module_data_in[0] scanchain_355/module_data_in[1]
+ scanchain_355/module_data_in[2] scanchain_355/module_data_in[3] scanchain_355/module_data_in[4]
+ scanchain_355/module_data_in[5] scanchain_355/module_data_in[6] scanchain_355/module_data_in[7]
+ scanchain_355/module_data_out[0] scanchain_355/module_data_out[1] scanchain_355/module_data_out[2]
+ scanchain_355/module_data_out[3] scanchain_355/module_data_out[4] scanchain_355/module_data_out[5]
+ scanchain_355/module_data_out[6] scanchain_355/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_344 scanchain_344/module_data_in[0] scanchain_344/module_data_in[1]
+ scanchain_344/module_data_in[2] scanchain_344/module_data_in[3] scanchain_344/module_data_in[4]
+ scanchain_344/module_data_in[5] scanchain_344/module_data_in[6] scanchain_344/module_data_in[7]
+ scanchain_344/module_data_out[0] scanchain_344/module_data_out[1] scanchain_344/module_data_out[2]
+ scanchain_344/module_data_out[3] scanchain_344/module_data_out[4] scanchain_344/module_data_out[5]
+ scanchain_344/module_data_out[6] scanchain_344/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_322 scanchain_322/module_data_in[0] scanchain_322/module_data_in[1]
+ scanchain_322/module_data_in[2] scanchain_322/module_data_in[3] scanchain_322/module_data_in[4]
+ scanchain_322/module_data_in[5] scanchain_322/module_data_in[6] scanchain_322/module_data_in[7]
+ scanchain_322/module_data_out[0] scanchain_322/module_data_out[1] scanchain_322/module_data_out[2]
+ scanchain_322/module_data_out[3] scanchain_322/module_data_out[4] scanchain_322/module_data_out[5]
+ scanchain_322/module_data_out[6] scanchain_322/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_333 scanchain_333/module_data_in[0] scanchain_333/module_data_in[1]
+ scanchain_333/module_data_in[2] scanchain_333/module_data_in[3] scanchain_333/module_data_in[4]
+ scanchain_333/module_data_in[5] scanchain_333/module_data_in[6] scanchain_333/module_data_in[7]
+ scanchain_333/module_data_out[0] scanchain_333/module_data_out[1] scanchain_333/module_data_out[2]
+ scanchain_333/module_data_out[3] scanchain_333/module_data_out[4] scanchain_333/module_data_out[5]
+ scanchain_333/module_data_out[6] scanchain_333/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_311 scanchain_311/module_data_in[0] scanchain_311/module_data_in[1]
+ scanchain_311/module_data_in[2] scanchain_311/module_data_in[3] scanchain_311/module_data_in[4]
+ scanchain_311/module_data_in[5] scanchain_311/module_data_in[6] scanchain_311/module_data_in[7]
+ scanchain_311/module_data_out[0] scanchain_311/module_data_out[1] scanchain_311/module_data_out[2]
+ scanchain_311/module_data_out[3] scanchain_311/module_data_out[4] scanchain_311/module_data_out[5]
+ scanchain_311/module_data_out[6] scanchain_311/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_300 scanchain_300/module_data_in[0] scanchain_300/module_data_in[1]
+ scanchain_300/module_data_in[2] scanchain_300/module_data_in[3] scanchain_300/module_data_in[4]
+ scanchain_300/module_data_in[5] scanchain_300/module_data_in[6] scanchain_300/module_data_in[7]
+ scanchain_300/module_data_out[0] scanchain_300/module_data_out[1] scanchain_300/module_data_out[2]
+ scanchain_300/module_data_out[3] scanchain_300/module_data_out[4] scanchain_300/module_data_out[5]
+ scanchain_300/module_data_out[6] scanchain_300/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_319 scanchain_319/clk_in scanchain_320/clk_in scanchain_319/data_in scanchain_320/data_in
+ scanchain_319/latch_enable_in scanchain_320/latch_enable_in scanchain_319/module_data_in[0]
+ scanchain_319/module_data_in[1] scanchain_319/module_data_in[2] scanchain_319/module_data_in[3]
+ scanchain_319/module_data_in[4] scanchain_319/module_data_in[5] scanchain_319/module_data_in[6]
+ scanchain_319/module_data_in[7] scanchain_319/module_data_out[0] scanchain_319/module_data_out[1]
+ scanchain_319/module_data_out[2] scanchain_319/module_data_out[3] scanchain_319/module_data_out[4]
+ scanchain_319/module_data_out[5] scanchain_319/module_data_out[6] scanchain_319/module_data_out[7]
+ scanchain_319/scan_select_in scanchain_320/scan_select_in vccd1 vssd1 scanchain
Xscanchain_308 scanchain_308/clk_in scanchain_309/clk_in scanchain_308/data_in scanchain_309/data_in
+ scanchain_308/latch_enable_in scanchain_309/latch_enable_in scanchain_308/module_data_in[0]
+ scanchain_308/module_data_in[1] scanchain_308/module_data_in[2] scanchain_308/module_data_in[3]
+ scanchain_308/module_data_in[4] scanchain_308/module_data_in[5] scanchain_308/module_data_in[6]
+ scanchain_308/module_data_in[7] scanchain_308/module_data_out[0] scanchain_308/module_data_out[1]
+ scanchain_308/module_data_out[2] scanchain_308/module_data_out[3] scanchain_308/module_data_out[4]
+ scanchain_308/module_data_out[5] scanchain_308/module_data_out[6] scanchain_308/module_data_out[7]
+ scanchain_308/scan_select_in scanchain_309/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_196 scanchain_196/module_data_in[0] scanchain_196/module_data_in[1]
+ scanchain_196/module_data_in[2] scanchain_196/module_data_in[3] scanchain_196/module_data_in[4]
+ scanchain_196/module_data_in[5] scanchain_196/module_data_in[6] scanchain_196/module_data_in[7]
+ scanchain_196/module_data_out[0] scanchain_196/module_data_out[1] scanchain_196/module_data_out[2]
+ scanchain_196/module_data_out[3] scanchain_196/module_data_out[4] scanchain_196/module_data_out[5]
+ scanchain_196/module_data_out[6] scanchain_196/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_105 scanchain_105/clk_in scanchain_106/clk_in scanchain_105/data_in scanchain_106/data_in
+ scanchain_105/latch_enable_in scanchain_106/latch_enable_in scanchain_105/module_data_in[0]
+ scanchain_105/module_data_in[1] scanchain_105/module_data_in[2] scanchain_105/module_data_in[3]
+ scanchain_105/module_data_in[4] scanchain_105/module_data_in[5] scanchain_105/module_data_in[6]
+ scanchain_105/module_data_in[7] scanchain_105/module_data_out[0] scanchain_105/module_data_out[1]
+ scanchain_105/module_data_out[2] scanchain_105/module_data_out[3] scanchain_105/module_data_out[4]
+ scanchain_105/module_data_out[5] scanchain_105/module_data_out[6] scanchain_105/module_data_out[7]
+ scanchain_105/scan_select_in scanchain_106/scan_select_in vccd1 vssd1 scanchain
Xscanchain_116 scanchain_116/clk_in scanchain_117/clk_in scanchain_116/data_in scanchain_117/data_in
+ scanchain_116/latch_enable_in scanchain_117/latch_enable_in scanchain_116/module_data_in[0]
+ scanchain_116/module_data_in[1] scanchain_116/module_data_in[2] scanchain_116/module_data_in[3]
+ scanchain_116/module_data_in[4] scanchain_116/module_data_in[5] scanchain_116/module_data_in[6]
+ scanchain_116/module_data_in[7] scanchain_116/module_data_out[0] scanchain_116/module_data_out[1]
+ scanchain_116/module_data_out[2] scanchain_116/module_data_out[3] scanchain_116/module_data_out[4]
+ scanchain_116/module_data_out[5] scanchain_116/module_data_out[6] scanchain_116/module_data_out[7]
+ scanchain_116/scan_select_in scanchain_117/scan_select_in vccd1 vssd1 scanchain
Xscanchain_127 scanchain_127/clk_in scanchain_128/clk_in scanchain_127/data_in scanchain_128/data_in
+ scanchain_127/latch_enable_in scanchain_128/latch_enable_in scanchain_127/module_data_in[0]
+ scanchain_127/module_data_in[1] scanchain_127/module_data_in[2] scanchain_127/module_data_in[3]
+ scanchain_127/module_data_in[4] scanchain_127/module_data_in[5] scanchain_127/module_data_in[6]
+ scanchain_127/module_data_in[7] scanchain_127/module_data_out[0] scanchain_127/module_data_out[1]
+ scanchain_127/module_data_out[2] scanchain_127/module_data_out[3] scanchain_127/module_data_out[4]
+ scanchain_127/module_data_out[5] scanchain_127/module_data_out[6] scanchain_127/module_data_out[7]
+ scanchain_127/scan_select_in scanchain_128/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_130 scanchain_130/module_data_in[0] scanchain_130/module_data_in[1]
+ scanchain_130/module_data_in[2] scanchain_130/module_data_in[3] scanchain_130/module_data_in[4]
+ scanchain_130/module_data_in[5] scanchain_130/module_data_in[6] scanchain_130/module_data_in[7]
+ scanchain_130/module_data_out[0] scanchain_130/module_data_out[1] scanchain_130/module_data_out[2]
+ scanchain_130/module_data_out[3] scanchain_130/module_data_out[4] scanchain_130/module_data_out[5]
+ scanchain_130/module_data_out[6] scanchain_130/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_149 scanchain_149/clk_in scanchain_150/clk_in scanchain_149/data_in scanchain_150/data_in
+ scanchain_149/latch_enable_in scanchain_150/latch_enable_in scanchain_149/module_data_in[0]
+ scanchain_149/module_data_in[1] scanchain_149/module_data_in[2] scanchain_149/module_data_in[3]
+ scanchain_149/module_data_in[4] scanchain_149/module_data_in[5] scanchain_149/module_data_in[6]
+ scanchain_149/module_data_in[7] scanchain_149/module_data_out[0] scanchain_149/module_data_out[1]
+ scanchain_149/module_data_out[2] scanchain_149/module_data_out[3] scanchain_149/module_data_out[4]
+ scanchain_149/module_data_out[5] scanchain_149/module_data_out[6] scanchain_149/module_data_out[7]
+ scanchain_149/scan_select_in scanchain_150/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_141 scanchain_141/module_data_in[0] scanchain_141/module_data_in[1]
+ scanchain_141/module_data_in[2] scanchain_141/module_data_in[3] scanchain_141/module_data_in[4]
+ scanchain_141/module_data_in[5] scanchain_141/module_data_in[6] scanchain_141/module_data_in[7]
+ scanchain_141/module_data_out[0] scanchain_141/module_data_out[1] scanchain_141/module_data_out[2]
+ scanchain_141/module_data_out[3] scanchain_141/module_data_out[4] scanchain_141/module_data_out[5]
+ scanchain_141/module_data_out[6] scanchain_141/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_138 scanchain_138/clk_in scanchain_139/clk_in scanchain_138/data_in scanchain_139/data_in
+ scanchain_138/latch_enable_in scanchain_139/latch_enable_in scanchain_138/module_data_in[0]
+ scanchain_138/module_data_in[1] scanchain_138/module_data_in[2] scanchain_138/module_data_in[3]
+ scanchain_138/module_data_in[4] scanchain_138/module_data_in[5] scanchain_138/module_data_in[6]
+ scanchain_138/module_data_in[7] scanchain_138/module_data_out[0] scanchain_138/module_data_out[1]
+ scanchain_138/module_data_out[2] scanchain_138/module_data_out[3] scanchain_138/module_data_out[4]
+ scanchain_138/module_data_out[5] scanchain_138/module_data_out[6] scanchain_138/module_data_out[7]
+ scanchain_138/scan_select_in scanchain_139/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_152 scanchain_152/module_data_in[0] scanchain_152/module_data_in[1]
+ scanchain_152/module_data_in[2] scanchain_152/module_data_in[3] scanchain_152/module_data_in[4]
+ scanchain_152/module_data_in[5] scanchain_152/module_data_in[6] scanchain_152/module_data_in[7]
+ scanchain_152/module_data_out[0] scanchain_152/module_data_out[1] scanchain_152/module_data_out[2]
+ scanchain_152/module_data_out[3] scanchain_152/module_data_out[4] scanchain_152/module_data_out[5]
+ scanchain_152/module_data_out[6] scanchain_152/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_163 scanchain_163/module_data_in[0] scanchain_163/module_data_in[1]
+ scanchain_163/module_data_in[2] scanchain_163/module_data_in[3] scanchain_163/module_data_in[4]
+ scanchain_163/module_data_in[5] scanchain_163/module_data_in[6] scanchain_163/module_data_in[7]
+ scanchain_163/module_data_out[0] scanchain_163/module_data_out[1] scanchain_163/module_data_out[2]
+ scanchain_163/module_data_out[3] scanchain_163/module_data_out[4] scanchain_163/module_data_out[5]
+ scanchain_163/module_data_out[6] scanchain_163/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_185 scanchain_185/module_data_in[0] scanchain_185/module_data_in[1]
+ scanchain_185/module_data_in[2] scanchain_185/module_data_in[3] scanchain_185/module_data_in[4]
+ scanchain_185/module_data_in[5] scanchain_185/module_data_in[6] scanchain_185/module_data_in[7]
+ scanchain_185/module_data_out[0] scanchain_185/module_data_out[1] scanchain_185/module_data_out[2]
+ scanchain_185/module_data_out[3] scanchain_185/module_data_out[4] scanchain_185/module_data_out[5]
+ scanchain_185/module_data_out[6] scanchain_185/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_174 scanchain_174/module_data_in[0] scanchain_174/module_data_in[1]
+ scanchain_174/module_data_in[2] scanchain_174/module_data_in[3] scanchain_174/module_data_in[4]
+ scanchain_174/module_data_in[5] scanchain_174/module_data_in[6] scanchain_174/module_data_in[7]
+ scanchain_174/module_data_out[0] scanchain_174/module_data_out[1] scanchain_174/module_data_out[2]
+ scanchain_174/module_data_out[3] scanchain_174/module_data_out[4] scanchain_174/module_data_out[5]
+ scanchain_174/module_data_out[6] scanchain_174/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xtholin_avalonsemi_5401_14 scanchain_14/module_data_in[0] scanchain_14/module_data_in[1]
+ scanchain_14/module_data_in[2] scanchain_14/module_data_in[3] scanchain_14/module_data_in[4]
+ scanchain_14/module_data_in[5] scanchain_14/module_data_in[6] scanchain_14/module_data_in[7]
+ scanchain_14/module_data_out[0] scanchain_14/module_data_out[1] scanchain_14/module_data_out[2]
+ scanchain_14/module_data_out[3] scanchain_14/module_data_out[4] scanchain_14/module_data_out[5]
+ scanchain_14/module_data_out[6] scanchain_14/module_data_out[7] vccd1 vssd1 tholin_avalonsemi_5401
Xmm21_LEDMatrixTop_26 mm21_LEDMatrixTop_26/io_in[0] mm21_LEDMatrixTop_26/io_in[1]
+ mm21_LEDMatrixTop_26/io_in[2] mm21_LEDMatrixTop_26/io_in[3] mm21_LEDMatrixTop_26/io_in[4]
+ mm21_LEDMatrixTop_26/io_in[5] mm21_LEDMatrixTop_26/io_in[6] mm21_LEDMatrixTop_26/io_in[7]
+ mm21_LEDMatrixTop_26/io_out[0] mm21_LEDMatrixTop_26/io_out[1] mm21_LEDMatrixTop_26/io_out[2]
+ mm21_LEDMatrixTop_26/io_out[3] mm21_LEDMatrixTop_26/io_out[4] mm21_LEDMatrixTop_26/io_out[5]
+ mm21_LEDMatrixTop_26/io_out[6] mm21_LEDMatrixTop_26/io_out[7] vccd1 vssd1 mm21_LEDMatrixTop
Xuser_module_339501025136214612_345 scanchain_345/module_data_in[0] scanchain_345/module_data_in[1]
+ scanchain_345/module_data_in[2] scanchain_345/module_data_in[3] scanchain_345/module_data_in[4]
+ scanchain_345/module_data_in[5] scanchain_345/module_data_in[6] scanchain_345/module_data_in[7]
+ scanchain_345/module_data_out[0] scanchain_345/module_data_out[1] scanchain_345/module_data_out[2]
+ scanchain_345/module_data_out[3] scanchain_345/module_data_out[4] scanchain_345/module_data_out[5]
+ scanchain_345/module_data_out[6] scanchain_345/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_323 scanchain_323/module_data_in[0] scanchain_323/module_data_in[1]
+ scanchain_323/module_data_in[2] scanchain_323/module_data_in[3] scanchain_323/module_data_in[4]
+ scanchain_323/module_data_in[5] scanchain_323/module_data_in[6] scanchain_323/module_data_in[7]
+ scanchain_323/module_data_out[0] scanchain_323/module_data_out[1] scanchain_323/module_data_out[2]
+ scanchain_323/module_data_out[3] scanchain_323/module_data_out[4] scanchain_323/module_data_out[5]
+ scanchain_323/module_data_out[6] scanchain_323/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_334 scanchain_334/module_data_in[0] scanchain_334/module_data_in[1]
+ scanchain_334/module_data_in[2] scanchain_334/module_data_in[3] scanchain_334/module_data_in[4]
+ scanchain_334/module_data_in[5] scanchain_334/module_data_in[6] scanchain_334/module_data_in[7]
+ scanchain_334/module_data_out[0] scanchain_334/module_data_out[1] scanchain_334/module_data_out[2]
+ scanchain_334/module_data_out[3] scanchain_334/module_data_out[4] scanchain_334/module_data_out[5]
+ scanchain_334/module_data_out[6] scanchain_334/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_312 scanchain_312/module_data_in[0] scanchain_312/module_data_in[1]
+ scanchain_312/module_data_in[2] scanchain_312/module_data_in[3] scanchain_312/module_data_in[4]
+ scanchain_312/module_data_in[5] scanchain_312/module_data_in[6] scanchain_312/module_data_in[7]
+ scanchain_312/module_data_out[0] scanchain_312/module_data_out[1] scanchain_312/module_data_out[2]
+ scanchain_312/module_data_out[3] scanchain_312/module_data_out[4] scanchain_312/module_data_out[5]
+ scanchain_312/module_data_out[6] scanchain_312/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_301 scanchain_301/module_data_in[0] scanchain_301/module_data_in[1]
+ scanchain_301/module_data_in[2] scanchain_301/module_data_in[3] scanchain_301/module_data_in[4]
+ scanchain_301/module_data_in[5] scanchain_301/module_data_in[6] scanchain_301/module_data_in[7]
+ scanchain_301/module_data_out[0] scanchain_301/module_data_out[1] scanchain_301/module_data_out[2]
+ scanchain_301/module_data_out[3] scanchain_301/module_data_out[4] scanchain_301/module_data_out[5]
+ scanchain_301/module_data_out[6] scanchain_301/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_389 scanchain_389/module_data_in[0] scanchain_389/module_data_in[1]
+ scanchain_389/module_data_in[2] scanchain_389/module_data_in[3] scanchain_389/module_data_in[4]
+ scanchain_389/module_data_in[5] scanchain_389/module_data_in[6] scanchain_389/module_data_in[7]
+ scanchain_389/module_data_out[0] scanchain_389/module_data_out[1] scanchain_389/module_data_out[2]
+ scanchain_389/module_data_out[3] scanchain_389/module_data_out[4] scanchain_389/module_data_out[5]
+ scanchain_389/module_data_out[6] scanchain_389/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_378 scanchain_378/module_data_in[0] scanchain_378/module_data_in[1]
+ scanchain_378/module_data_in[2] scanchain_378/module_data_in[3] scanchain_378/module_data_in[4]
+ scanchain_378/module_data_in[5] scanchain_378/module_data_in[6] scanchain_378/module_data_in[7]
+ scanchain_378/module_data_out[0] scanchain_378/module_data_out[1] scanchain_378/module_data_out[2]
+ scanchain_378/module_data_out[3] scanchain_378/module_data_out[4] scanchain_378/module_data_out[5]
+ scanchain_378/module_data_out[6] scanchain_378/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_367 scanchain_367/module_data_in[0] scanchain_367/module_data_in[1]
+ scanchain_367/module_data_in[2] scanchain_367/module_data_in[3] scanchain_367/module_data_in[4]
+ scanchain_367/module_data_in[5] scanchain_367/module_data_in[6] scanchain_367/module_data_in[7]
+ scanchain_367/module_data_out[0] scanchain_367/module_data_out[1] scanchain_367/module_data_out[2]
+ scanchain_367/module_data_out[3] scanchain_367/module_data_out[4] scanchain_367/module_data_out[5]
+ scanchain_367/module_data_out[6] scanchain_367/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_356 scanchain_356/module_data_in[0] scanchain_356/module_data_in[1]
+ scanchain_356/module_data_in[2] scanchain_356/module_data_in[3] scanchain_356/module_data_in[4]
+ scanchain_356/module_data_in[5] scanchain_356/module_data_in[6] scanchain_356/module_data_in[7]
+ scanchain_356/module_data_out[0] scanchain_356/module_data_out[1] scanchain_356/module_data_out[2]
+ scanchain_356/module_data_out[3] scanchain_356/module_data_out[4] scanchain_356/module_data_out[5]
+ scanchain_356/module_data_out[6] scanchain_356/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_309 scanchain_309/clk_in scanchain_310/clk_in scanchain_309/data_in scanchain_310/data_in
+ scanchain_309/latch_enable_in scanchain_310/latch_enable_in scanchain_309/module_data_in[0]
+ scanchain_309/module_data_in[1] scanchain_309/module_data_in[2] scanchain_309/module_data_in[3]
+ scanchain_309/module_data_in[4] scanchain_309/module_data_in[5] scanchain_309/module_data_in[6]
+ scanchain_309/module_data_in[7] scanchain_309/module_data_out[0] scanchain_309/module_data_out[1]
+ scanchain_309/module_data_out[2] scanchain_309/module_data_out[3] scanchain_309/module_data_out[4]
+ scanchain_309/module_data_out[5] scanchain_309/module_data_out[6] scanchain_309/module_data_out[7]
+ scanchain_309/scan_select_in scanchain_310/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_197 scanchain_197/module_data_in[0] scanchain_197/module_data_in[1]
+ scanchain_197/module_data_in[2] scanchain_197/module_data_in[3] scanchain_197/module_data_in[4]
+ scanchain_197/module_data_in[5] scanchain_197/module_data_in[6] scanchain_197/module_data_in[7]
+ scanchain_197/module_data_out[0] scanchain_197/module_data_out[1] scanchain_197/module_data_out[2]
+ scanchain_197/module_data_out[3] scanchain_197/module_data_out[4] scanchain_197/module_data_out[5]
+ scanchain_197/module_data_out[6] scanchain_197/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_120 scanchain_120/module_data_in[0] scanchain_120/module_data_in[1]
+ scanchain_120/module_data_in[2] scanchain_120/module_data_in[3] scanchain_120/module_data_in[4]
+ scanchain_120/module_data_in[5] scanchain_120/module_data_in[6] scanchain_120/module_data_in[7]
+ scanchain_120/module_data_out[0] scanchain_120/module_data_out[1] scanchain_120/module_data_out[2]
+ scanchain_120/module_data_out[3] scanchain_120/module_data_out[4] scanchain_120/module_data_out[5]
+ scanchain_120/module_data_out[6] scanchain_120/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_142 scanchain_142/module_data_in[0] scanchain_142/module_data_in[1]
+ scanchain_142/module_data_in[2] scanchain_142/module_data_in[3] scanchain_142/module_data_in[4]
+ scanchain_142/module_data_in[5] scanchain_142/module_data_in[6] scanchain_142/module_data_in[7]
+ scanchain_142/module_data_out[0] scanchain_142/module_data_out[1] scanchain_142/module_data_out[2]
+ scanchain_142/module_data_out[3] scanchain_142/module_data_out[4] scanchain_142/module_data_out[5]
+ scanchain_142/module_data_out[6] scanchain_142/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_131 scanchain_131/module_data_in[0] scanchain_131/module_data_in[1]
+ scanchain_131/module_data_in[2] scanchain_131/module_data_in[3] scanchain_131/module_data_in[4]
+ scanchain_131/module_data_in[5] scanchain_131/module_data_in[6] scanchain_131/module_data_in[7]
+ scanchain_131/module_data_out[0] scanchain_131/module_data_out[1] scanchain_131/module_data_out[2]
+ scanchain_131/module_data_out[3] scanchain_131/module_data_out[4] scanchain_131/module_data_out[5]
+ scanchain_131/module_data_out[6] scanchain_131/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_153 scanchain_153/module_data_in[0] scanchain_153/module_data_in[1]
+ scanchain_153/module_data_in[2] scanchain_153/module_data_in[3] scanchain_153/module_data_in[4]
+ scanchain_153/module_data_in[5] scanchain_153/module_data_in[6] scanchain_153/module_data_in[7]
+ scanchain_153/module_data_out[0] scanchain_153/module_data_out[1] scanchain_153/module_data_out[2]
+ scanchain_153/module_data_out[3] scanchain_153/module_data_out[4] scanchain_153/module_data_out[5]
+ scanchain_153/module_data_out[6] scanchain_153/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_164 scanchain_164/module_data_in[0] scanchain_164/module_data_in[1]
+ scanchain_164/module_data_in[2] scanchain_164/module_data_in[3] scanchain_164/module_data_in[4]
+ scanchain_164/module_data_in[5] scanchain_164/module_data_in[6] scanchain_164/module_data_in[7]
+ scanchain_164/module_data_out[0] scanchain_164/module_data_out[1] scanchain_164/module_data_out[2]
+ scanchain_164/module_data_out[3] scanchain_164/module_data_out[4] scanchain_164/module_data_out[5]
+ scanchain_164/module_data_out[6] scanchain_164/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_186 scanchain_186/module_data_in[0] scanchain_186/module_data_in[1]
+ scanchain_186/module_data_in[2] scanchain_186/module_data_in[3] scanchain_186/module_data_in[4]
+ scanchain_186/module_data_in[5] scanchain_186/module_data_in[6] scanchain_186/module_data_in[7]
+ scanchain_186/module_data_out[0] scanchain_186/module_data_out[1] scanchain_186/module_data_out[2]
+ scanchain_186/module_data_out[3] scanchain_186/module_data_out[4] scanchain_186/module_data_out[5]
+ scanchain_186/module_data_out[6] scanchain_186/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_175 scanchain_175/module_data_in[0] scanchain_175/module_data_in[1]
+ scanchain_175/module_data_in[2] scanchain_175/module_data_in[3] scanchain_175/module_data_in[4]
+ scanchain_175/module_data_in[5] scanchain_175/module_data_in[6] scanchain_175/module_data_in[7]
+ scanchain_175/module_data_out[0] scanchain_175/module_data_out[1] scanchain_175/module_data_out[2]
+ scanchain_175/module_data_out[3] scanchain_175/module_data_out[4] scanchain_175/module_data_out[5]
+ scanchain_175/module_data_out[6] scanchain_175/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_106 scanchain_106/clk_in scanchain_107/clk_in scanchain_106/data_in scanchain_107/data_in
+ scanchain_106/latch_enable_in scanchain_107/latch_enable_in scanchain_106/module_data_in[0]
+ scanchain_106/module_data_in[1] scanchain_106/module_data_in[2] scanchain_106/module_data_in[3]
+ scanchain_106/module_data_in[4] scanchain_106/module_data_in[5] scanchain_106/module_data_in[6]
+ scanchain_106/module_data_in[7] scanchain_106/module_data_out[0] scanchain_106/module_data_out[1]
+ scanchain_106/module_data_out[2] scanchain_106/module_data_out[3] scanchain_106/module_data_out[4]
+ scanchain_106/module_data_out[5] scanchain_106/module_data_out[6] scanchain_106/module_data_out[7]
+ scanchain_106/scan_select_in scanchain_107/scan_select_in vccd1 vssd1 scanchain
Xscanchain_117 scanchain_117/clk_in scanchain_118/clk_in scanchain_117/data_in scanchain_118/data_in
+ scanchain_117/latch_enable_in scanchain_118/latch_enable_in scanchain_117/module_data_in[0]
+ scanchain_117/module_data_in[1] scanchain_117/module_data_in[2] scanchain_117/module_data_in[3]
+ scanchain_117/module_data_in[4] scanchain_117/module_data_in[5] scanchain_117/module_data_in[6]
+ scanchain_117/module_data_in[7] scanchain_117/module_data_out[0] scanchain_117/module_data_out[1]
+ scanchain_117/module_data_out[2] scanchain_117/module_data_out[3] scanchain_117/module_data_out[4]
+ scanchain_117/module_data_out[5] scanchain_117/module_data_out[6] scanchain_117/module_data_out[7]
+ scanchain_117/scan_select_in scanchain_118/scan_select_in vccd1 vssd1 scanchain
Xscanchain_128 scanchain_128/clk_in scanchain_129/clk_in scanchain_128/data_in scanchain_129/data_in
+ scanchain_128/latch_enable_in scanchain_129/latch_enable_in scanchain_128/module_data_in[0]
+ scanchain_128/module_data_in[1] scanchain_128/module_data_in[2] scanchain_128/module_data_in[3]
+ scanchain_128/module_data_in[4] scanchain_128/module_data_in[5] scanchain_128/module_data_in[6]
+ scanchain_128/module_data_in[7] scanchain_128/module_data_out[0] scanchain_128/module_data_out[1]
+ scanchain_128/module_data_out[2] scanchain_128/module_data_out[3] scanchain_128/module_data_out[4]
+ scanchain_128/module_data_out[5] scanchain_128/module_data_out[6] scanchain_128/module_data_out[7]
+ scanchain_128/scan_select_in scanchain_129/scan_select_in vccd1 vssd1 scanchain
Xscanchain_139 scanchain_139/clk_in scanchain_140/clk_in scanchain_139/data_in scanchain_140/data_in
+ scanchain_139/latch_enable_in scanchain_140/latch_enable_in scanchain_139/module_data_in[0]
+ scanchain_139/module_data_in[1] scanchain_139/module_data_in[2] scanchain_139/module_data_in[3]
+ scanchain_139/module_data_in[4] scanchain_139/module_data_in[5] scanchain_139/module_data_in[6]
+ scanchain_139/module_data_in[7] scanchain_139/module_data_out[0] scanchain_139/module_data_out[1]
+ scanchain_139/module_data_out[2] scanchain_139/module_data_out[3] scanchain_139/module_data_out[4]
+ scanchain_139/module_data_out[5] scanchain_139/module_data_out[6] scanchain_139/module_data_out[7]
+ scanchain_139/scan_select_in scanchain_140/scan_select_in vccd1 vssd1 scanchain
Xscanchain_470 scanchain_470/clk_in scanchain_471/clk_in scanchain_470/data_in scanchain_471/data_in
+ scanchain_470/latch_enable_in scanchain_471/latch_enable_in scanchain_470/module_data_in[0]
+ scanchain_470/module_data_in[1] scanchain_470/module_data_in[2] scanchain_470/module_data_in[3]
+ scanchain_470/module_data_in[4] scanchain_470/module_data_in[5] scanchain_470/module_data_in[6]
+ scanchain_470/module_data_in[7] scanchain_470/module_data_out[0] scanchain_470/module_data_out[1]
+ scanchain_470/module_data_out[2] scanchain_470/module_data_out[3] scanchain_470/module_data_out[4]
+ scanchain_470/module_data_out[5] scanchain_470/module_data_out[6] scanchain_470/module_data_out[7]
+ scanchain_470/scan_select_in scanchain_471/scan_select_in vccd1 vssd1 scanchain
Xuser_module_346553315158393428_16 scanchain_16/module_data_in[0] scanchain_16/module_data_in[1]
+ scanchain_16/module_data_in[2] scanchain_16/module_data_in[3] scanchain_16/module_data_in[4]
+ scanchain_16/module_data_in[5] scanchain_16/module_data_in[6] scanchain_16/module_data_in[7]
+ scanchain_16/module_data_out[0] scanchain_16/module_data_out[1] scanchain_16/module_data_out[2]
+ scanchain_16/module_data_out[3] scanchain_16/module_data_out[4] scanchain_16/module_data_out[5]
+ scanchain_16/module_data_out[6] scanchain_16/module_data_out[7] vccd1 vssd1 user_module_346553315158393428
Xuser_module_341541108650607187_47 scanchain_47/module_data_in[0] scanchain_47/module_data_in[1]
+ scanchain_47/module_data_in[2] scanchain_47/module_data_in[3] scanchain_47/module_data_in[4]
+ scanchain_47/module_data_in[5] scanchain_47/module_data_in[6] scanchain_47/module_data_in[7]
+ scanchain_47/module_data_out[0] scanchain_47/module_data_out[1] scanchain_47/module_data_out[2]
+ scanchain_47/module_data_out[3] scanchain_47/module_data_out[4] scanchain_47/module_data_out[5]
+ scanchain_47/module_data_out[6] scanchain_47/module_data_out[7] vccd1 vssd1 user_module_341541108650607187
Xuser_module_339501025136214612_379 scanchain_379/module_data_in[0] scanchain_379/module_data_in[1]
+ scanchain_379/module_data_in[2] scanchain_379/module_data_in[3] scanchain_379/module_data_in[4]
+ scanchain_379/module_data_in[5] scanchain_379/module_data_in[6] scanchain_379/module_data_in[7]
+ scanchain_379/module_data_out[0] scanchain_379/module_data_out[1] scanchain_379/module_data_out[2]
+ scanchain_379/module_data_out[3] scanchain_379/module_data_out[4] scanchain_379/module_data_out[5]
+ scanchain_379/module_data_out[6] scanchain_379/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_368 scanchain_368/module_data_in[0] scanchain_368/module_data_in[1]
+ scanchain_368/module_data_in[2] scanchain_368/module_data_in[3] scanchain_368/module_data_in[4]
+ scanchain_368/module_data_in[5] scanchain_368/module_data_in[6] scanchain_368/module_data_in[7]
+ scanchain_368/module_data_out[0] scanchain_368/module_data_out[1] scanchain_368/module_data_out[2]
+ scanchain_368/module_data_out[3] scanchain_368/module_data_out[4] scanchain_368/module_data_out[5]
+ scanchain_368/module_data_out[6] scanchain_368/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_357 scanchain_357/module_data_in[0] scanchain_357/module_data_in[1]
+ scanchain_357/module_data_in[2] scanchain_357/module_data_in[3] scanchain_357/module_data_in[4]
+ scanchain_357/module_data_in[5] scanchain_357/module_data_in[6] scanchain_357/module_data_in[7]
+ scanchain_357/module_data_out[0] scanchain_357/module_data_out[1] scanchain_357/module_data_out[2]
+ scanchain_357/module_data_out[3] scanchain_357/module_data_out[4] scanchain_357/module_data_out[5]
+ scanchain_357/module_data_out[6] scanchain_357/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_346 scanchain_346/module_data_in[0] scanchain_346/module_data_in[1]
+ scanchain_346/module_data_in[2] scanchain_346/module_data_in[3] scanchain_346/module_data_in[4]
+ scanchain_346/module_data_in[5] scanchain_346/module_data_in[6] scanchain_346/module_data_in[7]
+ scanchain_346/module_data_out[0] scanchain_346/module_data_out[1] scanchain_346/module_data_out[2]
+ scanchain_346/module_data_out[3] scanchain_346/module_data_out[4] scanchain_346/module_data_out[5]
+ scanchain_346/module_data_out[6] scanchain_346/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_324 scanchain_324/module_data_in[0] scanchain_324/module_data_in[1]
+ scanchain_324/module_data_in[2] scanchain_324/module_data_in[3] scanchain_324/module_data_in[4]
+ scanchain_324/module_data_in[5] scanchain_324/module_data_in[6] scanchain_324/module_data_in[7]
+ scanchain_324/module_data_out[0] scanchain_324/module_data_out[1] scanchain_324/module_data_out[2]
+ scanchain_324/module_data_out[3] scanchain_324/module_data_out[4] scanchain_324/module_data_out[5]
+ scanchain_324/module_data_out[6] scanchain_324/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_335 scanchain_335/module_data_in[0] scanchain_335/module_data_in[1]
+ scanchain_335/module_data_in[2] scanchain_335/module_data_in[3] scanchain_335/module_data_in[4]
+ scanchain_335/module_data_in[5] scanchain_335/module_data_in[6] scanchain_335/module_data_in[7]
+ scanchain_335/module_data_out[0] scanchain_335/module_data_out[1] scanchain_335/module_data_out[2]
+ scanchain_335/module_data_out[3] scanchain_335/module_data_out[4] scanchain_335/module_data_out[5]
+ scanchain_335/module_data_out[6] scanchain_335/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_313 scanchain_313/module_data_in[0] scanchain_313/module_data_in[1]
+ scanchain_313/module_data_in[2] scanchain_313/module_data_in[3] scanchain_313/module_data_in[4]
+ scanchain_313/module_data_in[5] scanchain_313/module_data_in[6] scanchain_313/module_data_in[7]
+ scanchain_313/module_data_out[0] scanchain_313/module_data_out[1] scanchain_313/module_data_out[2]
+ scanchain_313/module_data_out[3] scanchain_313/module_data_out[4] scanchain_313/module_data_out[5]
+ scanchain_313/module_data_out[6] scanchain_313/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_302 scanchain_302/module_data_in[0] scanchain_302/module_data_in[1]
+ scanchain_302/module_data_in[2] scanchain_302/module_data_in[3] scanchain_302/module_data_in[4]
+ scanchain_302/module_data_in[5] scanchain_302/module_data_in[6] scanchain_302/module_data_in[7]
+ scanchain_302/module_data_out[0] scanchain_302/module_data_out[1] scanchain_302/module_data_out[2]
+ scanchain_302/module_data_out[3] scanchain_302/module_data_out[4] scanchain_302/module_data_out[5]
+ scanchain_302/module_data_out[6] scanchain_302/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_198 scanchain_198/module_data_in[0] scanchain_198/module_data_in[1]
+ scanchain_198/module_data_in[2] scanchain_198/module_data_in[3] scanchain_198/module_data_in[4]
+ scanchain_198/module_data_in[5] scanchain_198/module_data_in[6] scanchain_198/module_data_in[7]
+ scanchain_198/module_data_out[0] scanchain_198/module_data_out[1] scanchain_198/module_data_out[2]
+ scanchain_198/module_data_out[3] scanchain_198/module_data_out[4] scanchain_198/module_data_out[5]
+ scanchain_198/module_data_out[6] scanchain_198/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_110 scanchain_110/module_data_in[0] scanchain_110/module_data_in[1]
+ scanchain_110/module_data_in[2] scanchain_110/module_data_in[3] scanchain_110/module_data_in[4]
+ scanchain_110/module_data_in[5] scanchain_110/module_data_in[6] scanchain_110/module_data_in[7]
+ scanchain_110/module_data_out[0] scanchain_110/module_data_out[1] scanchain_110/module_data_out[2]
+ scanchain_110/module_data_out[3] scanchain_110/module_data_out[4] scanchain_110/module_data_out[5]
+ scanchain_110/module_data_out[6] scanchain_110/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_121 scanchain_121/module_data_in[0] scanchain_121/module_data_in[1]
+ scanchain_121/module_data_in[2] scanchain_121/module_data_in[3] scanchain_121/module_data_in[4]
+ scanchain_121/module_data_in[5] scanchain_121/module_data_in[6] scanchain_121/module_data_in[7]
+ scanchain_121/module_data_out[0] scanchain_121/module_data_out[1] scanchain_121/module_data_out[2]
+ scanchain_121/module_data_out[3] scanchain_121/module_data_out[4] scanchain_121/module_data_out[5]
+ scanchain_121/module_data_out[6] scanchain_121/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_143 scanchain_143/module_data_in[0] scanchain_143/module_data_in[1]
+ scanchain_143/module_data_in[2] scanchain_143/module_data_in[3] scanchain_143/module_data_in[4]
+ scanchain_143/module_data_in[5] scanchain_143/module_data_in[6] scanchain_143/module_data_in[7]
+ scanchain_143/module_data_out[0] scanchain_143/module_data_out[1] scanchain_143/module_data_out[2]
+ scanchain_143/module_data_out[3] scanchain_143/module_data_out[4] scanchain_143/module_data_out[5]
+ scanchain_143/module_data_out[6] scanchain_143/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_132 scanchain_132/module_data_in[0] scanchain_132/module_data_in[1]
+ scanchain_132/module_data_in[2] scanchain_132/module_data_in[3] scanchain_132/module_data_in[4]
+ scanchain_132/module_data_in[5] scanchain_132/module_data_in[6] scanchain_132/module_data_in[7]
+ scanchain_132/module_data_out[0] scanchain_132/module_data_out[1] scanchain_132/module_data_out[2]
+ scanchain_132/module_data_out[3] scanchain_132/module_data_out[4] scanchain_132/module_data_out[5]
+ scanchain_132/module_data_out[6] scanchain_132/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_154 scanchain_154/module_data_in[0] scanchain_154/module_data_in[1]
+ scanchain_154/module_data_in[2] scanchain_154/module_data_in[3] scanchain_154/module_data_in[4]
+ scanchain_154/module_data_in[5] scanchain_154/module_data_in[6] scanchain_154/module_data_in[7]
+ scanchain_154/module_data_out[0] scanchain_154/module_data_out[1] scanchain_154/module_data_out[2]
+ scanchain_154/module_data_out[3] scanchain_154/module_data_out[4] scanchain_154/module_data_out[5]
+ scanchain_154/module_data_out[6] scanchain_154/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_165 scanchain_165/module_data_in[0] scanchain_165/module_data_in[1]
+ scanchain_165/module_data_in[2] scanchain_165/module_data_in[3] scanchain_165/module_data_in[4]
+ scanchain_165/module_data_in[5] scanchain_165/module_data_in[6] scanchain_165/module_data_in[7]
+ scanchain_165/module_data_out[0] scanchain_165/module_data_out[1] scanchain_165/module_data_out[2]
+ scanchain_165/module_data_out[3] scanchain_165/module_data_out[4] scanchain_165/module_data_out[5]
+ scanchain_165/module_data_out[6] scanchain_165/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_187 scanchain_187/module_data_in[0] scanchain_187/module_data_in[1]
+ scanchain_187/module_data_in[2] scanchain_187/module_data_in[3] scanchain_187/module_data_in[4]
+ scanchain_187/module_data_in[5] scanchain_187/module_data_in[6] scanchain_187/module_data_in[7]
+ scanchain_187/module_data_out[0] scanchain_187/module_data_out[1] scanchain_187/module_data_out[2]
+ scanchain_187/module_data_out[3] scanchain_187/module_data_out[4] scanchain_187/module_data_out[5]
+ scanchain_187/module_data_out[6] scanchain_187/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_176 scanchain_176/module_data_in[0] scanchain_176/module_data_in[1]
+ scanchain_176/module_data_in[2] scanchain_176/module_data_in[3] scanchain_176/module_data_in[4]
+ scanchain_176/module_data_in[5] scanchain_176/module_data_in[6] scanchain_176/module_data_in[7]
+ scanchain_176/module_data_out[0] scanchain_176/module_data_out[1] scanchain_176/module_data_out[2]
+ scanchain_176/module_data_out[3] scanchain_176/module_data_out[4] scanchain_176/module_data_out[5]
+ scanchain_176/module_data_out[6] scanchain_176/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_107 scanchain_107/clk_in scanchain_108/clk_in scanchain_107/data_in scanchain_108/data_in
+ scanchain_107/latch_enable_in scanchain_108/latch_enable_in scanchain_107/module_data_in[0]
+ scanchain_107/module_data_in[1] scanchain_107/module_data_in[2] scanchain_107/module_data_in[3]
+ scanchain_107/module_data_in[4] scanchain_107/module_data_in[5] scanchain_107/module_data_in[6]
+ scanchain_107/module_data_in[7] scanchain_107/module_data_out[0] scanchain_107/module_data_out[1]
+ scanchain_107/module_data_out[2] scanchain_107/module_data_out[3] scanchain_107/module_data_out[4]
+ scanchain_107/module_data_out[5] scanchain_107/module_data_out[6] scanchain_107/module_data_out[7]
+ scanchain_107/scan_select_in scanchain_108/scan_select_in vccd1 vssd1 scanchain
Xscanchain_118 scanchain_118/clk_in scanchain_119/clk_in scanchain_118/data_in scanchain_119/data_in
+ scanchain_118/latch_enable_in scanchain_119/latch_enable_in scanchain_118/module_data_in[0]
+ scanchain_118/module_data_in[1] scanchain_118/module_data_in[2] scanchain_118/module_data_in[3]
+ scanchain_118/module_data_in[4] scanchain_118/module_data_in[5] scanchain_118/module_data_in[6]
+ scanchain_118/module_data_in[7] scanchain_118/module_data_out[0] scanchain_118/module_data_out[1]
+ scanchain_118/module_data_out[2] scanchain_118/module_data_out[3] scanchain_118/module_data_out[4]
+ scanchain_118/module_data_out[5] scanchain_118/module_data_out[6] scanchain_118/module_data_out[7]
+ scanchain_118/scan_select_in scanchain_119/scan_select_in vccd1 vssd1 scanchain
Xscanchain_129 scanchain_129/clk_in scanchain_130/clk_in scanchain_129/data_in scanchain_130/data_in
+ scanchain_129/latch_enable_in scanchain_130/latch_enable_in scanchain_129/module_data_in[0]
+ scanchain_129/module_data_in[1] scanchain_129/module_data_in[2] scanchain_129/module_data_in[3]
+ scanchain_129/module_data_in[4] scanchain_129/module_data_in[5] scanchain_129/module_data_in[6]
+ scanchain_129/module_data_in[7] scanchain_129/module_data_out[0] scanchain_129/module_data_out[1]
+ scanchain_129/module_data_out[2] scanchain_129/module_data_out[3] scanchain_129/module_data_out[4]
+ scanchain_129/module_data_out[5] scanchain_129/module_data_out[6] scanchain_129/module_data_out[7]
+ scanchain_129/scan_select_in scanchain_130/scan_select_in vccd1 vssd1 scanchain
Xscanchain_471 scanchain_471/clk_in scanchain_472/clk_in scanchain_471/data_in scanchain_472/data_in
+ scanchain_471/latch_enable_in scanchain_472/latch_enable_in scanchain_471/module_data_in[0]
+ scanchain_471/module_data_in[1] scanchain_471/module_data_in[2] scanchain_471/module_data_in[3]
+ scanchain_471/module_data_in[4] scanchain_471/module_data_in[5] scanchain_471/module_data_in[6]
+ scanchain_471/module_data_in[7] scanchain_471/module_data_out[0] scanchain_471/module_data_out[1]
+ scanchain_471/module_data_out[2] scanchain_471/module_data_out[3] scanchain_471/module_data_out[4]
+ scanchain_471/module_data_out[5] scanchain_471/module_data_out[6] scanchain_471/module_data_out[7]
+ scanchain_471/scan_select_in scanchain_472/scan_select_in vccd1 vssd1 scanchain
Xscanchain_460 scanchain_460/clk_in scanchain_461/clk_in scanchain_460/data_in scanchain_461/data_in
+ scanchain_460/latch_enable_in scanchain_461/latch_enable_in scanchain_460/module_data_in[0]
+ scanchain_460/module_data_in[1] scanchain_460/module_data_in[2] scanchain_460/module_data_in[3]
+ scanchain_460/module_data_in[4] scanchain_460/module_data_in[5] scanchain_460/module_data_in[6]
+ scanchain_460/module_data_in[7] scanchain_460/module_data_out[0] scanchain_460/module_data_out[1]
+ scanchain_460/module_data_out[2] scanchain_460/module_data_out[3] scanchain_460/module_data_out[4]
+ scanchain_460/module_data_out[5] scanchain_460/module_data_out[6] scanchain_460/module_data_out[7]
+ scanchain_460/scan_select_in scanchain_461/scan_select_in vccd1 vssd1 scanchain
Xscanchain_290 scanchain_290/clk_in scanchain_291/clk_in scanchain_290/data_in scanchain_291/data_in
+ scanchain_290/latch_enable_in scanchain_291/latch_enable_in scanchain_290/module_data_in[0]
+ scanchain_290/module_data_in[1] scanchain_290/module_data_in[2] scanchain_290/module_data_in[3]
+ scanchain_290/module_data_in[4] scanchain_290/module_data_in[5] scanchain_290/module_data_in[6]
+ scanchain_290/module_data_in[7] scanchain_290/module_data_out[0] scanchain_290/module_data_out[1]
+ scanchain_290/module_data_out[2] scanchain_290/module_data_out[3] scanchain_290/module_data_out[4]
+ scanchain_290/module_data_out[5] scanchain_290/module_data_out[6] scanchain_290/module_data_out[7]
+ scanchain_290/scan_select_in scanchain_291/scan_select_in vccd1 vssd1 scanchain
Xscanchain_0 scanchain_0/clk_in scanchain_1/clk_in scanchain_0/data_in scanchain_1/data_in
+ scanchain_0/latch_enable_in scanchain_1/latch_enable_in scanchain_0/module_data_in[0]
+ scanchain_0/module_data_in[1] scanchain_0/module_data_in[2] scanchain_0/module_data_in[3]
+ scanchain_0/module_data_in[4] scanchain_0/module_data_in[5] scanchain_0/module_data_in[6]
+ scanchain_0/module_data_in[7] scanchain_0/module_data_out[0] scanchain_0/module_data_out[1]
+ scanchain_0/module_data_out[2] scanchain_0/module_data_out[3] scanchain_0/module_data_out[4]
+ scanchain_0/module_data_out[5] scanchain_0/module_data_out[6] scanchain_0/module_data_out[7]
+ scanchain_0/scan_select_in scanchain_1/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_369 scanchain_369/module_data_in[0] scanchain_369/module_data_in[1]
+ scanchain_369/module_data_in[2] scanchain_369/module_data_in[3] scanchain_369/module_data_in[4]
+ scanchain_369/module_data_in[5] scanchain_369/module_data_in[6] scanchain_369/module_data_in[7]
+ scanchain_369/module_data_out[0] scanchain_369/module_data_out[1] scanchain_369/module_data_out[2]
+ scanchain_369/module_data_out[3] scanchain_369/module_data_out[4] scanchain_369/module_data_out[5]
+ scanchain_369/module_data_out[6] scanchain_369/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_358 scanchain_358/module_data_in[0] scanchain_358/module_data_in[1]
+ scanchain_358/module_data_in[2] scanchain_358/module_data_in[3] scanchain_358/module_data_in[4]
+ scanchain_358/module_data_in[5] scanchain_358/module_data_in[6] scanchain_358/module_data_in[7]
+ scanchain_358/module_data_out[0] scanchain_358/module_data_out[1] scanchain_358/module_data_out[2]
+ scanchain_358/module_data_out[3] scanchain_358/module_data_out[4] scanchain_358/module_data_out[5]
+ scanchain_358/module_data_out[6] scanchain_358/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_347 scanchain_347/module_data_in[0] scanchain_347/module_data_in[1]
+ scanchain_347/module_data_in[2] scanchain_347/module_data_in[3] scanchain_347/module_data_in[4]
+ scanchain_347/module_data_in[5] scanchain_347/module_data_in[6] scanchain_347/module_data_in[7]
+ scanchain_347/module_data_out[0] scanchain_347/module_data_out[1] scanchain_347/module_data_out[2]
+ scanchain_347/module_data_out[3] scanchain_347/module_data_out[4] scanchain_347/module_data_out[5]
+ scanchain_347/module_data_out[6] scanchain_347/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_325 scanchain_325/module_data_in[0] scanchain_325/module_data_in[1]
+ scanchain_325/module_data_in[2] scanchain_325/module_data_in[3] scanchain_325/module_data_in[4]
+ scanchain_325/module_data_in[5] scanchain_325/module_data_in[6] scanchain_325/module_data_in[7]
+ scanchain_325/module_data_out[0] scanchain_325/module_data_out[1] scanchain_325/module_data_out[2]
+ scanchain_325/module_data_out[3] scanchain_325/module_data_out[4] scanchain_325/module_data_out[5]
+ scanchain_325/module_data_out[6] scanchain_325/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_336 scanchain_336/module_data_in[0] scanchain_336/module_data_in[1]
+ scanchain_336/module_data_in[2] scanchain_336/module_data_in[3] scanchain_336/module_data_in[4]
+ scanchain_336/module_data_in[5] scanchain_336/module_data_in[6] scanchain_336/module_data_in[7]
+ scanchain_336/module_data_out[0] scanchain_336/module_data_out[1] scanchain_336/module_data_out[2]
+ scanchain_336/module_data_out[3] scanchain_336/module_data_out[4] scanchain_336/module_data_out[5]
+ scanchain_336/module_data_out[6] scanchain_336/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_314 scanchain_314/module_data_in[0] scanchain_314/module_data_in[1]
+ scanchain_314/module_data_in[2] scanchain_314/module_data_in[3] scanchain_314/module_data_in[4]
+ scanchain_314/module_data_in[5] scanchain_314/module_data_in[6] scanchain_314/module_data_in[7]
+ scanchain_314/module_data_out[0] scanchain_314/module_data_out[1] scanchain_314/module_data_out[2]
+ scanchain_314/module_data_out[3] scanchain_314/module_data_out[4] scanchain_314/module_data_out[5]
+ scanchain_314/module_data_out[6] scanchain_314/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_303 scanchain_303/module_data_in[0] scanchain_303/module_data_in[1]
+ scanchain_303/module_data_in[2] scanchain_303/module_data_in[3] scanchain_303/module_data_in[4]
+ scanchain_303/module_data_in[5] scanchain_303/module_data_in[6] scanchain_303/module_data_in[7]
+ scanchain_303/module_data_out[0] scanchain_303/module_data_out[1] scanchain_303/module_data_out[2]
+ scanchain_303/module_data_out[3] scanchain_303/module_data_out[4] scanchain_303/module_data_out[5]
+ scanchain_303/module_data_out[6] scanchain_303/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_100 scanchain_100/module_data_in[0] scanchain_100/module_data_in[1]
+ scanchain_100/module_data_in[2] scanchain_100/module_data_in[3] scanchain_100/module_data_in[4]
+ scanchain_100/module_data_in[5] scanchain_100/module_data_in[6] scanchain_100/module_data_in[7]
+ scanchain_100/module_data_out[0] scanchain_100/module_data_out[1] scanchain_100/module_data_out[2]
+ scanchain_100/module_data_out[3] scanchain_100/module_data_out[4] scanchain_100/module_data_out[5]
+ scanchain_100/module_data_out[6] scanchain_100/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_199 scanchain_199/module_data_in[0] scanchain_199/module_data_in[1]
+ scanchain_199/module_data_in[2] scanchain_199/module_data_in[3] scanchain_199/module_data_in[4]
+ scanchain_199/module_data_in[5] scanchain_199/module_data_in[6] scanchain_199/module_data_in[7]
+ scanchain_199/module_data_out[0] scanchain_199/module_data_out[1] scanchain_199/module_data_out[2]
+ scanchain_199/module_data_out[3] scanchain_199/module_data_out[4] scanchain_199/module_data_out[5]
+ scanchain_199/module_data_out[6] scanchain_199/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_111 scanchain_111/module_data_in[0] scanchain_111/module_data_in[1]
+ scanchain_111/module_data_in[2] scanchain_111/module_data_in[3] scanchain_111/module_data_in[4]
+ scanchain_111/module_data_in[5] scanchain_111/module_data_in[6] scanchain_111/module_data_in[7]
+ scanchain_111/module_data_out[0] scanchain_111/module_data_out[1] scanchain_111/module_data_out[2]
+ scanchain_111/module_data_out[3] scanchain_111/module_data_out[4] scanchain_111/module_data_out[5]
+ scanchain_111/module_data_out[6] scanchain_111/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_108 scanchain_108/clk_in scanchain_109/clk_in scanchain_108/data_in scanchain_109/data_in
+ scanchain_108/latch_enable_in scanchain_109/latch_enable_in scanchain_108/module_data_in[0]
+ scanchain_108/module_data_in[1] scanchain_108/module_data_in[2] scanchain_108/module_data_in[3]
+ scanchain_108/module_data_in[4] scanchain_108/module_data_in[5] scanchain_108/module_data_in[6]
+ scanchain_108/module_data_in[7] scanchain_108/module_data_out[0] scanchain_108/module_data_out[1]
+ scanchain_108/module_data_out[2] scanchain_108/module_data_out[3] scanchain_108/module_data_out[4]
+ scanchain_108/module_data_out[5] scanchain_108/module_data_out[6] scanchain_108/module_data_out[7]
+ scanchain_108/scan_select_in scanchain_109/scan_select_in vccd1 vssd1 scanchain
Xscanchain_119 scanchain_119/clk_in scanchain_120/clk_in scanchain_119/data_in scanchain_120/data_in
+ scanchain_119/latch_enable_in scanchain_120/latch_enable_in scanchain_119/module_data_in[0]
+ scanchain_119/module_data_in[1] scanchain_119/module_data_in[2] scanchain_119/module_data_in[3]
+ scanchain_119/module_data_in[4] scanchain_119/module_data_in[5] scanchain_119/module_data_in[6]
+ scanchain_119/module_data_in[7] scanchain_119/module_data_out[0] scanchain_119/module_data_out[1]
+ scanchain_119/module_data_out[2] scanchain_119/module_data_out[3] scanchain_119/module_data_out[4]
+ scanchain_119/module_data_out[5] scanchain_119/module_data_out[6] scanchain_119/module_data_out[7]
+ scanchain_119/scan_select_in scanchain_120/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_122 scanchain_122/module_data_in[0] scanchain_122/module_data_in[1]
+ scanchain_122/module_data_in[2] scanchain_122/module_data_in[3] scanchain_122/module_data_in[4]
+ scanchain_122/module_data_in[5] scanchain_122/module_data_in[6] scanchain_122/module_data_in[7]
+ scanchain_122/module_data_out[0] scanchain_122/module_data_out[1] scanchain_122/module_data_out[2]
+ scanchain_122/module_data_out[3] scanchain_122/module_data_out[4] scanchain_122/module_data_out[5]
+ scanchain_122/module_data_out[6] scanchain_122/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_144 scanchain_144/module_data_in[0] scanchain_144/module_data_in[1]
+ scanchain_144/module_data_in[2] scanchain_144/module_data_in[3] scanchain_144/module_data_in[4]
+ scanchain_144/module_data_in[5] scanchain_144/module_data_in[6] scanchain_144/module_data_in[7]
+ scanchain_144/module_data_out[0] scanchain_144/module_data_out[1] scanchain_144/module_data_out[2]
+ scanchain_144/module_data_out[3] scanchain_144/module_data_out[4] scanchain_144/module_data_out[5]
+ scanchain_144/module_data_out[6] scanchain_144/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_133 scanchain_133/module_data_in[0] scanchain_133/module_data_in[1]
+ scanchain_133/module_data_in[2] scanchain_133/module_data_in[3] scanchain_133/module_data_in[4]
+ scanchain_133/module_data_in[5] scanchain_133/module_data_in[6] scanchain_133/module_data_in[7]
+ scanchain_133/module_data_out[0] scanchain_133/module_data_out[1] scanchain_133/module_data_out[2]
+ scanchain_133/module_data_out[3] scanchain_133/module_data_out[4] scanchain_133/module_data_out[5]
+ scanchain_133/module_data_out[6] scanchain_133/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_155 scanchain_155/module_data_in[0] scanchain_155/module_data_in[1]
+ scanchain_155/module_data_in[2] scanchain_155/module_data_in[3] scanchain_155/module_data_in[4]
+ scanchain_155/module_data_in[5] scanchain_155/module_data_in[6] scanchain_155/module_data_in[7]
+ scanchain_155/module_data_out[0] scanchain_155/module_data_out[1] scanchain_155/module_data_out[2]
+ scanchain_155/module_data_out[3] scanchain_155/module_data_out[4] scanchain_155/module_data_out[5]
+ scanchain_155/module_data_out[6] scanchain_155/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_166 scanchain_166/module_data_in[0] scanchain_166/module_data_in[1]
+ scanchain_166/module_data_in[2] scanchain_166/module_data_in[3] scanchain_166/module_data_in[4]
+ scanchain_166/module_data_in[5] scanchain_166/module_data_in[6] scanchain_166/module_data_in[7]
+ scanchain_166/module_data_out[0] scanchain_166/module_data_out[1] scanchain_166/module_data_out[2]
+ scanchain_166/module_data_out[3] scanchain_166/module_data_out[4] scanchain_166/module_data_out[5]
+ scanchain_166/module_data_out[6] scanchain_166/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_177 scanchain_177/module_data_in[0] scanchain_177/module_data_in[1]
+ scanchain_177/module_data_in[2] scanchain_177/module_data_in[3] scanchain_177/module_data_in[4]
+ scanchain_177/module_data_in[5] scanchain_177/module_data_in[6] scanchain_177/module_data_in[7]
+ scanchain_177/module_data_out[0] scanchain_177/module_data_out[1] scanchain_177/module_data_out[2]
+ scanchain_177/module_data_out[3] scanchain_177/module_data_out[4] scanchain_177/module_data_out[5]
+ scanchain_177/module_data_out[6] scanchain_177/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_188 scanchain_188/module_data_in[0] scanchain_188/module_data_in[1]
+ scanchain_188/module_data_in[2] scanchain_188/module_data_in[3] scanchain_188/module_data_in[4]
+ scanchain_188/module_data_in[5] scanchain_188/module_data_in[6] scanchain_188/module_data_in[7]
+ scanchain_188/module_data_out[0] scanchain_188/module_data_out[1] scanchain_188/module_data_out[2]
+ scanchain_188/module_data_out[3] scanchain_188/module_data_out[4] scanchain_188/module_data_out[5]
+ scanchain_188/module_data_out[6] scanchain_188/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xtholin_avalonsemi_tbb1143_24 scanchain_24/module_data_in[0] scanchain_24/module_data_in[1]
+ scanchain_24/module_data_in[2] scanchain_24/module_data_in[3] scanchain_24/module_data_in[4]
+ scanchain_24/module_data_in[5] scanchain_24/module_data_in[6] scanchain_24/module_data_in[7]
+ scanchain_24/module_data_out[0] scanchain_24/module_data_out[1] scanchain_24/module_data_out[2]
+ scanchain_24/module_data_out[3] scanchain_24/module_data_out[4] scanchain_24/module_data_out[5]
+ scanchain_24/module_data_out[6] scanchain_24/module_data_out[7] vccd1 vssd1 tholin_avalonsemi_tbb1143
Xscanchain_472 scanchain_472/clk_in scanchain_472/clk_out scanchain_472/data_in scanchain_472/data_out
+ scanchain_472/latch_enable_in scanchain_472/latch_enable_out scanchain_472/module_data_in[0]
+ scanchain_472/module_data_in[1] scanchain_472/module_data_in[2] scanchain_472/module_data_in[3]
+ scanchain_472/module_data_in[4] scanchain_472/module_data_in[5] scanchain_472/module_data_in[6]
+ scanchain_472/module_data_in[7] scanchain_472/module_data_out[0] scanchain_472/module_data_out[1]
+ scanchain_472/module_data_out[2] scanchain_472/module_data_out[3] scanchain_472/module_data_out[4]
+ scanchain_472/module_data_out[5] scanchain_472/module_data_out[6] scanchain_472/module_data_out[7]
+ scanchain_472/scan_select_in scanchain_472/scan_select_out vccd1 vssd1 scanchain
Xscanchain_461 scanchain_461/clk_in scanchain_462/clk_in scanchain_461/data_in scanchain_462/data_in
+ scanchain_461/latch_enable_in scanchain_462/latch_enable_in scanchain_461/module_data_in[0]
+ scanchain_461/module_data_in[1] scanchain_461/module_data_in[2] scanchain_461/module_data_in[3]
+ scanchain_461/module_data_in[4] scanchain_461/module_data_in[5] scanchain_461/module_data_in[6]
+ scanchain_461/module_data_in[7] scanchain_461/module_data_out[0] scanchain_461/module_data_out[1]
+ scanchain_461/module_data_out[2] scanchain_461/module_data_out[3] scanchain_461/module_data_out[4]
+ scanchain_461/module_data_out[5] scanchain_461/module_data_out[6] scanchain_461/module_data_out[7]
+ scanchain_461/scan_select_in scanchain_462/scan_select_in vccd1 vssd1 scanchain
Xscanchain_450 scanchain_450/clk_in scanchain_451/clk_in scanchain_450/data_in scanchain_451/data_in
+ scanchain_450/latch_enable_in scanchain_451/latch_enable_in scanchain_450/module_data_in[0]
+ scanchain_450/module_data_in[1] scanchain_450/module_data_in[2] scanchain_450/module_data_in[3]
+ scanchain_450/module_data_in[4] scanchain_450/module_data_in[5] scanchain_450/module_data_in[6]
+ scanchain_450/module_data_in[7] scanchain_450/module_data_out[0] scanchain_450/module_data_out[1]
+ scanchain_450/module_data_out[2] scanchain_450/module_data_out[3] scanchain_450/module_data_out[4]
+ scanchain_450/module_data_out[5] scanchain_450/module_data_out[6] scanchain_450/module_data_out[7]
+ scanchain_450/scan_select_in scanchain_451/scan_select_in vccd1 vssd1 scanchain
Xtomkeddie_top_tto_a_25 scanchain_25/module_data_in[0] scanchain_25/module_data_in[1]
+ scanchain_25/module_data_in[2] scanchain_25/module_data_in[3] scanchain_25/module_data_in[4]
+ scanchain_25/module_data_in[5] scanchain_25/module_data_in[6] scanchain_25/module_data_in[7]
+ scanchain_25/module_data_out[0] scanchain_25/module_data_out[1] scanchain_25/module_data_out[2]
+ scanchain_25/module_data_out[3] scanchain_25/module_data_out[4] scanchain_25/module_data_out[5]
+ scanchain_25/module_data_out[6] scanchain_25/module_data_out[7] vccd1 vssd1 tomkeddie_top_tto_a
Xscanchain_291 scanchain_291/clk_in scanchain_292/clk_in scanchain_291/data_in scanchain_292/data_in
+ scanchain_291/latch_enable_in scanchain_292/latch_enable_in scanchain_291/module_data_in[0]
+ scanchain_291/module_data_in[1] scanchain_291/module_data_in[2] scanchain_291/module_data_in[3]
+ scanchain_291/module_data_in[4] scanchain_291/module_data_in[5] scanchain_291/module_data_in[6]
+ scanchain_291/module_data_in[7] scanchain_291/module_data_out[0] scanchain_291/module_data_out[1]
+ scanchain_291/module_data_out[2] scanchain_291/module_data_out[3] scanchain_291/module_data_out[4]
+ scanchain_291/module_data_out[5] scanchain_291/module_data_out[6] scanchain_291/module_data_out[7]
+ scanchain_291/scan_select_in scanchain_292/scan_select_in vccd1 vssd1 scanchain
Xscanchain_280 scanchain_280/clk_in scanchain_281/clk_in scanchain_280/data_in scanchain_281/data_in
+ scanchain_280/latch_enable_in scanchain_281/latch_enable_in scanchain_280/module_data_in[0]
+ scanchain_280/module_data_in[1] scanchain_280/module_data_in[2] scanchain_280/module_data_in[3]
+ scanchain_280/module_data_in[4] scanchain_280/module_data_in[5] scanchain_280/module_data_in[6]
+ scanchain_280/module_data_in[7] scanchain_280/module_data_out[0] scanchain_280/module_data_out[1]
+ scanchain_280/module_data_out[2] scanchain_280/module_data_out[3] scanchain_280/module_data_out[4]
+ scanchain_280/module_data_out[5] scanchain_280/module_data_out[6] scanchain_280/module_data_out[7]
+ scanchain_280/scan_select_in scanchain_281/scan_select_in vccd1 vssd1 scanchain
Xscanchain_1 scanchain_1/clk_in scanchain_2/clk_in scanchain_1/data_in scanchain_2/data_in
+ scanchain_1/latch_enable_in scanchain_2/latch_enable_in fraserbc_simon_1/io_in[0]
+ fraserbc_simon_1/io_in[1] fraserbc_simon_1/io_in[2] fraserbc_simon_1/io_in[3] fraserbc_simon_1/io_in[4]
+ fraserbc_simon_1/io_in[5] fraserbc_simon_1/io_in[6] fraserbc_simon_1/io_in[7] fraserbc_simon_1/io_out[0]
+ fraserbc_simon_1/io_out[1] fraserbc_simon_1/io_out[2] fraserbc_simon_1/io_out[3]
+ fraserbc_simon_1/io_out[4] fraserbc_simon_1/io_out[5] fraserbc_simon_1/io_out[6]
+ fraserbc_simon_1/io_out[7] scanchain_1/scan_select_in scanchain_2/scan_select_in
+ vccd1 vssd1 scanchain
Xuser_module_339501025136214612_359 scanchain_359/module_data_in[0] scanchain_359/module_data_in[1]
+ scanchain_359/module_data_in[2] scanchain_359/module_data_in[3] scanchain_359/module_data_in[4]
+ scanchain_359/module_data_in[5] scanchain_359/module_data_in[6] scanchain_359/module_data_in[7]
+ scanchain_359/module_data_out[0] scanchain_359/module_data_out[1] scanchain_359/module_data_out[2]
+ scanchain_359/module_data_out[3] scanchain_359/module_data_out[4] scanchain_359/module_data_out[5]
+ scanchain_359/module_data_out[6] scanchain_359/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_348 scanchain_348/module_data_in[0] scanchain_348/module_data_in[1]
+ scanchain_348/module_data_in[2] scanchain_348/module_data_in[3] scanchain_348/module_data_in[4]
+ scanchain_348/module_data_in[5] scanchain_348/module_data_in[6] scanchain_348/module_data_in[7]
+ scanchain_348/module_data_out[0] scanchain_348/module_data_out[1] scanchain_348/module_data_out[2]
+ scanchain_348/module_data_out[3] scanchain_348/module_data_out[4] scanchain_348/module_data_out[5]
+ scanchain_348/module_data_out[6] scanchain_348/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_326 scanchain_326/module_data_in[0] scanchain_326/module_data_in[1]
+ scanchain_326/module_data_in[2] scanchain_326/module_data_in[3] scanchain_326/module_data_in[4]
+ scanchain_326/module_data_in[5] scanchain_326/module_data_in[6] scanchain_326/module_data_in[7]
+ scanchain_326/module_data_out[0] scanchain_326/module_data_out[1] scanchain_326/module_data_out[2]
+ scanchain_326/module_data_out[3] scanchain_326/module_data_out[4] scanchain_326/module_data_out[5]
+ scanchain_326/module_data_out[6] scanchain_326/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_337 scanchain_337/module_data_in[0] scanchain_337/module_data_in[1]
+ scanchain_337/module_data_in[2] scanchain_337/module_data_in[3] scanchain_337/module_data_in[4]
+ scanchain_337/module_data_in[5] scanchain_337/module_data_in[6] scanchain_337/module_data_in[7]
+ scanchain_337/module_data_out[0] scanchain_337/module_data_out[1] scanchain_337/module_data_out[2]
+ scanchain_337/module_data_out[3] scanchain_337/module_data_out[4] scanchain_337/module_data_out[5]
+ scanchain_337/module_data_out[6] scanchain_337/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_315 scanchain_315/module_data_in[0] scanchain_315/module_data_in[1]
+ scanchain_315/module_data_in[2] scanchain_315/module_data_in[3] scanchain_315/module_data_in[4]
+ scanchain_315/module_data_in[5] scanchain_315/module_data_in[6] scanchain_315/module_data_in[7]
+ scanchain_315/module_data_out[0] scanchain_315/module_data_out[1] scanchain_315/module_data_out[2]
+ scanchain_315/module_data_out[3] scanchain_315/module_data_out[4] scanchain_315/module_data_out[5]
+ scanchain_315/module_data_out[6] scanchain_315/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_304 scanchain_304/module_data_in[0] scanchain_304/module_data_in[1]
+ scanchain_304/module_data_in[2] scanchain_304/module_data_in[3] scanchain_304/module_data_in[4]
+ scanchain_304/module_data_in[5] scanchain_304/module_data_in[6] scanchain_304/module_data_in[7]
+ scanchain_304/module_data_out[0] scanchain_304/module_data_out[1] scanchain_304/module_data_out[2]
+ scanchain_304/module_data_out[3] scanchain_304/module_data_out[4] scanchain_304/module_data_out[5]
+ scanchain_304/module_data_out[6] scanchain_304/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_109 scanchain_109/clk_in scanchain_110/clk_in scanchain_109/data_in scanchain_110/data_in
+ scanchain_109/latch_enable_in scanchain_110/latch_enable_in scanchain_109/module_data_in[0]
+ scanchain_109/module_data_in[1] scanchain_109/module_data_in[2] scanchain_109/module_data_in[3]
+ scanchain_109/module_data_in[4] scanchain_109/module_data_in[5] scanchain_109/module_data_in[6]
+ scanchain_109/module_data_in[7] scanchain_109/module_data_out[0] scanchain_109/module_data_out[1]
+ scanchain_109/module_data_out[2] scanchain_109/module_data_out[3] scanchain_109/module_data_out[4]
+ scanchain_109/module_data_out[5] scanchain_109/module_data_out[6] scanchain_109/module_data_out[7]
+ scanchain_109/scan_select_in scanchain_110/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_101 scanchain_101/module_data_in[0] scanchain_101/module_data_in[1]
+ scanchain_101/module_data_in[2] scanchain_101/module_data_in[3] scanchain_101/module_data_in[4]
+ scanchain_101/module_data_in[5] scanchain_101/module_data_in[6] scanchain_101/module_data_in[7]
+ scanchain_101/module_data_out[0] scanchain_101/module_data_out[1] scanchain_101/module_data_out[2]
+ scanchain_101/module_data_out[3] scanchain_101/module_data_out[4] scanchain_101/module_data_out[5]
+ scanchain_101/module_data_out[6] scanchain_101/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_112 scanchain_112/module_data_in[0] scanchain_112/module_data_in[1]
+ scanchain_112/module_data_in[2] scanchain_112/module_data_in[3] scanchain_112/module_data_in[4]
+ scanchain_112/module_data_in[5] scanchain_112/module_data_in[6] scanchain_112/module_data_in[7]
+ scanchain_112/module_data_out[0] scanchain_112/module_data_out[1] scanchain_112/module_data_out[2]
+ scanchain_112/module_data_out[3] scanchain_112/module_data_out[4] scanchain_112/module_data_out[5]
+ scanchain_112/module_data_out[6] scanchain_112/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_123 scanchain_123/module_data_in[0] scanchain_123/module_data_in[1]
+ scanchain_123/module_data_in[2] scanchain_123/module_data_in[3] scanchain_123/module_data_in[4]
+ scanchain_123/module_data_in[5] scanchain_123/module_data_in[6] scanchain_123/module_data_in[7]
+ scanchain_123/module_data_out[0] scanchain_123/module_data_out[1] scanchain_123/module_data_out[2]
+ scanchain_123/module_data_out[3] scanchain_123/module_data_out[4] scanchain_123/module_data_out[5]
+ scanchain_123/module_data_out[6] scanchain_123/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_145 scanchain_145/module_data_in[0] scanchain_145/module_data_in[1]
+ scanchain_145/module_data_in[2] scanchain_145/module_data_in[3] scanchain_145/module_data_in[4]
+ scanchain_145/module_data_in[5] scanchain_145/module_data_in[6] scanchain_145/module_data_in[7]
+ scanchain_145/module_data_out[0] scanchain_145/module_data_out[1] scanchain_145/module_data_out[2]
+ scanchain_145/module_data_out[3] scanchain_145/module_data_out[4] scanchain_145/module_data_out[5]
+ scanchain_145/module_data_out[6] scanchain_145/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_134 scanchain_134/module_data_in[0] scanchain_134/module_data_in[1]
+ scanchain_134/module_data_in[2] scanchain_134/module_data_in[3] scanchain_134/module_data_in[4]
+ scanchain_134/module_data_in[5] scanchain_134/module_data_in[6] scanchain_134/module_data_in[7]
+ scanchain_134/module_data_out[0] scanchain_134/module_data_out[1] scanchain_134/module_data_out[2]
+ scanchain_134/module_data_out[3] scanchain_134/module_data_out[4] scanchain_134/module_data_out[5]
+ scanchain_134/module_data_out[6] scanchain_134/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_156 scanchain_156/module_data_in[0] scanchain_156/module_data_in[1]
+ scanchain_156/module_data_in[2] scanchain_156/module_data_in[3] scanchain_156/module_data_in[4]
+ scanchain_156/module_data_in[5] scanchain_156/module_data_in[6] scanchain_156/module_data_in[7]
+ scanchain_156/module_data_out[0] scanchain_156/module_data_out[1] scanchain_156/module_data_out[2]
+ scanchain_156/module_data_out[3] scanchain_156/module_data_out[4] scanchain_156/module_data_out[5]
+ scanchain_156/module_data_out[6] scanchain_156/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_167 scanchain_167/module_data_in[0] scanchain_167/module_data_in[1]
+ scanchain_167/module_data_in[2] scanchain_167/module_data_in[3] scanchain_167/module_data_in[4]
+ scanchain_167/module_data_in[5] scanchain_167/module_data_in[6] scanchain_167/module_data_in[7]
+ scanchain_167/module_data_out[0] scanchain_167/module_data_out[1] scanchain_167/module_data_out[2]
+ scanchain_167/module_data_out[3] scanchain_167/module_data_out[4] scanchain_167/module_data_out[5]
+ scanchain_167/module_data_out[6] scanchain_167/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_178 scanchain_178/module_data_in[0] scanchain_178/module_data_in[1]
+ scanchain_178/module_data_in[2] scanchain_178/module_data_in[3] scanchain_178/module_data_in[4]
+ scanchain_178/module_data_in[5] scanchain_178/module_data_in[6] scanchain_178/module_data_in[7]
+ scanchain_178/module_data_out[0] scanchain_178/module_data_out[1] scanchain_178/module_data_out[2]
+ scanchain_178/module_data_out[3] scanchain_178/module_data_out[4] scanchain_178/module_data_out[5]
+ scanchain_178/module_data_out[6] scanchain_178/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_189 scanchain_189/module_data_in[0] scanchain_189/module_data_in[1]
+ scanchain_189/module_data_in[2] scanchain_189/module_data_in[3] scanchain_189/module_data_in[4]
+ scanchain_189/module_data_in[5] scanchain_189/module_data_in[6] scanchain_189/module_data_in[7]
+ scanchain_189/module_data_out[0] scanchain_189/module_data_out[1] scanchain_189/module_data_out[2]
+ scanchain_189/module_data_out[3] scanchain_189/module_data_out[4] scanchain_189/module_data_out[5]
+ scanchain_189/module_data_out[6] scanchain_189/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_462 scanchain_462/clk_in scanchain_463/clk_in scanchain_462/data_in scanchain_463/data_in
+ scanchain_462/latch_enable_in scanchain_463/latch_enable_in scanchain_462/module_data_in[0]
+ scanchain_462/module_data_in[1] scanchain_462/module_data_in[2] scanchain_462/module_data_in[3]
+ scanchain_462/module_data_in[4] scanchain_462/module_data_in[5] scanchain_462/module_data_in[6]
+ scanchain_462/module_data_in[7] scanchain_462/module_data_out[0] scanchain_462/module_data_out[1]
+ scanchain_462/module_data_out[2] scanchain_462/module_data_out[3] scanchain_462/module_data_out[4]
+ scanchain_462/module_data_out[5] scanchain_462/module_data_out[6] scanchain_462/module_data_out[7]
+ scanchain_462/scan_select_in scanchain_463/scan_select_in vccd1 vssd1 scanchain
Xscanchain_440 scanchain_440/clk_in scanchain_441/clk_in scanchain_440/data_in scanchain_441/data_in
+ scanchain_440/latch_enable_in scanchain_441/latch_enable_in scanchain_440/module_data_in[0]
+ scanchain_440/module_data_in[1] scanchain_440/module_data_in[2] scanchain_440/module_data_in[3]
+ scanchain_440/module_data_in[4] scanchain_440/module_data_in[5] scanchain_440/module_data_in[6]
+ scanchain_440/module_data_in[7] scanchain_440/module_data_out[0] scanchain_440/module_data_out[1]
+ scanchain_440/module_data_out[2] scanchain_440/module_data_out[3] scanchain_440/module_data_out[4]
+ scanchain_440/module_data_out[5] scanchain_440/module_data_out[6] scanchain_440/module_data_out[7]
+ scanchain_440/scan_select_in scanchain_441/scan_select_in vccd1 vssd1 scanchain
Xscanchain_451 scanchain_451/clk_in scanchain_452/clk_in scanchain_451/data_in scanchain_452/data_in
+ scanchain_451/latch_enable_in scanchain_452/latch_enable_in scanchain_451/module_data_in[0]
+ scanchain_451/module_data_in[1] scanchain_451/module_data_in[2] scanchain_451/module_data_in[3]
+ scanchain_451/module_data_in[4] scanchain_451/module_data_in[5] scanchain_451/module_data_in[6]
+ scanchain_451/module_data_in[7] scanchain_451/module_data_out[0] scanchain_451/module_data_out[1]
+ scanchain_451/module_data_out[2] scanchain_451/module_data_out[3] scanchain_451/module_data_out[4]
+ scanchain_451/module_data_out[5] scanchain_451/module_data_out[6] scanchain_451/module_data_out[7]
+ scanchain_451/scan_select_in scanchain_452/scan_select_in vccd1 vssd1 scanchain
Xscanchain_270 scanchain_270/clk_in scanchain_271/clk_in scanchain_270/data_in scanchain_271/data_in
+ scanchain_270/latch_enable_in scanchain_271/latch_enable_in scanchain_270/module_data_in[0]
+ scanchain_270/module_data_in[1] scanchain_270/module_data_in[2] scanchain_270/module_data_in[3]
+ scanchain_270/module_data_in[4] scanchain_270/module_data_in[5] scanchain_270/module_data_in[6]
+ scanchain_270/module_data_in[7] scanchain_270/module_data_out[0] scanchain_270/module_data_out[1]
+ scanchain_270/module_data_out[2] scanchain_270/module_data_out[3] scanchain_270/module_data_out[4]
+ scanchain_270/module_data_out[5] scanchain_270/module_data_out[6] scanchain_270/module_data_out[7]
+ scanchain_270/scan_select_in scanchain_271/scan_select_in vccd1 vssd1 scanchain
Xscanchain_292 scanchain_292/clk_in scanchain_293/clk_in scanchain_292/data_in scanchain_293/data_in
+ scanchain_292/latch_enable_in scanchain_293/latch_enable_in scanchain_292/module_data_in[0]
+ scanchain_292/module_data_in[1] scanchain_292/module_data_in[2] scanchain_292/module_data_in[3]
+ scanchain_292/module_data_in[4] scanchain_292/module_data_in[5] scanchain_292/module_data_in[6]
+ scanchain_292/module_data_in[7] scanchain_292/module_data_out[0] scanchain_292/module_data_out[1]
+ scanchain_292/module_data_out[2] scanchain_292/module_data_out[3] scanchain_292/module_data_out[4]
+ scanchain_292/module_data_out[5] scanchain_292/module_data_out[6] scanchain_292/module_data_out[7]
+ scanchain_292/scan_select_in scanchain_293/scan_select_in vccd1 vssd1 scanchain
Xscanchain_281 scanchain_281/clk_in scanchain_282/clk_in scanchain_281/data_in scanchain_282/data_in
+ scanchain_281/latch_enable_in scanchain_282/latch_enable_in scanchain_281/module_data_in[0]
+ scanchain_281/module_data_in[1] scanchain_281/module_data_in[2] scanchain_281/module_data_in[3]
+ scanchain_281/module_data_in[4] scanchain_281/module_data_in[5] scanchain_281/module_data_in[6]
+ scanchain_281/module_data_in[7] scanchain_281/module_data_out[0] scanchain_281/module_data_out[1]
+ scanchain_281/module_data_out[2] scanchain_281/module_data_out[3] scanchain_281/module_data_out[4]
+ scanchain_281/module_data_out[5] scanchain_281/module_data_out[6] scanchain_281/module_data_out[7]
+ scanchain_281/scan_select_in scanchain_282/scan_select_in vccd1 vssd1 scanchain
Xscanchain_2 scanchain_2/clk_in scanchain_3/clk_in scanchain_2/data_in scanchain_3/data_in
+ scanchain_2/latch_enable_in scanchain_3/latch_enable_in tomkeddie_top_tto_2/io_in[0]
+ tomkeddie_top_tto_2/io_in[1] tomkeddie_top_tto_2/io_in[2] tomkeddie_top_tto_2/io_in[3]
+ tomkeddie_top_tto_2/io_in[4] tomkeddie_top_tto_2/io_in[5] tomkeddie_top_tto_2/io_in[6]
+ tomkeddie_top_tto_2/io_in[7] tomkeddie_top_tto_2/io_out[0] tomkeddie_top_tto_2/io_out[1]
+ tomkeddie_top_tto_2/io_out[2] tomkeddie_top_tto_2/io_out[3] tomkeddie_top_tto_2/io_out[4]
+ tomkeddie_top_tto_2/io_out[5] tomkeddie_top_tto_2/io_out[6] tomkeddie_top_tto_2/io_out[7]
+ scanchain_2/scan_select_in scanchain_3/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_349 scanchain_349/module_data_in[0] scanchain_349/module_data_in[1]
+ scanchain_349/module_data_in[2] scanchain_349/module_data_in[3] scanchain_349/module_data_in[4]
+ scanchain_349/module_data_in[5] scanchain_349/module_data_in[6] scanchain_349/module_data_in[7]
+ scanchain_349/module_data_out[0] scanchain_349/module_data_out[1] scanchain_349/module_data_out[2]
+ scanchain_349/module_data_out[3] scanchain_349/module_data_out[4] scanchain_349/module_data_out[5]
+ scanchain_349/module_data_out[6] scanchain_349/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_327 scanchain_327/module_data_in[0] scanchain_327/module_data_in[1]
+ scanchain_327/module_data_in[2] scanchain_327/module_data_in[3] scanchain_327/module_data_in[4]
+ scanchain_327/module_data_in[5] scanchain_327/module_data_in[6] scanchain_327/module_data_in[7]
+ scanchain_327/module_data_out[0] scanchain_327/module_data_out[1] scanchain_327/module_data_out[2]
+ scanchain_327/module_data_out[3] scanchain_327/module_data_out[4] scanchain_327/module_data_out[5]
+ scanchain_327/module_data_out[6] scanchain_327/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_338 scanchain_338/module_data_in[0] scanchain_338/module_data_in[1]
+ scanchain_338/module_data_in[2] scanchain_338/module_data_in[3] scanchain_338/module_data_in[4]
+ scanchain_338/module_data_in[5] scanchain_338/module_data_in[6] scanchain_338/module_data_in[7]
+ scanchain_338/module_data_out[0] scanchain_338/module_data_out[1] scanchain_338/module_data_out[2]
+ scanchain_338/module_data_out[3] scanchain_338/module_data_out[4] scanchain_338/module_data_out[5]
+ scanchain_338/module_data_out[6] scanchain_338/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_316 scanchain_316/module_data_in[0] scanchain_316/module_data_in[1]
+ scanchain_316/module_data_in[2] scanchain_316/module_data_in[3] scanchain_316/module_data_in[4]
+ scanchain_316/module_data_in[5] scanchain_316/module_data_in[6] scanchain_316/module_data_in[7]
+ scanchain_316/module_data_out[0] scanchain_316/module_data_out[1] scanchain_316/module_data_out[2]
+ scanchain_316/module_data_out[3] scanchain_316/module_data_out[4] scanchain_316/module_data_out[5]
+ scanchain_316/module_data_out[6] scanchain_316/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_305 scanchain_305/module_data_in[0] scanchain_305/module_data_in[1]
+ scanchain_305/module_data_in[2] scanchain_305/module_data_in[3] scanchain_305/module_data_in[4]
+ scanchain_305/module_data_in[5] scanchain_305/module_data_in[6] scanchain_305/module_data_in[7]
+ scanchain_305/module_data_out[0] scanchain_305/module_data_out[1] scanchain_305/module_data_out[2]
+ scanchain_305/module_data_out[3] scanchain_305/module_data_out[4] scanchain_305/module_data_out[5]
+ scanchain_305/module_data_out[6] scanchain_305/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xtop_42 top_42/io_in[0] top_42/io_in[1] top_42/io_in[2] top_42/io_in[3] top_42/io_in[4]
+ top_42/io_in[5] top_42/io_in[6] top_42/io_in[7] top_42/io_out[0] top_42/io_out[1]
+ top_42/io_out[2] top_42/io_out[3] top_42/io_out[4] top_42/io_out[5] top_42/io_out[6]
+ top_42/io_out[7] vccd1 vssd1 top
Xuser_module_339501025136214612_102 scanchain_102/module_data_in[0] scanchain_102/module_data_in[1]
+ scanchain_102/module_data_in[2] scanchain_102/module_data_in[3] scanchain_102/module_data_in[4]
+ scanchain_102/module_data_in[5] scanchain_102/module_data_in[6] scanchain_102/module_data_in[7]
+ scanchain_102/module_data_out[0] scanchain_102/module_data_out[1] scanchain_102/module_data_out[2]
+ scanchain_102/module_data_out[3] scanchain_102/module_data_out[4] scanchain_102/module_data_out[5]
+ scanchain_102/module_data_out[6] scanchain_102/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_113 scanchain_113/module_data_in[0] scanchain_113/module_data_in[1]
+ scanchain_113/module_data_in[2] scanchain_113/module_data_in[3] scanchain_113/module_data_in[4]
+ scanchain_113/module_data_in[5] scanchain_113/module_data_in[6] scanchain_113/module_data_in[7]
+ scanchain_113/module_data_out[0] scanchain_113/module_data_out[1] scanchain_113/module_data_out[2]
+ scanchain_113/module_data_out[3] scanchain_113/module_data_out[4] scanchain_113/module_data_out[5]
+ scanchain_113/module_data_out[6] scanchain_113/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_124 scanchain_124/module_data_in[0] scanchain_124/module_data_in[1]
+ scanchain_124/module_data_in[2] scanchain_124/module_data_in[3] scanchain_124/module_data_in[4]
+ scanchain_124/module_data_in[5] scanchain_124/module_data_in[6] scanchain_124/module_data_in[7]
+ scanchain_124/module_data_out[0] scanchain_124/module_data_out[1] scanchain_124/module_data_out[2]
+ scanchain_124/module_data_out[3] scanchain_124/module_data_out[4] scanchain_124/module_data_out[5]
+ scanchain_124/module_data_out[6] scanchain_124/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_146 scanchain_146/module_data_in[0] scanchain_146/module_data_in[1]
+ scanchain_146/module_data_in[2] scanchain_146/module_data_in[3] scanchain_146/module_data_in[4]
+ scanchain_146/module_data_in[5] scanchain_146/module_data_in[6] scanchain_146/module_data_in[7]
+ scanchain_146/module_data_out[0] scanchain_146/module_data_out[1] scanchain_146/module_data_out[2]
+ scanchain_146/module_data_out[3] scanchain_146/module_data_out[4] scanchain_146/module_data_out[5]
+ scanchain_146/module_data_out[6] scanchain_146/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_135 scanchain_135/module_data_in[0] scanchain_135/module_data_in[1]
+ scanchain_135/module_data_in[2] scanchain_135/module_data_in[3] scanchain_135/module_data_in[4]
+ scanchain_135/module_data_in[5] scanchain_135/module_data_in[6] scanchain_135/module_data_in[7]
+ scanchain_135/module_data_out[0] scanchain_135/module_data_out[1] scanchain_135/module_data_out[2]
+ scanchain_135/module_data_out[3] scanchain_135/module_data_out[4] scanchain_135/module_data_out[5]
+ scanchain_135/module_data_out[6] scanchain_135/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_157 scanchain_157/module_data_in[0] scanchain_157/module_data_in[1]
+ scanchain_157/module_data_in[2] scanchain_157/module_data_in[3] scanchain_157/module_data_in[4]
+ scanchain_157/module_data_in[5] scanchain_157/module_data_in[6] scanchain_157/module_data_in[7]
+ scanchain_157/module_data_out[0] scanchain_157/module_data_out[1] scanchain_157/module_data_out[2]
+ scanchain_157/module_data_out[3] scanchain_157/module_data_out[4] scanchain_157/module_data_out[5]
+ scanchain_157/module_data_out[6] scanchain_157/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_168 scanchain_168/module_data_in[0] scanchain_168/module_data_in[1]
+ scanchain_168/module_data_in[2] scanchain_168/module_data_in[3] scanchain_168/module_data_in[4]
+ scanchain_168/module_data_in[5] scanchain_168/module_data_in[6] scanchain_168/module_data_in[7]
+ scanchain_168/module_data_out[0] scanchain_168/module_data_out[1] scanchain_168/module_data_out[2]
+ scanchain_168/module_data_out[3] scanchain_168/module_data_out[4] scanchain_168/module_data_out[5]
+ scanchain_168/module_data_out[6] scanchain_168/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_179 scanchain_179/module_data_in[0] scanchain_179/module_data_in[1]
+ scanchain_179/module_data_in[2] scanchain_179/module_data_in[3] scanchain_179/module_data_in[4]
+ scanchain_179/module_data_in[5] scanchain_179/module_data_in[6] scanchain_179/module_data_in[7]
+ scanchain_179/module_data_out[0] scanchain_179/module_data_out[1] scanchain_179/module_data_out[2]
+ scanchain_179/module_data_out[3] scanchain_179/module_data_out[4] scanchain_179/module_data_out[5]
+ scanchain_179/module_data_out[6] scanchain_179/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_463 scanchain_463/clk_in scanchain_464/clk_in scanchain_463/data_in scanchain_464/data_in
+ scanchain_463/latch_enable_in scanchain_464/latch_enable_in scanchain_463/module_data_in[0]
+ scanchain_463/module_data_in[1] scanchain_463/module_data_in[2] scanchain_463/module_data_in[3]
+ scanchain_463/module_data_in[4] scanchain_463/module_data_in[5] scanchain_463/module_data_in[6]
+ scanchain_463/module_data_in[7] scanchain_463/module_data_out[0] scanchain_463/module_data_out[1]
+ scanchain_463/module_data_out[2] scanchain_463/module_data_out[3] scanchain_463/module_data_out[4]
+ scanchain_463/module_data_out[5] scanchain_463/module_data_out[6] scanchain_463/module_data_out[7]
+ scanchain_463/scan_select_in scanchain_464/scan_select_in vccd1 vssd1 scanchain
Xscanchain_441 scanchain_441/clk_in scanchain_442/clk_in scanchain_441/data_in scanchain_442/data_in
+ scanchain_441/latch_enable_in scanchain_442/latch_enable_in scanchain_441/module_data_in[0]
+ scanchain_441/module_data_in[1] scanchain_441/module_data_in[2] scanchain_441/module_data_in[3]
+ scanchain_441/module_data_in[4] scanchain_441/module_data_in[5] scanchain_441/module_data_in[6]
+ scanchain_441/module_data_in[7] scanchain_441/module_data_out[0] scanchain_441/module_data_out[1]
+ scanchain_441/module_data_out[2] scanchain_441/module_data_out[3] scanchain_441/module_data_out[4]
+ scanchain_441/module_data_out[5] scanchain_441/module_data_out[6] scanchain_441/module_data_out[7]
+ scanchain_441/scan_select_in scanchain_442/scan_select_in vccd1 vssd1 scanchain
Xscanchain_452 scanchain_452/clk_in scanchain_453/clk_in scanchain_452/data_in scanchain_453/data_in
+ scanchain_452/latch_enable_in scanchain_453/latch_enable_in scanchain_452/module_data_in[0]
+ scanchain_452/module_data_in[1] scanchain_452/module_data_in[2] scanchain_452/module_data_in[3]
+ scanchain_452/module_data_in[4] scanchain_452/module_data_in[5] scanchain_452/module_data_in[6]
+ scanchain_452/module_data_in[7] scanchain_452/module_data_out[0] scanchain_452/module_data_out[1]
+ scanchain_452/module_data_out[2] scanchain_452/module_data_out[3] scanchain_452/module_data_out[4]
+ scanchain_452/module_data_out[5] scanchain_452/module_data_out[6] scanchain_452/module_data_out[7]
+ scanchain_452/scan_select_in scanchain_453/scan_select_in vccd1 vssd1 scanchain
Xscanchain_430 scanchain_430/clk_in scanchain_431/clk_in scanchain_430/data_in scanchain_431/data_in
+ scanchain_430/latch_enable_in scanchain_431/latch_enable_in scanchain_430/module_data_in[0]
+ scanchain_430/module_data_in[1] scanchain_430/module_data_in[2] scanchain_430/module_data_in[3]
+ scanchain_430/module_data_in[4] scanchain_430/module_data_in[5] scanchain_430/module_data_in[6]
+ scanchain_430/module_data_in[7] scanchain_430/module_data_out[0] scanchain_430/module_data_out[1]
+ scanchain_430/module_data_out[2] scanchain_430/module_data_out[3] scanchain_430/module_data_out[4]
+ scanchain_430/module_data_out[5] scanchain_430/module_data_out[6] scanchain_430/module_data_out[7]
+ scanchain_430/scan_select_in scanchain_431/scan_select_in vccd1 vssd1 scanchain
Xscanchain_293 scanchain_293/clk_in scanchain_294/clk_in scanchain_293/data_in scanchain_294/data_in
+ scanchain_293/latch_enable_in scanchain_294/latch_enable_in scanchain_293/module_data_in[0]
+ scanchain_293/module_data_in[1] scanchain_293/module_data_in[2] scanchain_293/module_data_in[3]
+ scanchain_293/module_data_in[4] scanchain_293/module_data_in[5] scanchain_293/module_data_in[6]
+ scanchain_293/module_data_in[7] scanchain_293/module_data_out[0] scanchain_293/module_data_out[1]
+ scanchain_293/module_data_out[2] scanchain_293/module_data_out[3] scanchain_293/module_data_out[4]
+ scanchain_293/module_data_out[5] scanchain_293/module_data_out[6] scanchain_293/module_data_out[7]
+ scanchain_293/scan_select_in scanchain_294/scan_select_in vccd1 vssd1 scanchain
Xscanchain_282 scanchain_282/clk_in scanchain_283/clk_in scanchain_282/data_in scanchain_283/data_in
+ scanchain_282/latch_enable_in scanchain_283/latch_enable_in scanchain_282/module_data_in[0]
+ scanchain_282/module_data_in[1] scanchain_282/module_data_in[2] scanchain_282/module_data_in[3]
+ scanchain_282/module_data_in[4] scanchain_282/module_data_in[5] scanchain_282/module_data_in[6]
+ scanchain_282/module_data_in[7] scanchain_282/module_data_out[0] scanchain_282/module_data_out[1]
+ scanchain_282/module_data_out[2] scanchain_282/module_data_out[3] scanchain_282/module_data_out[4]
+ scanchain_282/module_data_out[5] scanchain_282/module_data_out[6] scanchain_282/module_data_out[7]
+ scanchain_282/scan_select_in scanchain_283/scan_select_in vccd1 vssd1 scanchain
Xscanchain_271 scanchain_271/clk_in scanchain_272/clk_in scanchain_271/data_in scanchain_272/data_in
+ scanchain_271/latch_enable_in scanchain_272/latch_enable_in scanchain_271/module_data_in[0]
+ scanchain_271/module_data_in[1] scanchain_271/module_data_in[2] scanchain_271/module_data_in[3]
+ scanchain_271/module_data_in[4] scanchain_271/module_data_in[5] scanchain_271/module_data_in[6]
+ scanchain_271/module_data_in[7] scanchain_271/module_data_out[0] scanchain_271/module_data_out[1]
+ scanchain_271/module_data_out[2] scanchain_271/module_data_out[3] scanchain_271/module_data_out[4]
+ scanchain_271/module_data_out[5] scanchain_271/module_data_out[6] scanchain_271/module_data_out[7]
+ scanchain_271/scan_select_in scanchain_272/scan_select_in vccd1 vssd1 scanchain
Xscanchain_260 scanchain_260/clk_in scanchain_261/clk_in scanchain_260/data_in scanchain_261/data_in
+ scanchain_260/latch_enable_in scanchain_261/latch_enable_in scanchain_260/module_data_in[0]
+ scanchain_260/module_data_in[1] scanchain_260/module_data_in[2] scanchain_260/module_data_in[3]
+ scanchain_260/module_data_in[4] scanchain_260/module_data_in[5] scanchain_260/module_data_in[6]
+ scanchain_260/module_data_in[7] scanchain_260/module_data_out[0] scanchain_260/module_data_out[1]
+ scanchain_260/module_data_out[2] scanchain_260/module_data_out[3] scanchain_260/module_data_out[4]
+ scanchain_260/module_data_out[5] scanchain_260/module_data_out[6] scanchain_260/module_data_out[7]
+ scanchain_260/scan_select_in scanchain_261/scan_select_in vccd1 vssd1 scanchain
Xscanchain_3 scanchain_3/clk_in scanchain_4/clk_in scanchain_3/data_in scanchain_4/data_in
+ scanchain_3/latch_enable_in scanchain_4/latch_enable_in chrisruk_matrix_3/io_in[0]
+ chrisruk_matrix_3/io_in[1] chrisruk_matrix_3/io_in[2] chrisruk_matrix_3/io_in[3]
+ chrisruk_matrix_3/io_in[4] chrisruk_matrix_3/io_in[5] chrisruk_matrix_3/io_in[6]
+ chrisruk_matrix_3/io_in[7] chrisruk_matrix_3/io_out[0] chrisruk_matrix_3/io_out[1]
+ chrisruk_matrix_3/io_out[2] chrisruk_matrix_3/io_out[3] chrisruk_matrix_3/io_out[4]
+ chrisruk_matrix_3/io_out[5] chrisruk_matrix_3/io_out[6] chrisruk_matrix_3/io_out[7]
+ scanchain_3/scan_select_in scanchain_4/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_328 scanchain_328/module_data_in[0] scanchain_328/module_data_in[1]
+ scanchain_328/module_data_in[2] scanchain_328/module_data_in[3] scanchain_328/module_data_in[4]
+ scanchain_328/module_data_in[5] scanchain_328/module_data_in[6] scanchain_328/module_data_in[7]
+ scanchain_328/module_data_out[0] scanchain_328/module_data_out[1] scanchain_328/module_data_out[2]
+ scanchain_328/module_data_out[3] scanchain_328/module_data_out[4] scanchain_328/module_data_out[5]
+ scanchain_328/module_data_out[6] scanchain_328/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_339 scanchain_339/module_data_in[0] scanchain_339/module_data_in[1]
+ scanchain_339/module_data_in[2] scanchain_339/module_data_in[3] scanchain_339/module_data_in[4]
+ scanchain_339/module_data_in[5] scanchain_339/module_data_in[6] scanchain_339/module_data_in[7]
+ scanchain_339/module_data_out[0] scanchain_339/module_data_out[1] scanchain_339/module_data_out[2]
+ scanchain_339/module_data_out[3] scanchain_339/module_data_out[4] scanchain_339/module_data_out[5]
+ scanchain_339/module_data_out[6] scanchain_339/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_317 scanchain_317/module_data_in[0] scanchain_317/module_data_in[1]
+ scanchain_317/module_data_in[2] scanchain_317/module_data_in[3] scanchain_317/module_data_in[4]
+ scanchain_317/module_data_in[5] scanchain_317/module_data_in[6] scanchain_317/module_data_in[7]
+ scanchain_317/module_data_out[0] scanchain_317/module_data_out[1] scanchain_317/module_data_out[2]
+ scanchain_317/module_data_out[3] scanchain_317/module_data_out[4] scanchain_317/module_data_out[5]
+ scanchain_317/module_data_out[6] scanchain_317/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_306 scanchain_306/module_data_in[0] scanchain_306/module_data_in[1]
+ scanchain_306/module_data_in[2] scanchain_306/module_data_in[3] scanchain_306/module_data_in[4]
+ scanchain_306/module_data_in[5] scanchain_306/module_data_in[6] scanchain_306/module_data_in[7]
+ scanchain_306/module_data_out[0] scanchain_306/module_data_out[1] scanchain_306/module_data_out[2]
+ scanchain_306/module_data_out[3] scanchain_306/module_data_out[4] scanchain_306/module_data_out[5]
+ scanchain_306/module_data_out[6] scanchain_306/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_348242239268323922_37 scanchain_37/module_data_in[0] scanchain_37/module_data_in[1]
+ scanchain_37/module_data_in[2] scanchain_37/module_data_in[3] scanchain_37/module_data_in[4]
+ scanchain_37/module_data_in[5] scanchain_37/module_data_in[6] scanchain_37/module_data_in[7]
+ scanchain_37/module_data_out[0] scanchain_37/module_data_out[1] scanchain_37/module_data_out[2]
+ scanchain_37/module_data_out[3] scanchain_37/module_data_out[4] scanchain_37/module_data_out[5]
+ scanchain_37/module_data_out[6] scanchain_37/module_data_out[7] vccd1 vssd1 user_module_348242239268323922
Xuser_module_339501025136214612_103 scanchain_103/module_data_in[0] scanchain_103/module_data_in[1]
+ scanchain_103/module_data_in[2] scanchain_103/module_data_in[3] scanchain_103/module_data_in[4]
+ scanchain_103/module_data_in[5] scanchain_103/module_data_in[6] scanchain_103/module_data_in[7]
+ scanchain_103/module_data_out[0] scanchain_103/module_data_out[1] scanchain_103/module_data_out[2]
+ scanchain_103/module_data_out[3] scanchain_103/module_data_out[4] scanchain_103/module_data_out[5]
+ scanchain_103/module_data_out[6] scanchain_103/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_114 scanchain_114/module_data_in[0] scanchain_114/module_data_in[1]
+ scanchain_114/module_data_in[2] scanchain_114/module_data_in[3] scanchain_114/module_data_in[4]
+ scanchain_114/module_data_in[5] scanchain_114/module_data_in[6] scanchain_114/module_data_in[7]
+ scanchain_114/module_data_out[0] scanchain_114/module_data_out[1] scanchain_114/module_data_out[2]
+ scanchain_114/module_data_out[3] scanchain_114/module_data_out[4] scanchain_114/module_data_out[5]
+ scanchain_114/module_data_out[6] scanchain_114/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_125 scanchain_125/module_data_in[0] scanchain_125/module_data_in[1]
+ scanchain_125/module_data_in[2] scanchain_125/module_data_in[3] scanchain_125/module_data_in[4]
+ scanchain_125/module_data_in[5] scanchain_125/module_data_in[6] scanchain_125/module_data_in[7]
+ scanchain_125/module_data_out[0] scanchain_125/module_data_out[1] scanchain_125/module_data_out[2]
+ scanchain_125/module_data_out[3] scanchain_125/module_data_out[4] scanchain_125/module_data_out[5]
+ scanchain_125/module_data_out[6] scanchain_125/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_147 scanchain_147/module_data_in[0] scanchain_147/module_data_in[1]
+ scanchain_147/module_data_in[2] scanchain_147/module_data_in[3] scanchain_147/module_data_in[4]
+ scanchain_147/module_data_in[5] scanchain_147/module_data_in[6] scanchain_147/module_data_in[7]
+ scanchain_147/module_data_out[0] scanchain_147/module_data_out[1] scanchain_147/module_data_out[2]
+ scanchain_147/module_data_out[3] scanchain_147/module_data_out[4] scanchain_147/module_data_out[5]
+ scanchain_147/module_data_out[6] scanchain_147/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_136 scanchain_136/module_data_in[0] scanchain_136/module_data_in[1]
+ scanchain_136/module_data_in[2] scanchain_136/module_data_in[3] scanchain_136/module_data_in[4]
+ scanchain_136/module_data_in[5] scanchain_136/module_data_in[6] scanchain_136/module_data_in[7]
+ scanchain_136/module_data_out[0] scanchain_136/module_data_out[1] scanchain_136/module_data_out[2]
+ scanchain_136/module_data_out[3] scanchain_136/module_data_out[4] scanchain_136/module_data_out[5]
+ scanchain_136/module_data_out[6] scanchain_136/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_158 scanchain_158/module_data_in[0] scanchain_158/module_data_in[1]
+ scanchain_158/module_data_in[2] scanchain_158/module_data_in[3] scanchain_158/module_data_in[4]
+ scanchain_158/module_data_in[5] scanchain_158/module_data_in[6] scanchain_158/module_data_in[7]
+ scanchain_158/module_data_out[0] scanchain_158/module_data_out[1] scanchain_158/module_data_out[2]
+ scanchain_158/module_data_out[3] scanchain_158/module_data_out[4] scanchain_158/module_data_out[5]
+ scanchain_158/module_data_out[6] scanchain_158/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_169 scanchain_169/module_data_in[0] scanchain_169/module_data_in[1]
+ scanchain_169/module_data_in[2] scanchain_169/module_data_in[3] scanchain_169/module_data_in[4]
+ scanchain_169/module_data_in[5] scanchain_169/module_data_in[6] scanchain_169/module_data_in[7]
+ scanchain_169/module_data_out[0] scanchain_169/module_data_out[1] scanchain_169/module_data_out[2]
+ scanchain_169/module_data_out[3] scanchain_169/module_data_out[4] scanchain_169/module_data_out[5]
+ scanchain_169/module_data_out[6] scanchain_169/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_464 scanchain_464/clk_in scanchain_465/clk_in scanchain_464/data_in scanchain_465/data_in
+ scanchain_464/latch_enable_in scanchain_465/latch_enable_in scanchain_464/module_data_in[0]
+ scanchain_464/module_data_in[1] scanchain_464/module_data_in[2] scanchain_464/module_data_in[3]
+ scanchain_464/module_data_in[4] scanchain_464/module_data_in[5] scanchain_464/module_data_in[6]
+ scanchain_464/module_data_in[7] scanchain_464/module_data_out[0] scanchain_464/module_data_out[1]
+ scanchain_464/module_data_out[2] scanchain_464/module_data_out[3] scanchain_464/module_data_out[4]
+ scanchain_464/module_data_out[5] scanchain_464/module_data_out[6] scanchain_464/module_data_out[7]
+ scanchain_464/scan_select_in scanchain_465/scan_select_in vccd1 vssd1 scanchain
Xscanchain_442 scanchain_442/clk_in scanchain_443/clk_in scanchain_442/data_in scanchain_443/data_in
+ scanchain_442/latch_enable_in scanchain_443/latch_enable_in scanchain_442/module_data_in[0]
+ scanchain_442/module_data_in[1] scanchain_442/module_data_in[2] scanchain_442/module_data_in[3]
+ scanchain_442/module_data_in[4] scanchain_442/module_data_in[5] scanchain_442/module_data_in[6]
+ scanchain_442/module_data_in[7] scanchain_442/module_data_out[0] scanchain_442/module_data_out[1]
+ scanchain_442/module_data_out[2] scanchain_442/module_data_out[3] scanchain_442/module_data_out[4]
+ scanchain_442/module_data_out[5] scanchain_442/module_data_out[6] scanchain_442/module_data_out[7]
+ scanchain_442/scan_select_in scanchain_443/scan_select_in vccd1 vssd1 scanchain
Xscanchain_453 scanchain_453/clk_in scanchain_454/clk_in scanchain_453/data_in scanchain_454/data_in
+ scanchain_453/latch_enable_in scanchain_454/latch_enable_in scanchain_453/module_data_in[0]
+ scanchain_453/module_data_in[1] scanchain_453/module_data_in[2] scanchain_453/module_data_in[3]
+ scanchain_453/module_data_in[4] scanchain_453/module_data_in[5] scanchain_453/module_data_in[6]
+ scanchain_453/module_data_in[7] scanchain_453/module_data_out[0] scanchain_453/module_data_out[1]
+ scanchain_453/module_data_out[2] scanchain_453/module_data_out[3] scanchain_453/module_data_out[4]
+ scanchain_453/module_data_out[5] scanchain_453/module_data_out[6] scanchain_453/module_data_out[7]
+ scanchain_453/scan_select_in scanchain_454/scan_select_in vccd1 vssd1 scanchain
Xscanchain_431 scanchain_431/clk_in scanchain_432/clk_in scanchain_431/data_in scanchain_432/data_in
+ scanchain_431/latch_enable_in scanchain_432/latch_enable_in scanchain_431/module_data_in[0]
+ scanchain_431/module_data_in[1] scanchain_431/module_data_in[2] scanchain_431/module_data_in[3]
+ scanchain_431/module_data_in[4] scanchain_431/module_data_in[5] scanchain_431/module_data_in[6]
+ scanchain_431/module_data_in[7] scanchain_431/module_data_out[0] scanchain_431/module_data_out[1]
+ scanchain_431/module_data_out[2] scanchain_431/module_data_out[3] scanchain_431/module_data_out[4]
+ scanchain_431/module_data_out[5] scanchain_431/module_data_out[6] scanchain_431/module_data_out[7]
+ scanchain_431/scan_select_in scanchain_432/scan_select_in vccd1 vssd1 scanchain
Xscanchain_420 scanchain_420/clk_in scanchain_421/clk_in scanchain_420/data_in scanchain_421/data_in
+ scanchain_420/latch_enable_in scanchain_421/latch_enable_in scanchain_420/module_data_in[0]
+ scanchain_420/module_data_in[1] scanchain_420/module_data_in[2] scanchain_420/module_data_in[3]
+ scanchain_420/module_data_in[4] scanchain_420/module_data_in[5] scanchain_420/module_data_in[6]
+ scanchain_420/module_data_in[7] scanchain_420/module_data_out[0] scanchain_420/module_data_out[1]
+ scanchain_420/module_data_out[2] scanchain_420/module_data_out[3] scanchain_420/module_data_out[4]
+ scanchain_420/module_data_out[5] scanchain_420/module_data_out[6] scanchain_420/module_data_out[7]
+ scanchain_420/scan_select_in scanchain_421/scan_select_in vccd1 vssd1 scanchain
Xscanchain_283 scanchain_283/clk_in scanchain_284/clk_in scanchain_283/data_in scanchain_284/data_in
+ scanchain_283/latch_enable_in scanchain_284/latch_enable_in scanchain_283/module_data_in[0]
+ scanchain_283/module_data_in[1] scanchain_283/module_data_in[2] scanchain_283/module_data_in[3]
+ scanchain_283/module_data_in[4] scanchain_283/module_data_in[5] scanchain_283/module_data_in[6]
+ scanchain_283/module_data_in[7] scanchain_283/module_data_out[0] scanchain_283/module_data_out[1]
+ scanchain_283/module_data_out[2] scanchain_283/module_data_out[3] scanchain_283/module_data_out[4]
+ scanchain_283/module_data_out[5] scanchain_283/module_data_out[6] scanchain_283/module_data_out[7]
+ scanchain_283/scan_select_in scanchain_284/scan_select_in vccd1 vssd1 scanchain
Xscanchain_294 scanchain_294/clk_in scanchain_295/clk_in scanchain_294/data_in scanchain_295/data_in
+ scanchain_294/latch_enable_in scanchain_295/latch_enable_in scanchain_294/module_data_in[0]
+ scanchain_294/module_data_in[1] scanchain_294/module_data_in[2] scanchain_294/module_data_in[3]
+ scanchain_294/module_data_in[4] scanchain_294/module_data_in[5] scanchain_294/module_data_in[6]
+ scanchain_294/module_data_in[7] scanchain_294/module_data_out[0] scanchain_294/module_data_out[1]
+ scanchain_294/module_data_out[2] scanchain_294/module_data_out[3] scanchain_294/module_data_out[4]
+ scanchain_294/module_data_out[5] scanchain_294/module_data_out[6] scanchain_294/module_data_out[7]
+ scanchain_294/scan_select_in scanchain_295/scan_select_in vccd1 vssd1 scanchain
Xscanchain_272 scanchain_272/clk_in scanchain_273/clk_in scanchain_272/data_in scanchain_273/data_in
+ scanchain_272/latch_enable_in scanchain_273/latch_enable_in scanchain_272/module_data_in[0]
+ scanchain_272/module_data_in[1] scanchain_272/module_data_in[2] scanchain_272/module_data_in[3]
+ scanchain_272/module_data_in[4] scanchain_272/module_data_in[5] scanchain_272/module_data_in[6]
+ scanchain_272/module_data_in[7] scanchain_272/module_data_out[0] scanchain_272/module_data_out[1]
+ scanchain_272/module_data_out[2] scanchain_272/module_data_out[3] scanchain_272/module_data_out[4]
+ scanchain_272/module_data_out[5] scanchain_272/module_data_out[6] scanchain_272/module_data_out[7]
+ scanchain_272/scan_select_in scanchain_273/scan_select_in vccd1 vssd1 scanchain
Xscanchain_250 scanchain_250/clk_in scanchain_251/clk_in scanchain_250/data_in scanchain_251/data_in
+ scanchain_250/latch_enable_in scanchain_251/latch_enable_in scanchain_250/module_data_in[0]
+ scanchain_250/module_data_in[1] scanchain_250/module_data_in[2] scanchain_250/module_data_in[3]
+ scanchain_250/module_data_in[4] scanchain_250/module_data_in[5] scanchain_250/module_data_in[6]
+ scanchain_250/module_data_in[7] scanchain_250/module_data_out[0] scanchain_250/module_data_out[1]
+ scanchain_250/module_data_out[2] scanchain_250/module_data_out[3] scanchain_250/module_data_out[4]
+ scanchain_250/module_data_out[5] scanchain_250/module_data_out[6] scanchain_250/module_data_out[7]
+ scanchain_250/scan_select_in scanchain_251/scan_select_in vccd1 vssd1 scanchain
Xscanchain_261 scanchain_261/clk_in scanchain_262/clk_in scanchain_261/data_in scanchain_262/data_in
+ scanchain_261/latch_enable_in scanchain_262/latch_enable_in scanchain_261/module_data_in[0]
+ scanchain_261/module_data_in[1] scanchain_261/module_data_in[2] scanchain_261/module_data_in[3]
+ scanchain_261/module_data_in[4] scanchain_261/module_data_in[5] scanchain_261/module_data_in[6]
+ scanchain_261/module_data_in[7] scanchain_261/module_data_out[0] scanchain_261/module_data_out[1]
+ scanchain_261/module_data_out[2] scanchain_261/module_data_out[3] scanchain_261/module_data_out[4]
+ scanchain_261/module_data_out[5] scanchain_261/module_data_out[6] scanchain_261/module_data_out[7]
+ scanchain_261/scan_select_in scanchain_262/scan_select_in vccd1 vssd1 scanchain
Xscanchain_4 scanchain_4/clk_in scanchain_5/clk_in scanchain_4/data_in scanchain_5/data_in
+ scanchain_4/latch_enable_in scanchain_5/latch_enable_in loxodes_sequencer_4/io_in[0]
+ loxodes_sequencer_4/io_in[1] loxodes_sequencer_4/io_in[2] loxodes_sequencer_4/io_in[3]
+ loxodes_sequencer_4/io_in[4] loxodes_sequencer_4/io_in[5] loxodes_sequencer_4/io_in[6]
+ loxodes_sequencer_4/io_in[7] loxodes_sequencer_4/io_out[0] loxodes_sequencer_4/io_out[1]
+ loxodes_sequencer_4/io_out[2] loxodes_sequencer_4/io_out[3] loxodes_sequencer_4/io_out[4]
+ loxodes_sequencer_4/io_out[5] loxodes_sequencer_4/io_out[6] loxodes_sequencer_4/io_out[7]
+ scanchain_4/scan_select_in scanchain_5/scan_select_in vccd1 vssd1 scanchain
Xmoyes0_top_module_39 moyes0_top_module_39/io_in[0] moyes0_top_module_39/io_in[1]
+ moyes0_top_module_39/io_in[2] moyes0_top_module_39/io_in[3] moyes0_top_module_39/io_in[4]
+ moyes0_top_module_39/io_in[5] moyes0_top_module_39/io_in[6] moyes0_top_module_39/io_in[7]
+ moyes0_top_module_39/io_out[0] moyes0_top_module_39/io_out[1] moyes0_top_module_39/io_out[2]
+ moyes0_top_module_39/io_out[3] moyes0_top_module_39/io_out[4] moyes0_top_module_39/io_out[5]
+ moyes0_top_module_39/io_out[6] moyes0_top_module_39/io_out[7] vccd1 vssd1 moyes0_top_module
Xuser_module_339501025136214612_329 scanchain_329/module_data_in[0] scanchain_329/module_data_in[1]
+ scanchain_329/module_data_in[2] scanchain_329/module_data_in[3] scanchain_329/module_data_in[4]
+ scanchain_329/module_data_in[5] scanchain_329/module_data_in[6] scanchain_329/module_data_in[7]
+ scanchain_329/module_data_out[0] scanchain_329/module_data_out[1] scanchain_329/module_data_out[2]
+ scanchain_329/module_data_out[3] scanchain_329/module_data_out[4] scanchain_329/module_data_out[5]
+ scanchain_329/module_data_out[6] scanchain_329/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_318 scanchain_318/module_data_in[0] scanchain_318/module_data_in[1]
+ scanchain_318/module_data_in[2] scanchain_318/module_data_in[3] scanchain_318/module_data_in[4]
+ scanchain_318/module_data_in[5] scanchain_318/module_data_in[6] scanchain_318/module_data_in[7]
+ scanchain_318/module_data_out[0] scanchain_318/module_data_out[1] scanchain_318/module_data_out[2]
+ scanchain_318/module_data_out[3] scanchain_318/module_data_out[4] scanchain_318/module_data_out[5]
+ scanchain_318/module_data_out[6] scanchain_318/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_307 scanchain_307/module_data_in[0] scanchain_307/module_data_in[1]
+ scanchain_307/module_data_in[2] scanchain_307/module_data_in[3] scanchain_307/module_data_in[4]
+ scanchain_307/module_data_in[5] scanchain_307/module_data_in[6] scanchain_307/module_data_in[7]
+ scanchain_307/module_data_out[0] scanchain_307/module_data_out[1] scanchain_307/module_data_out[2]
+ scanchain_307/module_data_out[3] scanchain_307/module_data_out[4] scanchain_307/module_data_out[5]
+ scanchain_307/module_data_out[6] scanchain_307/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_104 scanchain_104/module_data_in[0] scanchain_104/module_data_in[1]
+ scanchain_104/module_data_in[2] scanchain_104/module_data_in[3] scanchain_104/module_data_in[4]
+ scanchain_104/module_data_in[5] scanchain_104/module_data_in[6] scanchain_104/module_data_in[7]
+ scanchain_104/module_data_out[0] scanchain_104/module_data_out[1] scanchain_104/module_data_out[2]
+ scanchain_104/module_data_out[3] scanchain_104/module_data_out[4] scanchain_104/module_data_out[5]
+ scanchain_104/module_data_out[6] scanchain_104/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_115 scanchain_115/module_data_in[0] scanchain_115/module_data_in[1]
+ scanchain_115/module_data_in[2] scanchain_115/module_data_in[3] scanchain_115/module_data_in[4]
+ scanchain_115/module_data_in[5] scanchain_115/module_data_in[6] scanchain_115/module_data_in[7]
+ scanchain_115/module_data_out[0] scanchain_115/module_data_out[1] scanchain_115/module_data_out[2]
+ scanchain_115/module_data_out[3] scanchain_115/module_data_out[4] scanchain_115/module_data_out[5]
+ scanchain_115/module_data_out[6] scanchain_115/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_126 scanchain_126/module_data_in[0] scanchain_126/module_data_in[1]
+ scanchain_126/module_data_in[2] scanchain_126/module_data_in[3] scanchain_126/module_data_in[4]
+ scanchain_126/module_data_in[5] scanchain_126/module_data_in[6] scanchain_126/module_data_in[7]
+ scanchain_126/module_data_out[0] scanchain_126/module_data_out[1] scanchain_126/module_data_out[2]
+ scanchain_126/module_data_out[3] scanchain_126/module_data_out[4] scanchain_126/module_data_out[5]
+ scanchain_126/module_data_out[6] scanchain_126/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_148 scanchain_148/module_data_in[0] scanchain_148/module_data_in[1]
+ scanchain_148/module_data_in[2] scanchain_148/module_data_in[3] scanchain_148/module_data_in[4]
+ scanchain_148/module_data_in[5] scanchain_148/module_data_in[6] scanchain_148/module_data_in[7]
+ scanchain_148/module_data_out[0] scanchain_148/module_data_out[1] scanchain_148/module_data_out[2]
+ scanchain_148/module_data_out[3] scanchain_148/module_data_out[4] scanchain_148/module_data_out[5]
+ scanchain_148/module_data_out[6] scanchain_148/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_137 scanchain_137/module_data_in[0] scanchain_137/module_data_in[1]
+ scanchain_137/module_data_in[2] scanchain_137/module_data_in[3] scanchain_137/module_data_in[4]
+ scanchain_137/module_data_in[5] scanchain_137/module_data_in[6] scanchain_137/module_data_in[7]
+ scanchain_137/module_data_out[0] scanchain_137/module_data_out[1] scanchain_137/module_data_out[2]
+ scanchain_137/module_data_out[3] scanchain_137/module_data_out[4] scanchain_137/module_data_out[5]
+ scanchain_137/module_data_out[6] scanchain_137/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_159 scanchain_159/module_data_in[0] scanchain_159/module_data_in[1]
+ scanchain_159/module_data_in[2] scanchain_159/module_data_in[3] scanchain_159/module_data_in[4]
+ scanchain_159/module_data_in[5] scanchain_159/module_data_in[6] scanchain_159/module_data_in[7]
+ scanchain_159/module_data_out[0] scanchain_159/module_data_out[1] scanchain_159/module_data_out[2]
+ scanchain_159/module_data_out[3] scanchain_159/module_data_out[4] scanchain_159/module_data_out[5]
+ scanchain_159/module_data_out[6] scanchain_159/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xflygoat_tt02_play_tune_53 scanchain_53/module_data_in[0] scanchain_53/module_data_in[1]
+ scanchain_53/module_data_in[2] scanchain_53/module_data_in[3] scanchain_53/module_data_in[4]
+ scanchain_53/module_data_in[5] scanchain_53/module_data_in[6] scanchain_53/module_data_in[7]
+ scanchain_53/module_data_out[0] scanchain_53/module_data_out[1] scanchain_53/module_data_out[2]
+ scanchain_53/module_data_out[3] scanchain_53/module_data_out[4] scanchain_53/module_data_out[5]
+ scanchain_53/module_data_out[6] scanchain_53/module_data_out[7] vccd1 vssd1 flygoat_tt02_play_tune
Xuser_module_348260124451668562_34 scanchain_34/module_data_in[0] scanchain_34/module_data_in[1]
+ scanchain_34/module_data_in[2] scanchain_34/module_data_in[3] scanchain_34/module_data_in[4]
+ scanchain_34/module_data_in[5] scanchain_34/module_data_in[6] scanchain_34/module_data_in[7]
+ scanchain_34/module_data_out[0] scanchain_34/module_data_out[1] scanchain_34/module_data_out[2]
+ scanchain_34/module_data_out[3] scanchain_34/module_data_out[4] scanchain_34/module_data_out[5]
+ scanchain_34/module_data_out[6] scanchain_34/module_data_out[7] vccd1 vssd1 user_module_348260124451668562
Xscanchain_465 scanchain_465/clk_in scanchain_466/clk_in scanchain_465/data_in scanchain_466/data_in
+ scanchain_465/latch_enable_in scanchain_466/latch_enable_in scanchain_465/module_data_in[0]
+ scanchain_465/module_data_in[1] scanchain_465/module_data_in[2] scanchain_465/module_data_in[3]
+ scanchain_465/module_data_in[4] scanchain_465/module_data_in[5] scanchain_465/module_data_in[6]
+ scanchain_465/module_data_in[7] scanchain_465/module_data_out[0] scanchain_465/module_data_out[1]
+ scanchain_465/module_data_out[2] scanchain_465/module_data_out[3] scanchain_465/module_data_out[4]
+ scanchain_465/module_data_out[5] scanchain_465/module_data_out[6] scanchain_465/module_data_out[7]
+ scanchain_465/scan_select_in scanchain_466/scan_select_in vccd1 vssd1 scanchain
Xscanchain_454 scanchain_454/clk_in scanchain_455/clk_in scanchain_454/data_in scanchain_455/data_in
+ scanchain_454/latch_enable_in scanchain_455/latch_enable_in scanchain_454/module_data_in[0]
+ scanchain_454/module_data_in[1] scanchain_454/module_data_in[2] scanchain_454/module_data_in[3]
+ scanchain_454/module_data_in[4] scanchain_454/module_data_in[5] scanchain_454/module_data_in[6]
+ scanchain_454/module_data_in[7] scanchain_454/module_data_out[0] scanchain_454/module_data_out[1]
+ scanchain_454/module_data_out[2] scanchain_454/module_data_out[3] scanchain_454/module_data_out[4]
+ scanchain_454/module_data_out[5] scanchain_454/module_data_out[6] scanchain_454/module_data_out[7]
+ scanchain_454/scan_select_in scanchain_455/scan_select_in vccd1 vssd1 scanchain
Xscanchain_443 scanchain_443/clk_in scanchain_444/clk_in scanchain_443/data_in scanchain_444/data_in
+ scanchain_443/latch_enable_in scanchain_444/latch_enable_in scanchain_443/module_data_in[0]
+ scanchain_443/module_data_in[1] scanchain_443/module_data_in[2] scanchain_443/module_data_in[3]
+ scanchain_443/module_data_in[4] scanchain_443/module_data_in[5] scanchain_443/module_data_in[6]
+ scanchain_443/module_data_in[7] scanchain_443/module_data_out[0] scanchain_443/module_data_out[1]
+ scanchain_443/module_data_out[2] scanchain_443/module_data_out[3] scanchain_443/module_data_out[4]
+ scanchain_443/module_data_out[5] scanchain_443/module_data_out[6] scanchain_443/module_data_out[7]
+ scanchain_443/scan_select_in scanchain_444/scan_select_in vccd1 vssd1 scanchain
Xscanchain_432 scanchain_432/clk_in scanchain_433/clk_in scanchain_432/data_in scanchain_433/data_in
+ scanchain_432/latch_enable_in scanchain_433/latch_enable_in scanchain_432/module_data_in[0]
+ scanchain_432/module_data_in[1] scanchain_432/module_data_in[2] scanchain_432/module_data_in[3]
+ scanchain_432/module_data_in[4] scanchain_432/module_data_in[5] scanchain_432/module_data_in[6]
+ scanchain_432/module_data_in[7] scanchain_432/module_data_out[0] scanchain_432/module_data_out[1]
+ scanchain_432/module_data_out[2] scanchain_432/module_data_out[3] scanchain_432/module_data_out[4]
+ scanchain_432/module_data_out[5] scanchain_432/module_data_out[6] scanchain_432/module_data_out[7]
+ scanchain_432/scan_select_in scanchain_433/scan_select_in vccd1 vssd1 scanchain
Xscanchain_421 scanchain_421/clk_in scanchain_422/clk_in scanchain_421/data_in scanchain_422/data_in
+ scanchain_421/latch_enable_in scanchain_422/latch_enable_in scanchain_421/module_data_in[0]
+ scanchain_421/module_data_in[1] scanchain_421/module_data_in[2] scanchain_421/module_data_in[3]
+ scanchain_421/module_data_in[4] scanchain_421/module_data_in[5] scanchain_421/module_data_in[6]
+ scanchain_421/module_data_in[7] scanchain_421/module_data_out[0] scanchain_421/module_data_out[1]
+ scanchain_421/module_data_out[2] scanchain_421/module_data_out[3] scanchain_421/module_data_out[4]
+ scanchain_421/module_data_out[5] scanchain_421/module_data_out[6] scanchain_421/module_data_out[7]
+ scanchain_421/scan_select_in scanchain_422/scan_select_in vccd1 vssd1 scanchain
Xscanchain_410 scanchain_410/clk_in scanchain_411/clk_in scanchain_410/data_in scanchain_411/data_in
+ scanchain_410/latch_enable_in scanchain_411/latch_enable_in scanchain_410/module_data_in[0]
+ scanchain_410/module_data_in[1] scanchain_410/module_data_in[2] scanchain_410/module_data_in[3]
+ scanchain_410/module_data_in[4] scanchain_410/module_data_in[5] scanchain_410/module_data_in[6]
+ scanchain_410/module_data_in[7] scanchain_410/module_data_out[0] scanchain_410/module_data_out[1]
+ scanchain_410/module_data_out[2] scanchain_410/module_data_out[3] scanchain_410/module_data_out[4]
+ scanchain_410/module_data_out[5] scanchain_410/module_data_out[6] scanchain_410/module_data_out[7]
+ scanchain_410/scan_select_in scanchain_411/scan_select_in vccd1 vssd1 scanchain
Xtiny_fft_15 tiny_fft_15/io_in[0] tiny_fft_15/io_in[1] tiny_fft_15/io_in[2] tiny_fft_15/io_in[3]
+ tiny_fft_15/io_in[4] tiny_fft_15/io_in[5] tiny_fft_15/io_in[6] tiny_fft_15/io_in[7]
+ tiny_fft_15/io_out[0] tiny_fft_15/io_out[1] tiny_fft_15/io_out[2] tiny_fft_15/io_out[3]
+ tiny_fft_15/io_out[4] tiny_fft_15/io_out[5] tiny_fft_15/io_out[6] tiny_fft_15/io_out[7]
+ vccd1 vssd1 tiny_fft
Xscanchain_284 scanchain_284/clk_in scanchain_285/clk_in scanchain_284/data_in scanchain_285/data_in
+ scanchain_284/latch_enable_in scanchain_285/latch_enable_in scanchain_284/module_data_in[0]
+ scanchain_284/module_data_in[1] scanchain_284/module_data_in[2] scanchain_284/module_data_in[3]
+ scanchain_284/module_data_in[4] scanchain_284/module_data_in[5] scanchain_284/module_data_in[6]
+ scanchain_284/module_data_in[7] scanchain_284/module_data_out[0] scanchain_284/module_data_out[1]
+ scanchain_284/module_data_out[2] scanchain_284/module_data_out[3] scanchain_284/module_data_out[4]
+ scanchain_284/module_data_out[5] scanchain_284/module_data_out[6] scanchain_284/module_data_out[7]
+ scanchain_284/scan_select_in scanchain_285/scan_select_in vccd1 vssd1 scanchain
Xscanchain_295 scanchain_295/clk_in scanchain_296/clk_in scanchain_295/data_in scanchain_296/data_in
+ scanchain_295/latch_enable_in scanchain_296/latch_enable_in scanchain_295/module_data_in[0]
+ scanchain_295/module_data_in[1] scanchain_295/module_data_in[2] scanchain_295/module_data_in[3]
+ scanchain_295/module_data_in[4] scanchain_295/module_data_in[5] scanchain_295/module_data_in[6]
+ scanchain_295/module_data_in[7] scanchain_295/module_data_out[0] scanchain_295/module_data_out[1]
+ scanchain_295/module_data_out[2] scanchain_295/module_data_out[3] scanchain_295/module_data_out[4]
+ scanchain_295/module_data_out[5] scanchain_295/module_data_out[6] scanchain_295/module_data_out[7]
+ scanchain_295/scan_select_in scanchain_296/scan_select_in vccd1 vssd1 scanchain
Xscanchain_273 scanchain_273/clk_in scanchain_274/clk_in scanchain_273/data_in scanchain_274/data_in
+ scanchain_273/latch_enable_in scanchain_274/latch_enable_in scanchain_273/module_data_in[0]
+ scanchain_273/module_data_in[1] scanchain_273/module_data_in[2] scanchain_273/module_data_in[3]
+ scanchain_273/module_data_in[4] scanchain_273/module_data_in[5] scanchain_273/module_data_in[6]
+ scanchain_273/module_data_in[7] scanchain_273/module_data_out[0] scanchain_273/module_data_out[1]
+ scanchain_273/module_data_out[2] scanchain_273/module_data_out[3] scanchain_273/module_data_out[4]
+ scanchain_273/module_data_out[5] scanchain_273/module_data_out[6] scanchain_273/module_data_out[7]
+ scanchain_273/scan_select_in scanchain_274/scan_select_in vccd1 vssd1 scanchain
Xscanchain_251 scanchain_251/clk_in scanchain_252/clk_in scanchain_251/data_in scanchain_252/data_in
+ scanchain_251/latch_enable_in scanchain_252/latch_enable_in scanchain_251/module_data_in[0]
+ scanchain_251/module_data_in[1] scanchain_251/module_data_in[2] scanchain_251/module_data_in[3]
+ scanchain_251/module_data_in[4] scanchain_251/module_data_in[5] scanchain_251/module_data_in[6]
+ scanchain_251/module_data_in[7] scanchain_251/module_data_out[0] scanchain_251/module_data_out[1]
+ scanchain_251/module_data_out[2] scanchain_251/module_data_out[3] scanchain_251/module_data_out[4]
+ scanchain_251/module_data_out[5] scanchain_251/module_data_out[6] scanchain_251/module_data_out[7]
+ scanchain_251/scan_select_in scanchain_252/scan_select_in vccd1 vssd1 scanchain
Xscanchain_262 scanchain_262/clk_in scanchain_263/clk_in scanchain_262/data_in scanchain_263/data_in
+ scanchain_262/latch_enable_in scanchain_263/latch_enable_in scanchain_262/module_data_in[0]
+ scanchain_262/module_data_in[1] scanchain_262/module_data_in[2] scanchain_262/module_data_in[3]
+ scanchain_262/module_data_in[4] scanchain_262/module_data_in[5] scanchain_262/module_data_in[6]
+ scanchain_262/module_data_in[7] scanchain_262/module_data_out[0] scanchain_262/module_data_out[1]
+ scanchain_262/module_data_out[2] scanchain_262/module_data_out[3] scanchain_262/module_data_out[4]
+ scanchain_262/module_data_out[5] scanchain_262/module_data_out[6] scanchain_262/module_data_out[7]
+ scanchain_262/scan_select_in scanchain_263/scan_select_in vccd1 vssd1 scanchain
Xscanchain_240 scanchain_240/clk_in scanchain_241/clk_in scanchain_240/data_in scanchain_241/data_in
+ scanchain_240/latch_enable_in scanchain_241/latch_enable_in scanchain_240/module_data_in[0]
+ scanchain_240/module_data_in[1] scanchain_240/module_data_in[2] scanchain_240/module_data_in[3]
+ scanchain_240/module_data_in[4] scanchain_240/module_data_in[5] scanchain_240/module_data_in[6]
+ scanchain_240/module_data_in[7] scanchain_240/module_data_out[0] scanchain_240/module_data_out[1]
+ scanchain_240/module_data_out[2] scanchain_240/module_data_out[3] scanchain_240/module_data_out[4]
+ scanchain_240/module_data_out[5] scanchain_240/module_data_out[6] scanchain_240/module_data_out[7]
+ scanchain_240/scan_select_in scanchain_241/scan_select_in vccd1 vssd1 scanchain
Xscanchain_5 scanchain_5/clk_in scanchain_6/clk_in scanchain_5/data_in scanchain_6/data_in
+ scanchain_5/latch_enable_in scanchain_6/latch_enable_in migcorre_pwm_5/io_in[0]
+ migcorre_pwm_5/io_in[1] migcorre_pwm_5/io_in[2] migcorre_pwm_5/io_in[3] migcorre_pwm_5/io_in[4]
+ migcorre_pwm_5/io_in[5] migcorre_pwm_5/io_in[6] migcorre_pwm_5/io_in[7] migcorre_pwm_5/io_out[0]
+ migcorre_pwm_5/io_out[1] migcorre_pwm_5/io_out[2] migcorre_pwm_5/io_out[3] migcorre_pwm_5/io_out[4]
+ migcorre_pwm_5/io_out[5] migcorre_pwm_5/io_out[6] migcorre_pwm_5/io_out[7] scanchain_5/scan_select_in
+ scanchain_6/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_319 scanchain_319/module_data_in[0] scanchain_319/module_data_in[1]
+ scanchain_319/module_data_in[2] scanchain_319/module_data_in[3] scanchain_319/module_data_in[4]
+ scanchain_319/module_data_in[5] scanchain_319/module_data_in[6] scanchain_319/module_data_in[7]
+ scanchain_319/module_data_out[0] scanchain_319/module_data_out[1] scanchain_319/module_data_out[2]
+ scanchain_319/module_data_out[3] scanchain_319/module_data_out[4] scanchain_319/module_data_out[5]
+ scanchain_319/module_data_out[6] scanchain_319/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_308 scanchain_308/module_data_in[0] scanchain_308/module_data_in[1]
+ scanchain_308/module_data_in[2] scanchain_308/module_data_in[3] scanchain_308/module_data_in[4]
+ scanchain_308/module_data_in[5] scanchain_308/module_data_in[6] scanchain_308/module_data_in[7]
+ scanchain_308/module_data_out[0] scanchain_308/module_data_out[1] scanchain_308/module_data_out[2]
+ scanchain_308/module_data_out[3] scanchain_308/module_data_out[4] scanchain_308/module_data_out[5]
+ scanchain_308/module_data_out[6] scanchain_308/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_105 scanchain_105/module_data_in[0] scanchain_105/module_data_in[1]
+ scanchain_105/module_data_in[2] scanchain_105/module_data_in[3] scanchain_105/module_data_in[4]
+ scanchain_105/module_data_in[5] scanchain_105/module_data_in[6] scanchain_105/module_data_in[7]
+ scanchain_105/module_data_out[0] scanchain_105/module_data_out[1] scanchain_105/module_data_out[2]
+ scanchain_105/module_data_out[3] scanchain_105/module_data_out[4] scanchain_105/module_data_out[5]
+ scanchain_105/module_data_out[6] scanchain_105/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_116 scanchain_116/module_data_in[0] scanchain_116/module_data_in[1]
+ scanchain_116/module_data_in[2] scanchain_116/module_data_in[3] scanchain_116/module_data_in[4]
+ scanchain_116/module_data_in[5] scanchain_116/module_data_in[6] scanchain_116/module_data_in[7]
+ scanchain_116/module_data_out[0] scanchain_116/module_data_out[1] scanchain_116/module_data_out[2]
+ scanchain_116/module_data_out[3] scanchain_116/module_data_out[4] scanchain_116/module_data_out[5]
+ scanchain_116/module_data_out[6] scanchain_116/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_127 scanchain_127/module_data_in[0] scanchain_127/module_data_in[1]
+ scanchain_127/module_data_in[2] scanchain_127/module_data_in[3] scanchain_127/module_data_in[4]
+ scanchain_127/module_data_in[5] scanchain_127/module_data_in[6] scanchain_127/module_data_in[7]
+ scanchain_127/module_data_out[0] scanchain_127/module_data_out[1] scanchain_127/module_data_out[2]
+ scanchain_127/module_data_out[3] scanchain_127/module_data_out[4] scanchain_127/module_data_out[5]
+ scanchain_127/module_data_out[6] scanchain_127/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_149 scanchain_149/module_data_in[0] scanchain_149/module_data_in[1]
+ scanchain_149/module_data_in[2] scanchain_149/module_data_in[3] scanchain_149/module_data_in[4]
+ scanchain_149/module_data_in[5] scanchain_149/module_data_in[6] scanchain_149/module_data_in[7]
+ scanchain_149/module_data_out[0] scanchain_149/module_data_out[1] scanchain_149/module_data_out[2]
+ scanchain_149/module_data_out[3] scanchain_149/module_data_out[4] scanchain_149/module_data_out[5]
+ scanchain_149/module_data_out[6] scanchain_149/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_138 scanchain_138/module_data_in[0] scanchain_138/module_data_in[1]
+ scanchain_138/module_data_in[2] scanchain_138/module_data_in[3] scanchain_138/module_data_in[4]
+ scanchain_138/module_data_in[5] scanchain_138/module_data_in[6] scanchain_138/module_data_in[7]
+ scanchain_138/module_data_out[0] scanchain_138/module_data_out[1] scanchain_138/module_data_out[2]
+ scanchain_138/module_data_out[3] scanchain_138/module_data_out[4] scanchain_138/module_data_out[5]
+ scanchain_138/module_data_out[6] scanchain_138/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_400 scanchain_400/clk_in scanchain_401/clk_in scanchain_400/data_in scanchain_401/data_in
+ scanchain_400/latch_enable_in scanchain_401/latch_enable_in scanchain_400/module_data_in[0]
+ scanchain_400/module_data_in[1] scanchain_400/module_data_in[2] scanchain_400/module_data_in[3]
+ scanchain_400/module_data_in[4] scanchain_400/module_data_in[5] scanchain_400/module_data_in[6]
+ scanchain_400/module_data_in[7] scanchain_400/module_data_out[0] scanchain_400/module_data_out[1]
+ scanchain_400/module_data_out[2] scanchain_400/module_data_out[3] scanchain_400/module_data_out[4]
+ scanchain_400/module_data_out[5] scanchain_400/module_data_out[6] scanchain_400/module_data_out[7]
+ scanchain_400/scan_select_in scanchain_401/scan_select_in vccd1 vssd1 scanchain
Xscanchain_466 scanchain_466/clk_in scanchain_467/clk_in scanchain_466/data_in scanchain_467/data_in
+ scanchain_466/latch_enable_in scanchain_467/latch_enable_in scanchain_466/module_data_in[0]
+ scanchain_466/module_data_in[1] scanchain_466/module_data_in[2] scanchain_466/module_data_in[3]
+ scanchain_466/module_data_in[4] scanchain_466/module_data_in[5] scanchain_466/module_data_in[6]
+ scanchain_466/module_data_in[7] scanchain_466/module_data_out[0] scanchain_466/module_data_out[1]
+ scanchain_466/module_data_out[2] scanchain_466/module_data_out[3] scanchain_466/module_data_out[4]
+ scanchain_466/module_data_out[5] scanchain_466/module_data_out[6] scanchain_466/module_data_out[7]
+ scanchain_466/scan_select_in scanchain_467/scan_select_in vccd1 vssd1 scanchain
Xscanchain_455 scanchain_455/clk_in scanchain_456/clk_in scanchain_455/data_in scanchain_456/data_in
+ scanchain_455/latch_enable_in scanchain_456/latch_enable_in scanchain_455/module_data_in[0]
+ scanchain_455/module_data_in[1] scanchain_455/module_data_in[2] scanchain_455/module_data_in[3]
+ scanchain_455/module_data_in[4] scanchain_455/module_data_in[5] scanchain_455/module_data_in[6]
+ scanchain_455/module_data_in[7] scanchain_455/module_data_out[0] scanchain_455/module_data_out[1]
+ scanchain_455/module_data_out[2] scanchain_455/module_data_out[3] scanchain_455/module_data_out[4]
+ scanchain_455/module_data_out[5] scanchain_455/module_data_out[6] scanchain_455/module_data_out[7]
+ scanchain_455/scan_select_in scanchain_456/scan_select_in vccd1 vssd1 scanchain
Xscanchain_444 scanchain_444/clk_in scanchain_445/clk_in scanchain_444/data_in scanchain_445/data_in
+ scanchain_444/latch_enable_in scanchain_445/latch_enable_in scanchain_444/module_data_in[0]
+ scanchain_444/module_data_in[1] scanchain_444/module_data_in[2] scanchain_444/module_data_in[3]
+ scanchain_444/module_data_in[4] scanchain_444/module_data_in[5] scanchain_444/module_data_in[6]
+ scanchain_444/module_data_in[7] scanchain_444/module_data_out[0] scanchain_444/module_data_out[1]
+ scanchain_444/module_data_out[2] scanchain_444/module_data_out[3] scanchain_444/module_data_out[4]
+ scanchain_444/module_data_out[5] scanchain_444/module_data_out[6] scanchain_444/module_data_out[7]
+ scanchain_444/scan_select_in scanchain_445/scan_select_in vccd1 vssd1 scanchain
Xscanchain_433 scanchain_433/clk_in scanchain_434/clk_in scanchain_433/data_in scanchain_434/data_in
+ scanchain_433/latch_enable_in scanchain_434/latch_enable_in scanchain_433/module_data_in[0]
+ scanchain_433/module_data_in[1] scanchain_433/module_data_in[2] scanchain_433/module_data_in[3]
+ scanchain_433/module_data_in[4] scanchain_433/module_data_in[5] scanchain_433/module_data_in[6]
+ scanchain_433/module_data_in[7] scanchain_433/module_data_out[0] scanchain_433/module_data_out[1]
+ scanchain_433/module_data_out[2] scanchain_433/module_data_out[3] scanchain_433/module_data_out[4]
+ scanchain_433/module_data_out[5] scanchain_433/module_data_out[6] scanchain_433/module_data_out[7]
+ scanchain_433/scan_select_in scanchain_434/scan_select_in vccd1 vssd1 scanchain
Xscanchain_422 scanchain_422/clk_in scanchain_423/clk_in scanchain_422/data_in scanchain_423/data_in
+ scanchain_422/latch_enable_in scanchain_423/latch_enable_in scanchain_422/module_data_in[0]
+ scanchain_422/module_data_in[1] scanchain_422/module_data_in[2] scanchain_422/module_data_in[3]
+ scanchain_422/module_data_in[4] scanchain_422/module_data_in[5] scanchain_422/module_data_in[6]
+ scanchain_422/module_data_in[7] scanchain_422/module_data_out[0] scanchain_422/module_data_out[1]
+ scanchain_422/module_data_out[2] scanchain_422/module_data_out[3] scanchain_422/module_data_out[4]
+ scanchain_422/module_data_out[5] scanchain_422/module_data_out[6] scanchain_422/module_data_out[7]
+ scanchain_422/scan_select_in scanchain_423/scan_select_in vccd1 vssd1 scanchain
Xscanchain_411 scanchain_411/clk_in scanchain_412/clk_in scanchain_411/data_in scanchain_412/data_in
+ scanchain_411/latch_enable_in scanchain_412/latch_enable_in scanchain_411/module_data_in[0]
+ scanchain_411/module_data_in[1] scanchain_411/module_data_in[2] scanchain_411/module_data_in[3]
+ scanchain_411/module_data_in[4] scanchain_411/module_data_in[5] scanchain_411/module_data_in[6]
+ scanchain_411/module_data_in[7] scanchain_411/module_data_out[0] scanchain_411/module_data_out[1]
+ scanchain_411/module_data_out[2] scanchain_411/module_data_out[3] scanchain_411/module_data_out[4]
+ scanchain_411/module_data_out[5] scanchain_411/module_data_out[6] scanchain_411/module_data_out[7]
+ scanchain_411/scan_select_in scanchain_412/scan_select_in vccd1 vssd1 scanchain
Xscanchain_285 scanchain_285/clk_in scanchain_286/clk_in scanchain_285/data_in scanchain_286/data_in
+ scanchain_285/latch_enable_in scanchain_286/latch_enable_in scanchain_285/module_data_in[0]
+ scanchain_285/module_data_in[1] scanchain_285/module_data_in[2] scanchain_285/module_data_in[3]
+ scanchain_285/module_data_in[4] scanchain_285/module_data_in[5] scanchain_285/module_data_in[6]
+ scanchain_285/module_data_in[7] scanchain_285/module_data_out[0] scanchain_285/module_data_out[1]
+ scanchain_285/module_data_out[2] scanchain_285/module_data_out[3] scanchain_285/module_data_out[4]
+ scanchain_285/module_data_out[5] scanchain_285/module_data_out[6] scanchain_285/module_data_out[7]
+ scanchain_285/scan_select_in scanchain_286/scan_select_in vccd1 vssd1 scanchain
Xscanchain_296 scanchain_296/clk_in scanchain_297/clk_in scanchain_296/data_in scanchain_297/data_in
+ scanchain_296/latch_enable_in scanchain_297/latch_enable_in scanchain_296/module_data_in[0]
+ scanchain_296/module_data_in[1] scanchain_296/module_data_in[2] scanchain_296/module_data_in[3]
+ scanchain_296/module_data_in[4] scanchain_296/module_data_in[5] scanchain_296/module_data_in[6]
+ scanchain_296/module_data_in[7] scanchain_296/module_data_out[0] scanchain_296/module_data_out[1]
+ scanchain_296/module_data_out[2] scanchain_296/module_data_out[3] scanchain_296/module_data_out[4]
+ scanchain_296/module_data_out[5] scanchain_296/module_data_out[6] scanchain_296/module_data_out[7]
+ scanchain_296/scan_select_in scanchain_297/scan_select_in vccd1 vssd1 scanchain
Xscanchain_274 scanchain_274/clk_in scanchain_275/clk_in scanchain_274/data_in scanchain_275/data_in
+ scanchain_274/latch_enable_in scanchain_275/latch_enable_in scanchain_274/module_data_in[0]
+ scanchain_274/module_data_in[1] scanchain_274/module_data_in[2] scanchain_274/module_data_in[3]
+ scanchain_274/module_data_in[4] scanchain_274/module_data_in[5] scanchain_274/module_data_in[6]
+ scanchain_274/module_data_in[7] scanchain_274/module_data_out[0] scanchain_274/module_data_out[1]
+ scanchain_274/module_data_out[2] scanchain_274/module_data_out[3] scanchain_274/module_data_out[4]
+ scanchain_274/module_data_out[5] scanchain_274/module_data_out[6] scanchain_274/module_data_out[7]
+ scanchain_274/scan_select_in scanchain_275/scan_select_in vccd1 vssd1 scanchain
Xscanchain_252 scanchain_252/clk_in scanchain_253/clk_in scanchain_252/data_in scanchain_253/data_in
+ scanchain_252/latch_enable_in scanchain_253/latch_enable_in scanchain_252/module_data_in[0]
+ scanchain_252/module_data_in[1] scanchain_252/module_data_in[2] scanchain_252/module_data_in[3]
+ scanchain_252/module_data_in[4] scanchain_252/module_data_in[5] scanchain_252/module_data_in[6]
+ scanchain_252/module_data_in[7] scanchain_252/module_data_out[0] scanchain_252/module_data_out[1]
+ scanchain_252/module_data_out[2] scanchain_252/module_data_out[3] scanchain_252/module_data_out[4]
+ scanchain_252/module_data_out[5] scanchain_252/module_data_out[6] scanchain_252/module_data_out[7]
+ scanchain_252/scan_select_in scanchain_253/scan_select_in vccd1 vssd1 scanchain
Xscanchain_263 scanchain_263/clk_in scanchain_264/clk_in scanchain_263/data_in scanchain_264/data_in
+ scanchain_263/latch_enable_in scanchain_264/latch_enable_in scanchain_263/module_data_in[0]
+ scanchain_263/module_data_in[1] scanchain_263/module_data_in[2] scanchain_263/module_data_in[3]
+ scanchain_263/module_data_in[4] scanchain_263/module_data_in[5] scanchain_263/module_data_in[6]
+ scanchain_263/module_data_in[7] scanchain_263/module_data_out[0] scanchain_263/module_data_out[1]
+ scanchain_263/module_data_out[2] scanchain_263/module_data_out[3] scanchain_263/module_data_out[4]
+ scanchain_263/module_data_out[5] scanchain_263/module_data_out[6] scanchain_263/module_data_out[7]
+ scanchain_263/scan_select_in scanchain_264/scan_select_in vccd1 vssd1 scanchain
Xscanchain_241 scanchain_241/clk_in scanchain_242/clk_in scanchain_241/data_in scanchain_242/data_in
+ scanchain_241/latch_enable_in scanchain_242/latch_enable_in scanchain_241/module_data_in[0]
+ scanchain_241/module_data_in[1] scanchain_241/module_data_in[2] scanchain_241/module_data_in[3]
+ scanchain_241/module_data_in[4] scanchain_241/module_data_in[5] scanchain_241/module_data_in[6]
+ scanchain_241/module_data_in[7] scanchain_241/module_data_out[0] scanchain_241/module_data_out[1]
+ scanchain_241/module_data_out[2] scanchain_241/module_data_out[3] scanchain_241/module_data_out[4]
+ scanchain_241/module_data_out[5] scanchain_241/module_data_out[6] scanchain_241/module_data_out[7]
+ scanchain_241/scan_select_in scanchain_242/scan_select_in vccd1 vssd1 scanchain
Xscanchain_230 scanchain_230/clk_in scanchain_231/clk_in scanchain_230/data_in scanchain_231/data_in
+ scanchain_230/latch_enable_in scanchain_231/latch_enable_in scanchain_230/module_data_in[0]
+ scanchain_230/module_data_in[1] scanchain_230/module_data_in[2] scanchain_230/module_data_in[3]
+ scanchain_230/module_data_in[4] scanchain_230/module_data_in[5] scanchain_230/module_data_in[6]
+ scanchain_230/module_data_in[7] scanchain_230/module_data_out[0] scanchain_230/module_data_out[1]
+ scanchain_230/module_data_out[2] scanchain_230/module_data_out[3] scanchain_230/module_data_out[4]
+ scanchain_230/module_data_out[5] scanchain_230/module_data_out[6] scanchain_230/module_data_out[7]
+ scanchain_230/scan_select_in scanchain_231/scan_select_in vccd1 vssd1 scanchain
Xscanchain_6 scanchain_6/clk_in scanchain_7/clk_in scanchain_6/data_in scanchain_7/data_in
+ scanchain_6/latch_enable_in scanchain_7/latch_enable_in s4ga_6/io_in[0] s4ga_6/io_in[1]
+ s4ga_6/io_in[2] s4ga_6/io_in[3] s4ga_6/io_in[4] s4ga_6/io_in[5] s4ga_6/io_in[6]
+ s4ga_6/io_in[7] s4ga_6/io_out[0] s4ga_6/io_out[1] s4ga_6/io_out[2] s4ga_6/io_out[3]
+ s4ga_6/io_out[4] s4ga_6/io_out[5] s4ga_6/io_out[6] s4ga_6/io_out[7] scanchain_6/scan_select_in
+ scanchain_7/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_309 scanchain_309/module_data_in[0] scanchain_309/module_data_in[1]
+ scanchain_309/module_data_in[2] scanchain_309/module_data_in[3] scanchain_309/module_data_in[4]
+ scanchain_309/module_data_in[5] scanchain_309/module_data_in[6] scanchain_309/module_data_in[7]
+ scanchain_309/module_data_out[0] scanchain_309/module_data_out[1] scanchain_309/module_data_out[2]
+ scanchain_309/module_data_out[3] scanchain_309/module_data_out[4] scanchain_309/module_data_out[5]
+ scanchain_309/module_data_out[6] scanchain_309/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_90 scanchain_90/clk_in scanchain_91/clk_in scanchain_90/data_in scanchain_91/data_in
+ scanchain_90/latch_enable_in scanchain_91/latch_enable_in scanchain_90/module_data_in[0]
+ scanchain_90/module_data_in[1] scanchain_90/module_data_in[2] scanchain_90/module_data_in[3]
+ scanchain_90/module_data_in[4] scanchain_90/module_data_in[5] scanchain_90/module_data_in[6]
+ scanchain_90/module_data_in[7] scanchain_90/module_data_out[0] scanchain_90/module_data_out[1]
+ scanchain_90/module_data_out[2] scanchain_90/module_data_out[3] scanchain_90/module_data_out[4]
+ scanchain_90/module_data_out[5] scanchain_90/module_data_out[6] scanchain_90/module_data_out[7]
+ scanchain_90/scan_select_in scanchain_91/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_106 scanchain_106/module_data_in[0] scanchain_106/module_data_in[1]
+ scanchain_106/module_data_in[2] scanchain_106/module_data_in[3] scanchain_106/module_data_in[4]
+ scanchain_106/module_data_in[5] scanchain_106/module_data_in[6] scanchain_106/module_data_in[7]
+ scanchain_106/module_data_out[0] scanchain_106/module_data_out[1] scanchain_106/module_data_out[2]
+ scanchain_106/module_data_out[3] scanchain_106/module_data_out[4] scanchain_106/module_data_out[5]
+ scanchain_106/module_data_out[6] scanchain_106/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_117 scanchain_117/module_data_in[0] scanchain_117/module_data_in[1]
+ scanchain_117/module_data_in[2] scanchain_117/module_data_in[3] scanchain_117/module_data_in[4]
+ scanchain_117/module_data_in[5] scanchain_117/module_data_in[6] scanchain_117/module_data_in[7]
+ scanchain_117/module_data_out[0] scanchain_117/module_data_out[1] scanchain_117/module_data_out[2]
+ scanchain_117/module_data_out[3] scanchain_117/module_data_out[4] scanchain_117/module_data_out[5]
+ scanchain_117/module_data_out[6] scanchain_117/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_128 scanchain_128/module_data_in[0] scanchain_128/module_data_in[1]
+ scanchain_128/module_data_in[2] scanchain_128/module_data_in[3] scanchain_128/module_data_in[4]
+ scanchain_128/module_data_in[5] scanchain_128/module_data_in[6] scanchain_128/module_data_in[7]
+ scanchain_128/module_data_out[0] scanchain_128/module_data_out[1] scanchain_128/module_data_out[2]
+ scanchain_128/module_data_out[3] scanchain_128/module_data_out[4] scanchain_128/module_data_out[5]
+ scanchain_128/module_data_out[6] scanchain_128/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_139 scanchain_139/module_data_in[0] scanchain_139/module_data_in[1]
+ scanchain_139/module_data_in[2] scanchain_139/module_data_in[3] scanchain_139/module_data_in[4]
+ scanchain_139/module_data_in[5] scanchain_139/module_data_in[6] scanchain_139/module_data_in[7]
+ scanchain_139/module_data_out[0] scanchain_139/module_data_out[1] scanchain_139/module_data_out[2]
+ scanchain_139/module_data_out[3] scanchain_139/module_data_out[4] scanchain_139/module_data_out[5]
+ scanchain_139/module_data_out[6] scanchain_139/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xtt2_tholin_namebadge_55 scanchain_55/module_data_in[0] scanchain_55/module_data_in[1]
+ scanchain_55/module_data_in[2] scanchain_55/module_data_in[3] scanchain_55/module_data_in[4]
+ scanchain_55/module_data_in[5] scanchain_55/module_data_in[6] scanchain_55/module_data_in[7]
+ scanchain_55/module_data_out[0] scanchain_55/module_data_out[1] scanchain_55/module_data_out[2]
+ scanchain_55/module_data_out[3] scanchain_55/module_data_out[4] scanchain_55/module_data_out[5]
+ scanchain_55/module_data_out[6] scanchain_55/module_data_out[7] vccd1 vssd1 tt2_tholin_namebadge
Xuser_module_339501025136214612_470 scanchain_470/module_data_in[0] scanchain_470/module_data_in[1]
+ scanchain_470/module_data_in[2] scanchain_470/module_data_in[3] scanchain_470/module_data_in[4]
+ scanchain_470/module_data_in[5] scanchain_470/module_data_in[6] scanchain_470/module_data_in[7]
+ scanchain_470/module_data_out[0] scanchain_470/module_data_out[1] scanchain_470/module_data_out[2]
+ scanchain_470/module_data_out[3] scanchain_470/module_data_out[4] scanchain_470/module_data_out[5]
+ scanchain_470/module_data_out[6] scanchain_470/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_467 scanchain_467/clk_in scanchain_468/clk_in scanchain_467/data_in scanchain_468/data_in
+ scanchain_467/latch_enable_in scanchain_468/latch_enable_in scanchain_467/module_data_in[0]
+ scanchain_467/module_data_in[1] scanchain_467/module_data_in[2] scanchain_467/module_data_in[3]
+ scanchain_467/module_data_in[4] scanchain_467/module_data_in[5] scanchain_467/module_data_in[6]
+ scanchain_467/module_data_in[7] scanchain_467/module_data_out[0] scanchain_467/module_data_out[1]
+ scanchain_467/module_data_out[2] scanchain_467/module_data_out[3] scanchain_467/module_data_out[4]
+ scanchain_467/module_data_out[5] scanchain_467/module_data_out[6] scanchain_467/module_data_out[7]
+ scanchain_467/scan_select_in scanchain_468/scan_select_in vccd1 vssd1 scanchain
Xscanchain_456 scanchain_456/clk_in scanchain_457/clk_in scanchain_456/data_in scanchain_457/data_in
+ scanchain_456/latch_enable_in scanchain_457/latch_enable_in scanchain_456/module_data_in[0]
+ scanchain_456/module_data_in[1] scanchain_456/module_data_in[2] scanchain_456/module_data_in[3]
+ scanchain_456/module_data_in[4] scanchain_456/module_data_in[5] scanchain_456/module_data_in[6]
+ scanchain_456/module_data_in[7] scanchain_456/module_data_out[0] scanchain_456/module_data_out[1]
+ scanchain_456/module_data_out[2] scanchain_456/module_data_out[3] scanchain_456/module_data_out[4]
+ scanchain_456/module_data_out[5] scanchain_456/module_data_out[6] scanchain_456/module_data_out[7]
+ scanchain_456/scan_select_in scanchain_457/scan_select_in vccd1 vssd1 scanchain
Xscanchain_445 scanchain_445/clk_in scanchain_446/clk_in scanchain_445/data_in scanchain_446/data_in
+ scanchain_445/latch_enable_in scanchain_446/latch_enable_in scanchain_445/module_data_in[0]
+ scanchain_445/module_data_in[1] scanchain_445/module_data_in[2] scanchain_445/module_data_in[3]
+ scanchain_445/module_data_in[4] scanchain_445/module_data_in[5] scanchain_445/module_data_in[6]
+ scanchain_445/module_data_in[7] scanchain_445/module_data_out[0] scanchain_445/module_data_out[1]
+ scanchain_445/module_data_out[2] scanchain_445/module_data_out[3] scanchain_445/module_data_out[4]
+ scanchain_445/module_data_out[5] scanchain_445/module_data_out[6] scanchain_445/module_data_out[7]
+ scanchain_445/scan_select_in scanchain_446/scan_select_in vccd1 vssd1 scanchain
Xscanchain_434 scanchain_434/clk_in scanchain_435/clk_in scanchain_434/data_in scanchain_435/data_in
+ scanchain_434/latch_enable_in scanchain_435/latch_enable_in scanchain_434/module_data_in[0]
+ scanchain_434/module_data_in[1] scanchain_434/module_data_in[2] scanchain_434/module_data_in[3]
+ scanchain_434/module_data_in[4] scanchain_434/module_data_in[5] scanchain_434/module_data_in[6]
+ scanchain_434/module_data_in[7] scanchain_434/module_data_out[0] scanchain_434/module_data_out[1]
+ scanchain_434/module_data_out[2] scanchain_434/module_data_out[3] scanchain_434/module_data_out[4]
+ scanchain_434/module_data_out[5] scanchain_434/module_data_out[6] scanchain_434/module_data_out[7]
+ scanchain_434/scan_select_in scanchain_435/scan_select_in vccd1 vssd1 scanchain
Xscanchain_423 scanchain_423/clk_in scanchain_424/clk_in scanchain_423/data_in scanchain_424/data_in
+ scanchain_423/latch_enable_in scanchain_424/latch_enable_in scanchain_423/module_data_in[0]
+ scanchain_423/module_data_in[1] scanchain_423/module_data_in[2] scanchain_423/module_data_in[3]
+ scanchain_423/module_data_in[4] scanchain_423/module_data_in[5] scanchain_423/module_data_in[6]
+ scanchain_423/module_data_in[7] scanchain_423/module_data_out[0] scanchain_423/module_data_out[1]
+ scanchain_423/module_data_out[2] scanchain_423/module_data_out[3] scanchain_423/module_data_out[4]
+ scanchain_423/module_data_out[5] scanchain_423/module_data_out[6] scanchain_423/module_data_out[7]
+ scanchain_423/scan_select_in scanchain_424/scan_select_in vccd1 vssd1 scanchain
Xscanchain_401 scanchain_401/clk_in scanchain_402/clk_in scanchain_401/data_in scanchain_402/data_in
+ scanchain_401/latch_enable_in scanchain_402/latch_enable_in scanchain_401/module_data_in[0]
+ scanchain_401/module_data_in[1] scanchain_401/module_data_in[2] scanchain_401/module_data_in[3]
+ scanchain_401/module_data_in[4] scanchain_401/module_data_in[5] scanchain_401/module_data_in[6]
+ scanchain_401/module_data_in[7] scanchain_401/module_data_out[0] scanchain_401/module_data_out[1]
+ scanchain_401/module_data_out[2] scanchain_401/module_data_out[3] scanchain_401/module_data_out[4]
+ scanchain_401/module_data_out[5] scanchain_401/module_data_out[6] scanchain_401/module_data_out[7]
+ scanchain_401/scan_select_in scanchain_402/scan_select_in vccd1 vssd1 scanchain
Xscanchain_412 scanchain_412/clk_in scanchain_413/clk_in scanchain_412/data_in scanchain_413/data_in
+ scanchain_412/latch_enable_in scanchain_413/latch_enable_in scanchain_412/module_data_in[0]
+ scanchain_412/module_data_in[1] scanchain_412/module_data_in[2] scanchain_412/module_data_in[3]
+ scanchain_412/module_data_in[4] scanchain_412/module_data_in[5] scanchain_412/module_data_in[6]
+ scanchain_412/module_data_in[7] scanchain_412/module_data_out[0] scanchain_412/module_data_out[1]
+ scanchain_412/module_data_out[2] scanchain_412/module_data_out[3] scanchain_412/module_data_out[4]
+ scanchain_412/module_data_out[5] scanchain_412/module_data_out[6] scanchain_412/module_data_out[7]
+ scanchain_412/scan_select_in scanchain_413/scan_select_in vccd1 vssd1 scanchain
Xscanchain_275 scanchain_275/clk_in scanchain_276/clk_in scanchain_275/data_in scanchain_276/data_in
+ scanchain_275/latch_enable_in scanchain_276/latch_enable_in scanchain_275/module_data_in[0]
+ scanchain_275/module_data_in[1] scanchain_275/module_data_in[2] scanchain_275/module_data_in[3]
+ scanchain_275/module_data_in[4] scanchain_275/module_data_in[5] scanchain_275/module_data_in[6]
+ scanchain_275/module_data_in[7] scanchain_275/module_data_out[0] scanchain_275/module_data_out[1]
+ scanchain_275/module_data_out[2] scanchain_275/module_data_out[3] scanchain_275/module_data_out[4]
+ scanchain_275/module_data_out[5] scanchain_275/module_data_out[6] scanchain_275/module_data_out[7]
+ scanchain_275/scan_select_in scanchain_276/scan_select_in vccd1 vssd1 scanchain
Xscanchain_264 scanchain_264/clk_in scanchain_265/clk_in scanchain_264/data_in scanchain_265/data_in
+ scanchain_264/latch_enable_in scanchain_265/latch_enable_in scanchain_264/module_data_in[0]
+ scanchain_264/module_data_in[1] scanchain_264/module_data_in[2] scanchain_264/module_data_in[3]
+ scanchain_264/module_data_in[4] scanchain_264/module_data_in[5] scanchain_264/module_data_in[6]
+ scanchain_264/module_data_in[7] scanchain_264/module_data_out[0] scanchain_264/module_data_out[1]
+ scanchain_264/module_data_out[2] scanchain_264/module_data_out[3] scanchain_264/module_data_out[4]
+ scanchain_264/module_data_out[5] scanchain_264/module_data_out[6] scanchain_264/module_data_out[7]
+ scanchain_264/scan_select_in scanchain_265/scan_select_in vccd1 vssd1 scanchain
Xscanchain_253 scanchain_253/clk_in scanchain_254/clk_in scanchain_253/data_in scanchain_254/data_in
+ scanchain_253/latch_enable_in scanchain_254/latch_enable_in scanchain_253/module_data_in[0]
+ scanchain_253/module_data_in[1] scanchain_253/module_data_in[2] scanchain_253/module_data_in[3]
+ scanchain_253/module_data_in[4] scanchain_253/module_data_in[5] scanchain_253/module_data_in[6]
+ scanchain_253/module_data_in[7] scanchain_253/module_data_out[0] scanchain_253/module_data_out[1]
+ scanchain_253/module_data_out[2] scanchain_253/module_data_out[3] scanchain_253/module_data_out[4]
+ scanchain_253/module_data_out[5] scanchain_253/module_data_out[6] scanchain_253/module_data_out[7]
+ scanchain_253/scan_select_in scanchain_254/scan_select_in vccd1 vssd1 scanchain
Xscanchain_242 scanchain_242/clk_in scanchain_243/clk_in scanchain_242/data_in scanchain_243/data_in
+ scanchain_242/latch_enable_in scanchain_243/latch_enable_in scanchain_242/module_data_in[0]
+ scanchain_242/module_data_in[1] scanchain_242/module_data_in[2] scanchain_242/module_data_in[3]
+ scanchain_242/module_data_in[4] scanchain_242/module_data_in[5] scanchain_242/module_data_in[6]
+ scanchain_242/module_data_in[7] scanchain_242/module_data_out[0] scanchain_242/module_data_out[1]
+ scanchain_242/module_data_out[2] scanchain_242/module_data_out[3] scanchain_242/module_data_out[4]
+ scanchain_242/module_data_out[5] scanchain_242/module_data_out[6] scanchain_242/module_data_out[7]
+ scanchain_242/scan_select_in scanchain_243/scan_select_in vccd1 vssd1 scanchain
Xscanchain_231 scanchain_231/clk_in scanchain_232/clk_in scanchain_231/data_in scanchain_232/data_in
+ scanchain_231/latch_enable_in scanchain_232/latch_enable_in scanchain_231/module_data_in[0]
+ scanchain_231/module_data_in[1] scanchain_231/module_data_in[2] scanchain_231/module_data_in[3]
+ scanchain_231/module_data_in[4] scanchain_231/module_data_in[5] scanchain_231/module_data_in[6]
+ scanchain_231/module_data_in[7] scanchain_231/module_data_out[0] scanchain_231/module_data_out[1]
+ scanchain_231/module_data_out[2] scanchain_231/module_data_out[3] scanchain_231/module_data_out[4]
+ scanchain_231/module_data_out[5] scanchain_231/module_data_out[6] scanchain_231/module_data_out[7]
+ scanchain_231/scan_select_in scanchain_232/scan_select_in vccd1 vssd1 scanchain
Xscanchain_220 scanchain_220/clk_in scanchain_221/clk_in scanchain_220/data_in scanchain_221/data_in
+ scanchain_220/latch_enable_in scanchain_221/latch_enable_in scanchain_220/module_data_in[0]
+ scanchain_220/module_data_in[1] scanchain_220/module_data_in[2] scanchain_220/module_data_in[3]
+ scanchain_220/module_data_in[4] scanchain_220/module_data_in[5] scanchain_220/module_data_in[6]
+ scanchain_220/module_data_in[7] scanchain_220/module_data_out[0] scanchain_220/module_data_out[1]
+ scanchain_220/module_data_out[2] scanchain_220/module_data_out[3] scanchain_220/module_data_out[4]
+ scanchain_220/module_data_out[5] scanchain_220/module_data_out[6] scanchain_220/module_data_out[7]
+ scanchain_220/scan_select_in scanchain_221/scan_select_in vccd1 vssd1 scanchain
Xscanchain_286 scanchain_286/clk_in scanchain_287/clk_in scanchain_286/data_in scanchain_287/data_in
+ scanchain_286/latch_enable_in scanchain_287/latch_enable_in scanchain_286/module_data_in[0]
+ scanchain_286/module_data_in[1] scanchain_286/module_data_in[2] scanchain_286/module_data_in[3]
+ scanchain_286/module_data_in[4] scanchain_286/module_data_in[5] scanchain_286/module_data_in[6]
+ scanchain_286/module_data_in[7] scanchain_286/module_data_out[0] scanchain_286/module_data_out[1]
+ scanchain_286/module_data_out[2] scanchain_286/module_data_out[3] scanchain_286/module_data_out[4]
+ scanchain_286/module_data_out[5] scanchain_286/module_data_out[6] scanchain_286/module_data_out[7]
+ scanchain_286/scan_select_in scanchain_287/scan_select_in vccd1 vssd1 scanchain
Xscanchain_297 scanchain_297/clk_in scanchain_298/clk_in scanchain_297/data_in scanchain_298/data_in
+ scanchain_297/latch_enable_in scanchain_298/latch_enable_in scanchain_297/module_data_in[0]
+ scanchain_297/module_data_in[1] scanchain_297/module_data_in[2] scanchain_297/module_data_in[3]
+ scanchain_297/module_data_in[4] scanchain_297/module_data_in[5] scanchain_297/module_data_in[6]
+ scanchain_297/module_data_in[7] scanchain_297/module_data_out[0] scanchain_297/module_data_out[1]
+ scanchain_297/module_data_out[2] scanchain_297/module_data_out[3] scanchain_297/module_data_out[4]
+ scanchain_297/module_data_out[5] scanchain_297/module_data_out[6] scanchain_297/module_data_out[7]
+ scanchain_297/scan_select_in scanchain_298/scan_select_in vccd1 vssd1 scanchain
Xscanchain_7 scanchain_7/clk_in scanchain_8/clk_in scanchain_7/data_in scanchain_8/data_in
+ scanchain_7/latch_enable_in scanchain_8/latch_enable_in alu_top_7/io_in[0] alu_top_7/io_in[1]
+ alu_top_7/io_in[2] alu_top_7/io_in[3] alu_top_7/io_in[4] alu_top_7/io_in[5] alu_top_7/io_in[6]
+ alu_top_7/io_in[7] alu_top_7/io_out[0] alu_top_7/io_out[1] alu_top_7/io_out[2] alu_top_7/io_out[3]
+ alu_top_7/io_out[4] alu_top_7/io_out[5] alu_top_7/io_out[6] alu_top_7/io_out[7]
+ scanchain_7/scan_select_in scanchain_8/scan_select_in vccd1 vssd1 scanchain
Xtomkeddie_top_tto_2 tomkeddie_top_tto_2/io_in[0] tomkeddie_top_tto_2/io_in[1] tomkeddie_top_tto_2/io_in[2]
+ tomkeddie_top_tto_2/io_in[3] tomkeddie_top_tto_2/io_in[4] tomkeddie_top_tto_2/io_in[5]
+ tomkeddie_top_tto_2/io_in[6] tomkeddie_top_tto_2/io_in[7] tomkeddie_top_tto_2/io_out[0]
+ tomkeddie_top_tto_2/io_out[1] tomkeddie_top_tto_2/io_out[2] tomkeddie_top_tto_2/io_out[3]
+ tomkeddie_top_tto_2/io_out[4] tomkeddie_top_tto_2/io_out[5] tomkeddie_top_tto_2/io_out[6]
+ tomkeddie_top_tto_2/io_out[7] vccd1 vssd1 tomkeddie_top_tto
Xzoechip_31 zoechip_31/io_in[0] zoechip_31/io_in[1] zoechip_31/io_in[2] zoechip_31/io_in[3]
+ zoechip_31/io_in[4] zoechip_31/io_in[5] zoechip_31/io_in[6] zoechip_31/io_in[7]
+ zoechip_31/io_out[0] zoechip_31/io_out[1] zoechip_31/io_out[2] zoechip_31/io_out[3]
+ zoechip_31/io_out[4] zoechip_31/io_out[5] zoechip_31/io_out[6] zoechip_31/io_out[7]
+ vccd1 vssd1 zoechip
Xscanchain_80 scanchain_80/clk_in scanchain_81/clk_in scanchain_80/data_in scanchain_81/data_in
+ scanchain_80/latch_enable_in scanchain_81/latch_enable_in scanchain_80/module_data_in[0]
+ scanchain_80/module_data_in[1] scanchain_80/module_data_in[2] scanchain_80/module_data_in[3]
+ scanchain_80/module_data_in[4] scanchain_80/module_data_in[5] scanchain_80/module_data_in[6]
+ scanchain_80/module_data_in[7] scanchain_80/module_data_out[0] scanchain_80/module_data_out[1]
+ scanchain_80/module_data_out[2] scanchain_80/module_data_out[3] scanchain_80/module_data_out[4]
+ scanchain_80/module_data_out[5] scanchain_80/module_data_out[6] scanchain_80/module_data_out[7]
+ scanchain_80/scan_select_in scanchain_81/scan_select_in vccd1 vssd1 scanchain
Xscanchain_91 scanchain_91/clk_in scanchain_92/clk_in scanchain_91/data_in scanchain_92/data_in
+ scanchain_91/latch_enable_in scanchain_92/latch_enable_in scanchain_91/module_data_in[0]
+ scanchain_91/module_data_in[1] scanchain_91/module_data_in[2] scanchain_91/module_data_in[3]
+ scanchain_91/module_data_in[4] scanchain_91/module_data_in[5] scanchain_91/module_data_in[6]
+ scanchain_91/module_data_in[7] scanchain_91/module_data_out[0] scanchain_91/module_data_out[1]
+ scanchain_91/module_data_out[2] scanchain_91/module_data_out[3] scanchain_91/module_data_out[4]
+ scanchain_91/module_data_out[5] scanchain_91/module_data_out[6] scanchain_91/module_data_out[7]
+ scanchain_91/scan_select_in scanchain_92/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_107 scanchain_107/module_data_in[0] scanchain_107/module_data_in[1]
+ scanchain_107/module_data_in[2] scanchain_107/module_data_in[3] scanchain_107/module_data_in[4]
+ scanchain_107/module_data_in[5] scanchain_107/module_data_in[6] scanchain_107/module_data_in[7]
+ scanchain_107/module_data_out[0] scanchain_107/module_data_out[1] scanchain_107/module_data_out[2]
+ scanchain_107/module_data_out[3] scanchain_107/module_data_out[4] scanchain_107/module_data_out[5]
+ scanchain_107/module_data_out[6] scanchain_107/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_118 scanchain_118/module_data_in[0] scanchain_118/module_data_in[1]
+ scanchain_118/module_data_in[2] scanchain_118/module_data_in[3] scanchain_118/module_data_in[4]
+ scanchain_118/module_data_in[5] scanchain_118/module_data_in[6] scanchain_118/module_data_in[7]
+ scanchain_118/module_data_out[0] scanchain_118/module_data_out[1] scanchain_118/module_data_out[2]
+ scanchain_118/module_data_out[3] scanchain_118/module_data_out[4] scanchain_118/module_data_out[5]
+ scanchain_118/module_data_out[6] scanchain_118/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_129 scanchain_129/module_data_in[0] scanchain_129/module_data_in[1]
+ scanchain_129/module_data_in[2] scanchain_129/module_data_in[3] scanchain_129/module_data_in[4]
+ scanchain_129/module_data_in[5] scanchain_129/module_data_in[6] scanchain_129/module_data_in[7]
+ scanchain_129/module_data_out[0] scanchain_129/module_data_out[1] scanchain_129/module_data_out[2]
+ scanchain_129/module_data_out[3] scanchain_129/module_data_out[4] scanchain_129/module_data_out[5]
+ scanchain_129/module_data_out[6] scanchain_129/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xthezoq2_yafpga_38 thezoq2_yafpga_38/io_in[0] thezoq2_yafpga_38/io_in[1] thezoq2_yafpga_38/io_in[2]
+ thezoq2_yafpga_38/io_in[3] thezoq2_yafpga_38/io_in[4] thezoq2_yafpga_38/io_in[5]
+ thezoq2_yafpga_38/io_in[6] thezoq2_yafpga_38/io_in[7] thezoq2_yafpga_38/io_out[0]
+ thezoq2_yafpga_38/io_out[1] thezoq2_yafpga_38/io_out[2] thezoq2_yafpga_38/io_out[3]
+ thezoq2_yafpga_38/io_out[4] thezoq2_yafpga_38/io_out[5] thezoq2_yafpga_38/io_out[6]
+ thezoq2_yafpga_38/io_out[7] vccd1 vssd1 thezoq2_yafpga
Xuser_module_339501025136214612_471 scanchain_471/module_data_in[0] scanchain_471/module_data_in[1]
+ scanchain_471/module_data_in[2] scanchain_471/module_data_in[3] scanchain_471/module_data_in[4]
+ scanchain_471/module_data_in[5] scanchain_471/module_data_in[6] scanchain_471/module_data_in[7]
+ scanchain_471/module_data_out[0] scanchain_471/module_data_out[1] scanchain_471/module_data_out[2]
+ scanchain_471/module_data_out[3] scanchain_471/module_data_out[4] scanchain_471/module_data_out[5]
+ scanchain_471/module_data_out[6] scanchain_471/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_468 scanchain_468/clk_in scanchain_469/clk_in scanchain_468/data_in scanchain_469/data_in
+ scanchain_468/latch_enable_in scanchain_469/latch_enable_in scanchain_468/module_data_in[0]
+ scanchain_468/module_data_in[1] scanchain_468/module_data_in[2] scanchain_468/module_data_in[3]
+ scanchain_468/module_data_in[4] scanchain_468/module_data_in[5] scanchain_468/module_data_in[6]
+ scanchain_468/module_data_in[7] scanchain_468/module_data_out[0] scanchain_468/module_data_out[1]
+ scanchain_468/module_data_out[2] scanchain_468/module_data_out[3] scanchain_468/module_data_out[4]
+ scanchain_468/module_data_out[5] scanchain_468/module_data_out[6] scanchain_468/module_data_out[7]
+ scanchain_468/scan_select_in scanchain_469/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_460 scanchain_460/module_data_in[0] scanchain_460/module_data_in[1]
+ scanchain_460/module_data_in[2] scanchain_460/module_data_in[3] scanchain_460/module_data_in[4]
+ scanchain_460/module_data_in[5] scanchain_460/module_data_in[6] scanchain_460/module_data_in[7]
+ scanchain_460/module_data_out[0] scanchain_460/module_data_out[1] scanchain_460/module_data_out[2]
+ scanchain_460/module_data_out[3] scanchain_460/module_data_out[4] scanchain_460/module_data_out[5]
+ scanchain_460/module_data_out[6] scanchain_460/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_457 scanchain_457/clk_in scanchain_458/clk_in scanchain_457/data_in scanchain_458/data_in
+ scanchain_457/latch_enable_in scanchain_458/latch_enable_in scanchain_457/module_data_in[0]
+ scanchain_457/module_data_in[1] scanchain_457/module_data_in[2] scanchain_457/module_data_in[3]
+ scanchain_457/module_data_in[4] scanchain_457/module_data_in[5] scanchain_457/module_data_in[6]
+ scanchain_457/module_data_in[7] scanchain_457/module_data_out[0] scanchain_457/module_data_out[1]
+ scanchain_457/module_data_out[2] scanchain_457/module_data_out[3] scanchain_457/module_data_out[4]
+ scanchain_457/module_data_out[5] scanchain_457/module_data_out[6] scanchain_457/module_data_out[7]
+ scanchain_457/scan_select_in scanchain_458/scan_select_in vccd1 vssd1 scanchain
Xscanchain_435 scanchain_435/clk_in scanchain_436/clk_in scanchain_435/data_in scanchain_436/data_in
+ scanchain_435/latch_enable_in scanchain_436/latch_enable_in scanchain_435/module_data_in[0]
+ scanchain_435/module_data_in[1] scanchain_435/module_data_in[2] scanchain_435/module_data_in[3]
+ scanchain_435/module_data_in[4] scanchain_435/module_data_in[5] scanchain_435/module_data_in[6]
+ scanchain_435/module_data_in[7] scanchain_435/module_data_out[0] scanchain_435/module_data_out[1]
+ scanchain_435/module_data_out[2] scanchain_435/module_data_out[3] scanchain_435/module_data_out[4]
+ scanchain_435/module_data_out[5] scanchain_435/module_data_out[6] scanchain_435/module_data_out[7]
+ scanchain_435/scan_select_in scanchain_436/scan_select_in vccd1 vssd1 scanchain
Xscanchain_446 scanchain_446/clk_in scanchain_447/clk_in scanchain_446/data_in scanchain_447/data_in
+ scanchain_446/latch_enable_in scanchain_447/latch_enable_in scanchain_446/module_data_in[0]
+ scanchain_446/module_data_in[1] scanchain_446/module_data_in[2] scanchain_446/module_data_in[3]
+ scanchain_446/module_data_in[4] scanchain_446/module_data_in[5] scanchain_446/module_data_in[6]
+ scanchain_446/module_data_in[7] scanchain_446/module_data_out[0] scanchain_446/module_data_out[1]
+ scanchain_446/module_data_out[2] scanchain_446/module_data_out[3] scanchain_446/module_data_out[4]
+ scanchain_446/module_data_out[5] scanchain_446/module_data_out[6] scanchain_446/module_data_out[7]
+ scanchain_446/scan_select_in scanchain_447/scan_select_in vccd1 vssd1 scanchain
Xscanchain_424 scanchain_424/clk_in scanchain_425/clk_in scanchain_424/data_in scanchain_425/data_in
+ scanchain_424/latch_enable_in scanchain_425/latch_enable_in scanchain_424/module_data_in[0]
+ scanchain_424/module_data_in[1] scanchain_424/module_data_in[2] scanchain_424/module_data_in[3]
+ scanchain_424/module_data_in[4] scanchain_424/module_data_in[5] scanchain_424/module_data_in[6]
+ scanchain_424/module_data_in[7] scanchain_424/module_data_out[0] scanchain_424/module_data_out[1]
+ scanchain_424/module_data_out[2] scanchain_424/module_data_out[3] scanchain_424/module_data_out[4]
+ scanchain_424/module_data_out[5] scanchain_424/module_data_out[6] scanchain_424/module_data_out[7]
+ scanchain_424/scan_select_in scanchain_425/scan_select_in vccd1 vssd1 scanchain
Xscanchain_402 scanchain_402/clk_in scanchain_403/clk_in scanchain_402/data_in scanchain_403/data_in
+ scanchain_402/latch_enable_in scanchain_403/latch_enable_in scanchain_402/module_data_in[0]
+ scanchain_402/module_data_in[1] scanchain_402/module_data_in[2] scanchain_402/module_data_in[3]
+ scanchain_402/module_data_in[4] scanchain_402/module_data_in[5] scanchain_402/module_data_in[6]
+ scanchain_402/module_data_in[7] scanchain_402/module_data_out[0] scanchain_402/module_data_out[1]
+ scanchain_402/module_data_out[2] scanchain_402/module_data_out[3] scanchain_402/module_data_out[4]
+ scanchain_402/module_data_out[5] scanchain_402/module_data_out[6] scanchain_402/module_data_out[7]
+ scanchain_402/scan_select_in scanchain_403/scan_select_in vccd1 vssd1 scanchain
Xscanchain_413 scanchain_413/clk_in scanchain_414/clk_in scanchain_413/data_in scanchain_414/data_in
+ scanchain_413/latch_enable_in scanchain_414/latch_enable_in scanchain_413/module_data_in[0]
+ scanchain_413/module_data_in[1] scanchain_413/module_data_in[2] scanchain_413/module_data_in[3]
+ scanchain_413/module_data_in[4] scanchain_413/module_data_in[5] scanchain_413/module_data_in[6]
+ scanchain_413/module_data_in[7] scanchain_413/module_data_out[0] scanchain_413/module_data_out[1]
+ scanchain_413/module_data_out[2] scanchain_413/module_data_out[3] scanchain_413/module_data_out[4]
+ scanchain_413/module_data_out[5] scanchain_413/module_data_out[6] scanchain_413/module_data_out[7]
+ scanchain_413/scan_select_in scanchain_414/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_290 scanchain_290/module_data_in[0] scanchain_290/module_data_in[1]
+ scanchain_290/module_data_in[2] scanchain_290/module_data_in[3] scanchain_290/module_data_in[4]
+ scanchain_290/module_data_in[5] scanchain_290/module_data_in[6] scanchain_290/module_data_in[7]
+ scanchain_290/module_data_out[0] scanchain_290/module_data_out[1] scanchain_290/module_data_out[2]
+ scanchain_290/module_data_out[3] scanchain_290/module_data_out[4] scanchain_290/module_data_out[5]
+ scanchain_290/module_data_out[6] scanchain_290/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_287 scanchain_287/clk_in scanchain_288/clk_in scanchain_287/data_in scanchain_288/data_in
+ scanchain_287/latch_enable_in scanchain_288/latch_enable_in scanchain_287/module_data_in[0]
+ scanchain_287/module_data_in[1] scanchain_287/module_data_in[2] scanchain_287/module_data_in[3]
+ scanchain_287/module_data_in[4] scanchain_287/module_data_in[5] scanchain_287/module_data_in[6]
+ scanchain_287/module_data_in[7] scanchain_287/module_data_out[0] scanchain_287/module_data_out[1]
+ scanchain_287/module_data_out[2] scanchain_287/module_data_out[3] scanchain_287/module_data_out[4]
+ scanchain_287/module_data_out[5] scanchain_287/module_data_out[6] scanchain_287/module_data_out[7]
+ scanchain_287/scan_select_in scanchain_288/scan_select_in vccd1 vssd1 scanchain
Xscanchain_298 scanchain_298/clk_in scanchain_299/clk_in scanchain_298/data_in scanchain_299/data_in
+ scanchain_298/latch_enable_in scanchain_299/latch_enable_in scanchain_298/module_data_in[0]
+ scanchain_298/module_data_in[1] scanchain_298/module_data_in[2] scanchain_298/module_data_in[3]
+ scanchain_298/module_data_in[4] scanchain_298/module_data_in[5] scanchain_298/module_data_in[6]
+ scanchain_298/module_data_in[7] scanchain_298/module_data_out[0] scanchain_298/module_data_out[1]
+ scanchain_298/module_data_out[2] scanchain_298/module_data_out[3] scanchain_298/module_data_out[4]
+ scanchain_298/module_data_out[5] scanchain_298/module_data_out[6] scanchain_298/module_data_out[7]
+ scanchain_298/scan_select_in scanchain_299/scan_select_in vccd1 vssd1 scanchain
Xscanchain_276 scanchain_276/clk_in scanchain_277/clk_in scanchain_276/data_in scanchain_277/data_in
+ scanchain_276/latch_enable_in scanchain_277/latch_enable_in scanchain_276/module_data_in[0]
+ scanchain_276/module_data_in[1] scanchain_276/module_data_in[2] scanchain_276/module_data_in[3]
+ scanchain_276/module_data_in[4] scanchain_276/module_data_in[5] scanchain_276/module_data_in[6]
+ scanchain_276/module_data_in[7] scanchain_276/module_data_out[0] scanchain_276/module_data_out[1]
+ scanchain_276/module_data_out[2] scanchain_276/module_data_out[3] scanchain_276/module_data_out[4]
+ scanchain_276/module_data_out[5] scanchain_276/module_data_out[6] scanchain_276/module_data_out[7]
+ scanchain_276/scan_select_in scanchain_277/scan_select_in vccd1 vssd1 scanchain
Xscanchain_265 scanchain_265/clk_in scanchain_266/clk_in scanchain_265/data_in scanchain_266/data_in
+ scanchain_265/latch_enable_in scanchain_266/latch_enable_in scanchain_265/module_data_in[0]
+ scanchain_265/module_data_in[1] scanchain_265/module_data_in[2] scanchain_265/module_data_in[3]
+ scanchain_265/module_data_in[4] scanchain_265/module_data_in[5] scanchain_265/module_data_in[6]
+ scanchain_265/module_data_in[7] scanchain_265/module_data_out[0] scanchain_265/module_data_out[1]
+ scanchain_265/module_data_out[2] scanchain_265/module_data_out[3] scanchain_265/module_data_out[4]
+ scanchain_265/module_data_out[5] scanchain_265/module_data_out[6] scanchain_265/module_data_out[7]
+ scanchain_265/scan_select_in scanchain_266/scan_select_in vccd1 vssd1 scanchain
Xscanchain_254 scanchain_254/clk_in scanchain_255/clk_in scanchain_254/data_in scanchain_255/data_in
+ scanchain_254/latch_enable_in scanchain_255/latch_enable_in scanchain_254/module_data_in[0]
+ scanchain_254/module_data_in[1] scanchain_254/module_data_in[2] scanchain_254/module_data_in[3]
+ scanchain_254/module_data_in[4] scanchain_254/module_data_in[5] scanchain_254/module_data_in[6]
+ scanchain_254/module_data_in[7] scanchain_254/module_data_out[0] scanchain_254/module_data_out[1]
+ scanchain_254/module_data_out[2] scanchain_254/module_data_out[3] scanchain_254/module_data_out[4]
+ scanchain_254/module_data_out[5] scanchain_254/module_data_out[6] scanchain_254/module_data_out[7]
+ scanchain_254/scan_select_in scanchain_255/scan_select_in vccd1 vssd1 scanchain
Xscanchain_243 scanchain_243/clk_in scanchain_244/clk_in scanchain_243/data_in scanchain_244/data_in
+ scanchain_243/latch_enable_in scanchain_244/latch_enable_in scanchain_243/module_data_in[0]
+ scanchain_243/module_data_in[1] scanchain_243/module_data_in[2] scanchain_243/module_data_in[3]
+ scanchain_243/module_data_in[4] scanchain_243/module_data_in[5] scanchain_243/module_data_in[6]
+ scanchain_243/module_data_in[7] scanchain_243/module_data_out[0] scanchain_243/module_data_out[1]
+ scanchain_243/module_data_out[2] scanchain_243/module_data_out[3] scanchain_243/module_data_out[4]
+ scanchain_243/module_data_out[5] scanchain_243/module_data_out[6] scanchain_243/module_data_out[7]
+ scanchain_243/scan_select_in scanchain_244/scan_select_in vccd1 vssd1 scanchain
Xscanchain_232 scanchain_232/clk_in scanchain_233/clk_in scanchain_232/data_in scanchain_233/data_in
+ scanchain_232/latch_enable_in scanchain_233/latch_enable_in scanchain_232/module_data_in[0]
+ scanchain_232/module_data_in[1] scanchain_232/module_data_in[2] scanchain_232/module_data_in[3]
+ scanchain_232/module_data_in[4] scanchain_232/module_data_in[5] scanchain_232/module_data_in[6]
+ scanchain_232/module_data_in[7] scanchain_232/module_data_out[0] scanchain_232/module_data_out[1]
+ scanchain_232/module_data_out[2] scanchain_232/module_data_out[3] scanchain_232/module_data_out[4]
+ scanchain_232/module_data_out[5] scanchain_232/module_data_out[6] scanchain_232/module_data_out[7]
+ scanchain_232/scan_select_in scanchain_233/scan_select_in vccd1 vssd1 scanchain
Xscanchain_210 scanchain_210/clk_in scanchain_211/clk_in scanchain_210/data_in scanchain_211/data_in
+ scanchain_210/latch_enable_in scanchain_211/latch_enable_in scanchain_210/module_data_in[0]
+ scanchain_210/module_data_in[1] scanchain_210/module_data_in[2] scanchain_210/module_data_in[3]
+ scanchain_210/module_data_in[4] scanchain_210/module_data_in[5] scanchain_210/module_data_in[6]
+ scanchain_210/module_data_in[7] scanchain_210/module_data_out[0] scanchain_210/module_data_out[1]
+ scanchain_210/module_data_out[2] scanchain_210/module_data_out[3] scanchain_210/module_data_out[4]
+ scanchain_210/module_data_out[5] scanchain_210/module_data_out[6] scanchain_210/module_data_out[7]
+ scanchain_210/scan_select_in scanchain_211/scan_select_in vccd1 vssd1 scanchain
Xscanchain_221 scanchain_221/clk_in scanchain_222/clk_in scanchain_221/data_in scanchain_222/data_in
+ scanchain_221/latch_enable_in scanchain_222/latch_enable_in scanchain_221/module_data_in[0]
+ scanchain_221/module_data_in[1] scanchain_221/module_data_in[2] scanchain_221/module_data_in[3]
+ scanchain_221/module_data_in[4] scanchain_221/module_data_in[5] scanchain_221/module_data_in[6]
+ scanchain_221/module_data_in[7] scanchain_221/module_data_out[0] scanchain_221/module_data_out[1]
+ scanchain_221/module_data_out[2] scanchain_221/module_data_out[3] scanchain_221/module_data_out[4]
+ scanchain_221/module_data_out[5] scanchain_221/module_data_out[6] scanchain_221/module_data_out[7]
+ scanchain_221/scan_select_in scanchain_222/scan_select_in vccd1 vssd1 scanchain
Xscanchain_8 scanchain_8/clk_in scanchain_9/clk_in scanchain_8/data_in scanchain_9/data_in
+ scanchain_8/latch_enable_in scanchain_9/latch_enable_in aidan_McCoy_8/io_in[0] aidan_McCoy_8/io_in[1]
+ aidan_McCoy_8/io_in[2] aidan_McCoy_8/io_in[3] aidan_McCoy_8/io_in[4] aidan_McCoy_8/io_in[5]
+ aidan_McCoy_8/io_in[6] aidan_McCoy_8/io_in[7] aidan_McCoy_8/io_out[0] aidan_McCoy_8/io_out[1]
+ aidan_McCoy_8/io_out[2] aidan_McCoy_8/io_out[3] aidan_McCoy_8/io_out[4] aidan_McCoy_8/io_out[5]
+ aidan_McCoy_8/io_out[6] aidan_McCoy_8/io_out[7] scanchain_8/scan_select_in scanchain_9/scan_select_in
+ vccd1 vssd1 scanchain
Xuser_module_347594509754827347_19 scanchain_19/module_data_in[0] scanchain_19/module_data_in[1]
+ scanchain_19/module_data_in[2] scanchain_19/module_data_in[3] scanchain_19/module_data_in[4]
+ scanchain_19/module_data_in[5] scanchain_19/module_data_in[6] scanchain_19/module_data_in[7]
+ scanchain_19/module_data_out[0] scanchain_19/module_data_out[1] scanchain_19/module_data_out[2]
+ scanchain_19/module_data_out[3] scanchain_19/module_data_out[4] scanchain_19/module_data_out[5]
+ scanchain_19/module_data_out[6] scanchain_19/module_data_out[7] vccd1 vssd1 user_module_347594509754827347
Xscanchain_70 scanchain_70/clk_in scanchain_71/clk_in scanchain_70/data_in scanchain_71/data_in
+ scanchain_70/latch_enable_in scanchain_71/latch_enable_in scanchain_70/module_data_in[0]
+ scanchain_70/module_data_in[1] scanchain_70/module_data_in[2] scanchain_70/module_data_in[3]
+ scanchain_70/module_data_in[4] scanchain_70/module_data_in[5] scanchain_70/module_data_in[6]
+ scanchain_70/module_data_in[7] scanchain_70/module_data_out[0] scanchain_70/module_data_out[1]
+ scanchain_70/module_data_out[2] scanchain_70/module_data_out[3] scanchain_70/module_data_out[4]
+ scanchain_70/module_data_out[5] scanchain_70/module_data_out[6] scanchain_70/module_data_out[7]
+ scanchain_70/scan_select_in scanchain_71/scan_select_in vccd1 vssd1 scanchain
Xscanchain_81 scanchain_81/clk_in scanchain_82/clk_in scanchain_81/data_in scanchain_82/data_in
+ scanchain_81/latch_enable_in scanchain_82/latch_enable_in scanchain_81/module_data_in[0]
+ scanchain_81/module_data_in[1] scanchain_81/module_data_in[2] scanchain_81/module_data_in[3]
+ scanchain_81/module_data_in[4] scanchain_81/module_data_in[5] scanchain_81/module_data_in[6]
+ scanchain_81/module_data_in[7] scanchain_81/module_data_out[0] scanchain_81/module_data_out[1]
+ scanchain_81/module_data_out[2] scanchain_81/module_data_out[3] scanchain_81/module_data_out[4]
+ scanchain_81/module_data_out[5] scanchain_81/module_data_out[6] scanchain_81/module_data_out[7]
+ scanchain_81/scan_select_in scanchain_82/scan_select_in vccd1 vssd1 scanchain
Xscanchain_92 scanchain_92/clk_in scanchain_93/clk_in scanchain_92/data_in scanchain_93/data_in
+ scanchain_92/latch_enable_in scanchain_93/latch_enable_in scanchain_92/module_data_in[0]
+ scanchain_92/module_data_in[1] scanchain_92/module_data_in[2] scanchain_92/module_data_in[3]
+ scanchain_92/module_data_in[4] scanchain_92/module_data_in[5] scanchain_92/module_data_in[6]
+ scanchain_92/module_data_in[7] scanchain_92/module_data_out[0] scanchain_92/module_data_out[1]
+ scanchain_92/module_data_out[2] scanchain_92/module_data_out[3] scanchain_92/module_data_out[4]
+ scanchain_92/module_data_out[5] scanchain_92/module_data_out[6] scanchain_92/module_data_out[7]
+ scanchain_92/scan_select_in scanchain_93/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_108 scanchain_108/module_data_in[0] scanchain_108/module_data_in[1]
+ scanchain_108/module_data_in[2] scanchain_108/module_data_in[3] scanchain_108/module_data_in[4]
+ scanchain_108/module_data_in[5] scanchain_108/module_data_in[6] scanchain_108/module_data_in[7]
+ scanchain_108/module_data_out[0] scanchain_108/module_data_out[1] scanchain_108/module_data_out[2]
+ scanchain_108/module_data_out[3] scanchain_108/module_data_out[4] scanchain_108/module_data_out[5]
+ scanchain_108/module_data_out[6] scanchain_108/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_119 scanchain_119/module_data_in[0] scanchain_119/module_data_in[1]
+ scanchain_119/module_data_in[2] scanchain_119/module_data_in[3] scanchain_119/module_data_in[4]
+ scanchain_119/module_data_in[5] scanchain_119/module_data_in[6] scanchain_119/module_data_in[7]
+ scanchain_119/module_data_out[0] scanchain_119/module_data_out[1] scanchain_119/module_data_out[2]
+ scanchain_119/module_data_out[3] scanchain_119/module_data_out[4] scanchain_119/module_data_out[5]
+ scanchain_119/module_data_out[6] scanchain_119/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_472 scanchain_472/module_data_in[0] scanchain_472/module_data_in[1]
+ scanchain_472/module_data_in[2] scanchain_472/module_data_in[3] scanchain_472/module_data_in[4]
+ scanchain_472/module_data_in[5] scanchain_472/module_data_in[6] scanchain_472/module_data_in[7]
+ scanchain_472/module_data_out[0] scanchain_472/module_data_out[1] scanchain_472/module_data_out[2]
+ scanchain_472/module_data_out[3] scanchain_472/module_data_out[4] scanchain_472/module_data_out[5]
+ scanchain_472/module_data_out[6] scanchain_472/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_469 scanchain_469/clk_in scanchain_470/clk_in scanchain_469/data_in scanchain_470/data_in
+ scanchain_469/latch_enable_in scanchain_470/latch_enable_in scanchain_469/module_data_in[0]
+ scanchain_469/module_data_in[1] scanchain_469/module_data_in[2] scanchain_469/module_data_in[3]
+ scanchain_469/module_data_in[4] scanchain_469/module_data_in[5] scanchain_469/module_data_in[6]
+ scanchain_469/module_data_in[7] scanchain_469/module_data_out[0] scanchain_469/module_data_out[1]
+ scanchain_469/module_data_out[2] scanchain_469/module_data_out[3] scanchain_469/module_data_out[4]
+ scanchain_469/module_data_out[5] scanchain_469/module_data_out[6] scanchain_469/module_data_out[7]
+ scanchain_469/scan_select_in scanchain_470/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_461 scanchain_461/module_data_in[0] scanchain_461/module_data_in[1]
+ scanchain_461/module_data_in[2] scanchain_461/module_data_in[3] scanchain_461/module_data_in[4]
+ scanchain_461/module_data_in[5] scanchain_461/module_data_in[6] scanchain_461/module_data_in[7]
+ scanchain_461/module_data_out[0] scanchain_461/module_data_out[1] scanchain_461/module_data_out[2]
+ scanchain_461/module_data_out[3] scanchain_461/module_data_out[4] scanchain_461/module_data_out[5]
+ scanchain_461/module_data_out[6] scanchain_461/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_458 scanchain_458/clk_in scanchain_459/clk_in scanchain_458/data_in scanchain_459/data_in
+ scanchain_458/latch_enable_in scanchain_459/latch_enable_in scanchain_458/module_data_in[0]
+ scanchain_458/module_data_in[1] scanchain_458/module_data_in[2] scanchain_458/module_data_in[3]
+ scanchain_458/module_data_in[4] scanchain_458/module_data_in[5] scanchain_458/module_data_in[6]
+ scanchain_458/module_data_in[7] scanchain_458/module_data_out[0] scanchain_458/module_data_out[1]
+ scanchain_458/module_data_out[2] scanchain_458/module_data_out[3] scanchain_458/module_data_out[4]
+ scanchain_458/module_data_out[5] scanchain_458/module_data_out[6] scanchain_458/module_data_out[7]
+ scanchain_458/scan_select_in scanchain_459/scan_select_in vccd1 vssd1 scanchain
Xscanchain_436 scanchain_436/clk_in scanchain_437/clk_in scanchain_436/data_in scanchain_437/data_in
+ scanchain_436/latch_enable_in scanchain_437/latch_enable_in scanchain_436/module_data_in[0]
+ scanchain_436/module_data_in[1] scanchain_436/module_data_in[2] scanchain_436/module_data_in[3]
+ scanchain_436/module_data_in[4] scanchain_436/module_data_in[5] scanchain_436/module_data_in[6]
+ scanchain_436/module_data_in[7] scanchain_436/module_data_out[0] scanchain_436/module_data_out[1]
+ scanchain_436/module_data_out[2] scanchain_436/module_data_out[3] scanchain_436/module_data_out[4]
+ scanchain_436/module_data_out[5] scanchain_436/module_data_out[6] scanchain_436/module_data_out[7]
+ scanchain_436/scan_select_in scanchain_437/scan_select_in vccd1 vssd1 scanchain
Xscanchain_447 scanchain_447/clk_in scanchain_448/clk_in scanchain_447/data_in scanchain_448/data_in
+ scanchain_447/latch_enable_in scanchain_448/latch_enable_in scanchain_447/module_data_in[0]
+ scanchain_447/module_data_in[1] scanchain_447/module_data_in[2] scanchain_447/module_data_in[3]
+ scanchain_447/module_data_in[4] scanchain_447/module_data_in[5] scanchain_447/module_data_in[6]
+ scanchain_447/module_data_in[7] scanchain_447/module_data_out[0] scanchain_447/module_data_out[1]
+ scanchain_447/module_data_out[2] scanchain_447/module_data_out[3] scanchain_447/module_data_out[4]
+ scanchain_447/module_data_out[5] scanchain_447/module_data_out[6] scanchain_447/module_data_out[7]
+ scanchain_447/scan_select_in scanchain_448/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_450 scanchain_450/module_data_in[0] scanchain_450/module_data_in[1]
+ scanchain_450/module_data_in[2] scanchain_450/module_data_in[3] scanchain_450/module_data_in[4]
+ scanchain_450/module_data_in[5] scanchain_450/module_data_in[6] scanchain_450/module_data_in[7]
+ scanchain_450/module_data_out[0] scanchain_450/module_data_out[1] scanchain_450/module_data_out[2]
+ scanchain_450/module_data_out[3] scanchain_450/module_data_out[4] scanchain_450/module_data_out[5]
+ scanchain_450/module_data_out[6] scanchain_450/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_425 scanchain_425/clk_in scanchain_426/clk_in scanchain_425/data_in scanchain_426/data_in
+ scanchain_425/latch_enable_in scanchain_426/latch_enable_in scanchain_425/module_data_in[0]
+ scanchain_425/module_data_in[1] scanchain_425/module_data_in[2] scanchain_425/module_data_in[3]
+ scanchain_425/module_data_in[4] scanchain_425/module_data_in[5] scanchain_425/module_data_in[6]
+ scanchain_425/module_data_in[7] scanchain_425/module_data_out[0] scanchain_425/module_data_out[1]
+ scanchain_425/module_data_out[2] scanchain_425/module_data_out[3] scanchain_425/module_data_out[4]
+ scanchain_425/module_data_out[5] scanchain_425/module_data_out[6] scanchain_425/module_data_out[7]
+ scanchain_425/scan_select_in scanchain_426/scan_select_in vccd1 vssd1 scanchain
Xscanchain_403 scanchain_403/clk_in scanchain_404/clk_in scanchain_403/data_in scanchain_404/data_in
+ scanchain_403/latch_enable_in scanchain_404/latch_enable_in scanchain_403/module_data_in[0]
+ scanchain_403/module_data_in[1] scanchain_403/module_data_in[2] scanchain_403/module_data_in[3]
+ scanchain_403/module_data_in[4] scanchain_403/module_data_in[5] scanchain_403/module_data_in[6]
+ scanchain_403/module_data_in[7] scanchain_403/module_data_out[0] scanchain_403/module_data_out[1]
+ scanchain_403/module_data_out[2] scanchain_403/module_data_out[3] scanchain_403/module_data_out[4]
+ scanchain_403/module_data_out[5] scanchain_403/module_data_out[6] scanchain_403/module_data_out[7]
+ scanchain_403/scan_select_in scanchain_404/scan_select_in vccd1 vssd1 scanchain
Xscanchain_414 scanchain_414/clk_in scanchain_415/clk_in scanchain_414/data_in scanchain_415/data_in
+ scanchain_414/latch_enable_in scanchain_415/latch_enable_in scanchain_414/module_data_in[0]
+ scanchain_414/module_data_in[1] scanchain_414/module_data_in[2] scanchain_414/module_data_in[3]
+ scanchain_414/module_data_in[4] scanchain_414/module_data_in[5] scanchain_414/module_data_in[6]
+ scanchain_414/module_data_in[7] scanchain_414/module_data_out[0] scanchain_414/module_data_out[1]
+ scanchain_414/module_data_out[2] scanchain_414/module_data_out[3] scanchain_414/module_data_out[4]
+ scanchain_414/module_data_out[5] scanchain_414/module_data_out[6] scanchain_414/module_data_out[7]
+ scanchain_414/scan_select_in scanchain_415/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_291 scanchain_291/module_data_in[0] scanchain_291/module_data_in[1]
+ scanchain_291/module_data_in[2] scanchain_291/module_data_in[3] scanchain_291/module_data_in[4]
+ scanchain_291/module_data_in[5] scanchain_291/module_data_in[6] scanchain_291/module_data_in[7]
+ scanchain_291/module_data_out[0] scanchain_291/module_data_out[1] scanchain_291/module_data_out[2]
+ scanchain_291/module_data_out[3] scanchain_291/module_data_out[4] scanchain_291/module_data_out[5]
+ scanchain_291/module_data_out[6] scanchain_291/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_280 scanchain_280/module_data_in[0] scanchain_280/module_data_in[1]
+ scanchain_280/module_data_in[2] scanchain_280/module_data_in[3] scanchain_280/module_data_in[4]
+ scanchain_280/module_data_in[5] scanchain_280/module_data_in[6] scanchain_280/module_data_in[7]
+ scanchain_280/module_data_out[0] scanchain_280/module_data_out[1] scanchain_280/module_data_out[2]
+ scanchain_280/module_data_out[3] scanchain_280/module_data_out[4] scanchain_280/module_data_out[5]
+ scanchain_280/module_data_out[6] scanchain_280/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_288 scanchain_288/clk_in scanchain_289/clk_in scanchain_288/data_in scanchain_289/data_in
+ scanchain_288/latch_enable_in scanchain_289/latch_enable_in scanchain_288/module_data_in[0]
+ scanchain_288/module_data_in[1] scanchain_288/module_data_in[2] scanchain_288/module_data_in[3]
+ scanchain_288/module_data_in[4] scanchain_288/module_data_in[5] scanchain_288/module_data_in[6]
+ scanchain_288/module_data_in[7] scanchain_288/module_data_out[0] scanchain_288/module_data_out[1]
+ scanchain_288/module_data_out[2] scanchain_288/module_data_out[3] scanchain_288/module_data_out[4]
+ scanchain_288/module_data_out[5] scanchain_288/module_data_out[6] scanchain_288/module_data_out[7]
+ scanchain_288/scan_select_in scanchain_289/scan_select_in vccd1 vssd1 scanchain
Xscanchain_299 scanchain_299/clk_in scanchain_300/clk_in scanchain_299/data_in scanchain_300/data_in
+ scanchain_299/latch_enable_in scanchain_300/latch_enable_in scanchain_299/module_data_in[0]
+ scanchain_299/module_data_in[1] scanchain_299/module_data_in[2] scanchain_299/module_data_in[3]
+ scanchain_299/module_data_in[4] scanchain_299/module_data_in[5] scanchain_299/module_data_in[6]
+ scanchain_299/module_data_in[7] scanchain_299/module_data_out[0] scanchain_299/module_data_out[1]
+ scanchain_299/module_data_out[2] scanchain_299/module_data_out[3] scanchain_299/module_data_out[4]
+ scanchain_299/module_data_out[5] scanchain_299/module_data_out[6] scanchain_299/module_data_out[7]
+ scanchain_299/scan_select_in scanchain_300/scan_select_in vccd1 vssd1 scanchain
Xscanchain_277 scanchain_277/clk_in scanchain_278/clk_in scanchain_277/data_in scanchain_278/data_in
+ scanchain_277/latch_enable_in scanchain_278/latch_enable_in scanchain_277/module_data_in[0]
+ scanchain_277/module_data_in[1] scanchain_277/module_data_in[2] scanchain_277/module_data_in[3]
+ scanchain_277/module_data_in[4] scanchain_277/module_data_in[5] scanchain_277/module_data_in[6]
+ scanchain_277/module_data_in[7] scanchain_277/module_data_out[0] scanchain_277/module_data_out[1]
+ scanchain_277/module_data_out[2] scanchain_277/module_data_out[3] scanchain_277/module_data_out[4]
+ scanchain_277/module_data_out[5] scanchain_277/module_data_out[6] scanchain_277/module_data_out[7]
+ scanchain_277/scan_select_in scanchain_278/scan_select_in vccd1 vssd1 scanchain
Xscanchain_266 scanchain_266/clk_in scanchain_267/clk_in scanchain_266/data_in scanchain_267/data_in
+ scanchain_266/latch_enable_in scanchain_267/latch_enable_in scanchain_266/module_data_in[0]
+ scanchain_266/module_data_in[1] scanchain_266/module_data_in[2] scanchain_266/module_data_in[3]
+ scanchain_266/module_data_in[4] scanchain_266/module_data_in[5] scanchain_266/module_data_in[6]
+ scanchain_266/module_data_in[7] scanchain_266/module_data_out[0] scanchain_266/module_data_out[1]
+ scanchain_266/module_data_out[2] scanchain_266/module_data_out[3] scanchain_266/module_data_out[4]
+ scanchain_266/module_data_out[5] scanchain_266/module_data_out[6] scanchain_266/module_data_out[7]
+ scanchain_266/scan_select_in scanchain_267/scan_select_in vccd1 vssd1 scanchain
Xscanchain_255 scanchain_255/clk_in scanchain_256/clk_in scanchain_255/data_in scanchain_256/data_in
+ scanchain_255/latch_enable_in scanchain_256/latch_enable_in scanchain_255/module_data_in[0]
+ scanchain_255/module_data_in[1] scanchain_255/module_data_in[2] scanchain_255/module_data_in[3]
+ scanchain_255/module_data_in[4] scanchain_255/module_data_in[5] scanchain_255/module_data_in[6]
+ scanchain_255/module_data_in[7] scanchain_255/module_data_out[0] scanchain_255/module_data_out[1]
+ scanchain_255/module_data_out[2] scanchain_255/module_data_out[3] scanchain_255/module_data_out[4]
+ scanchain_255/module_data_out[5] scanchain_255/module_data_out[6] scanchain_255/module_data_out[7]
+ scanchain_255/scan_select_in scanchain_256/scan_select_in vccd1 vssd1 scanchain
Xscanchain_244 scanchain_244/clk_in scanchain_245/clk_in scanchain_244/data_in scanchain_245/data_in
+ scanchain_244/latch_enable_in scanchain_245/latch_enable_in scanchain_244/module_data_in[0]
+ scanchain_244/module_data_in[1] scanchain_244/module_data_in[2] scanchain_244/module_data_in[3]
+ scanchain_244/module_data_in[4] scanchain_244/module_data_in[5] scanchain_244/module_data_in[6]
+ scanchain_244/module_data_in[7] scanchain_244/module_data_out[0] scanchain_244/module_data_out[1]
+ scanchain_244/module_data_out[2] scanchain_244/module_data_out[3] scanchain_244/module_data_out[4]
+ scanchain_244/module_data_out[5] scanchain_244/module_data_out[6] scanchain_244/module_data_out[7]
+ scanchain_244/scan_select_in scanchain_245/scan_select_in vccd1 vssd1 scanchain
Xscanchain_233 scanchain_233/clk_in scanchain_234/clk_in scanchain_233/data_in scanchain_234/data_in
+ scanchain_233/latch_enable_in scanchain_234/latch_enable_in scanchain_233/module_data_in[0]
+ scanchain_233/module_data_in[1] scanchain_233/module_data_in[2] scanchain_233/module_data_in[3]
+ scanchain_233/module_data_in[4] scanchain_233/module_data_in[5] scanchain_233/module_data_in[6]
+ scanchain_233/module_data_in[7] scanchain_233/module_data_out[0] scanchain_233/module_data_out[1]
+ scanchain_233/module_data_out[2] scanchain_233/module_data_out[3] scanchain_233/module_data_out[4]
+ scanchain_233/module_data_out[5] scanchain_233/module_data_out[6] scanchain_233/module_data_out[7]
+ scanchain_233/scan_select_in scanchain_234/scan_select_in vccd1 vssd1 scanchain
Xscanchain_211 scanchain_211/clk_in scanchain_212/clk_in scanchain_211/data_in scanchain_212/data_in
+ scanchain_211/latch_enable_in scanchain_212/latch_enable_in scanchain_211/module_data_in[0]
+ scanchain_211/module_data_in[1] scanchain_211/module_data_in[2] scanchain_211/module_data_in[3]
+ scanchain_211/module_data_in[4] scanchain_211/module_data_in[5] scanchain_211/module_data_in[6]
+ scanchain_211/module_data_in[7] scanchain_211/module_data_out[0] scanchain_211/module_data_out[1]
+ scanchain_211/module_data_out[2] scanchain_211/module_data_out[3] scanchain_211/module_data_out[4]
+ scanchain_211/module_data_out[5] scanchain_211/module_data_out[6] scanchain_211/module_data_out[7]
+ scanchain_211/scan_select_in scanchain_212/scan_select_in vccd1 vssd1 scanchain
Xscanchain_222 scanchain_222/clk_in scanchain_223/clk_in scanchain_222/data_in scanchain_223/data_in
+ scanchain_222/latch_enable_in scanchain_223/latch_enable_in scanchain_222/module_data_in[0]
+ scanchain_222/module_data_in[1] scanchain_222/module_data_in[2] scanchain_222/module_data_in[3]
+ scanchain_222/module_data_in[4] scanchain_222/module_data_in[5] scanchain_222/module_data_in[6]
+ scanchain_222/module_data_in[7] scanchain_222/module_data_out[0] scanchain_222/module_data_out[1]
+ scanchain_222/module_data_out[2] scanchain_222/module_data_out[3] scanchain_222/module_data_out[4]
+ scanchain_222/module_data_out[5] scanchain_222/module_data_out[6] scanchain_222/module_data_out[7]
+ scanchain_222/scan_select_in scanchain_223/scan_select_in vccd1 vssd1 scanchain
Xscanchain_200 scanchain_200/clk_in scanchain_201/clk_in scanchain_200/data_in scanchain_201/data_in
+ scanchain_200/latch_enable_in scanchain_201/latch_enable_in scanchain_200/module_data_in[0]
+ scanchain_200/module_data_in[1] scanchain_200/module_data_in[2] scanchain_200/module_data_in[3]
+ scanchain_200/module_data_in[4] scanchain_200/module_data_in[5] scanchain_200/module_data_in[6]
+ scanchain_200/module_data_in[7] scanchain_200/module_data_out[0] scanchain_200/module_data_out[1]
+ scanchain_200/module_data_out[2] scanchain_200/module_data_out[3] scanchain_200/module_data_out[4]
+ scanchain_200/module_data_out[5] scanchain_200/module_data_out[6] scanchain_200/module_data_out[7]
+ scanchain_200/scan_select_in scanchain_201/scan_select_in vccd1 vssd1 scanchain
Xscanchain_9 scanchain_9/clk_in scanchain_9/clk_out scanchain_9/data_in scanchain_9/data_out
+ scanchain_9/latch_enable_in scanchain_9/latch_enable_out scanchain_9/module_data_in[0]
+ scanchain_9/module_data_in[1] scanchain_9/module_data_in[2] scanchain_9/module_data_in[3]
+ scanchain_9/module_data_in[4] scanchain_9/module_data_in[5] scanchain_9/module_data_in[6]
+ scanchain_9/module_data_in[7] scanchain_9/module_data_out[0] scanchain_9/module_data_out[1]
+ scanchain_9/module_data_out[2] scanchain_9/module_data_out[3] scanchain_9/module_data_out[4]
+ scanchain_9/module_data_out[5] scanchain_9/module_data_out[6] scanchain_9/module_data_out[7]
+ scanchain_9/scan_select_in scanchain_9/scan_select_out vccd1 vssd1 scanchain
Xs4ga_6 s4ga_6/io_in[0] s4ga_6/io_in[1] s4ga_6/io_in[2] s4ga_6/io_in[3] s4ga_6/io_in[4]
+ s4ga_6/io_in[5] s4ga_6/io_in[6] s4ga_6/io_in[7] s4ga_6/io_out[0] s4ga_6/io_out[1]
+ s4ga_6/io_out[2] s4ga_6/io_out[3] s4ga_6/io_out[4] s4ga_6/io_out[5] s4ga_6/io_out[6]
+ s4ga_6/io_out[7] vccd1 vssd1 s4ga
Xscanchain_71 scanchain_71/clk_in scanchain_72/clk_in scanchain_71/data_in scanchain_72/data_in
+ scanchain_71/latch_enable_in scanchain_72/latch_enable_in scanchain_71/module_data_in[0]
+ scanchain_71/module_data_in[1] scanchain_71/module_data_in[2] scanchain_71/module_data_in[3]
+ scanchain_71/module_data_in[4] scanchain_71/module_data_in[5] scanchain_71/module_data_in[6]
+ scanchain_71/module_data_in[7] scanchain_71/module_data_out[0] scanchain_71/module_data_out[1]
+ scanchain_71/module_data_out[2] scanchain_71/module_data_out[3] scanchain_71/module_data_out[4]
+ scanchain_71/module_data_out[5] scanchain_71/module_data_out[6] scanchain_71/module_data_out[7]
+ scanchain_71/scan_select_in scanchain_72/scan_select_in vccd1 vssd1 scanchain
Xscanchain_60 scanchain_60/clk_in scanchain_61/clk_in scanchain_60/data_in scanchain_61/data_in
+ scanchain_60/latch_enable_in scanchain_61/latch_enable_in scanchain_60/module_data_in[0]
+ scanchain_60/module_data_in[1] scanchain_60/module_data_in[2] scanchain_60/module_data_in[3]
+ scanchain_60/module_data_in[4] scanchain_60/module_data_in[5] scanchain_60/module_data_in[6]
+ scanchain_60/module_data_in[7] scanchain_60/module_data_out[0] scanchain_60/module_data_out[1]
+ scanchain_60/module_data_out[2] scanchain_60/module_data_out[3] scanchain_60/module_data_out[4]
+ scanchain_60/module_data_out[5] scanchain_60/module_data_out[6] scanchain_60/module_data_out[7]
+ scanchain_60/scan_select_in scanchain_61/scan_select_in vccd1 vssd1 scanchain
Xscanchain_82 scanchain_82/clk_in scanchain_83/clk_in scanchain_82/data_in scanchain_83/data_in
+ scanchain_82/latch_enable_in scanchain_83/latch_enable_in scanchain_82/module_data_in[0]
+ scanchain_82/module_data_in[1] scanchain_82/module_data_in[2] scanchain_82/module_data_in[3]
+ scanchain_82/module_data_in[4] scanchain_82/module_data_in[5] scanchain_82/module_data_in[6]
+ scanchain_82/module_data_in[7] scanchain_82/module_data_out[0] scanchain_82/module_data_out[1]
+ scanchain_82/module_data_out[2] scanchain_82/module_data_out[3] scanchain_82/module_data_out[4]
+ scanchain_82/module_data_out[5] scanchain_82/module_data_out[6] scanchain_82/module_data_out[7]
+ scanchain_82/scan_select_in scanchain_83/scan_select_in vccd1 vssd1 scanchain
Xscanchain_93 scanchain_93/clk_in scanchain_94/clk_in scanchain_93/data_in scanchain_94/data_in
+ scanchain_93/latch_enable_in scanchain_94/latch_enable_in scanchain_93/module_data_in[0]
+ scanchain_93/module_data_in[1] scanchain_93/module_data_in[2] scanchain_93/module_data_in[3]
+ scanchain_93/module_data_in[4] scanchain_93/module_data_in[5] scanchain_93/module_data_in[6]
+ scanchain_93/module_data_in[7] scanchain_93/module_data_out[0] scanchain_93/module_data_out[1]
+ scanchain_93/module_data_out[2] scanchain_93/module_data_out[3] scanchain_93/module_data_out[4]
+ scanchain_93/module_data_out[5] scanchain_93/module_data_out[6] scanchain_93/module_data_out[7]
+ scanchain_93/scan_select_in scanchain_94/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_109 scanchain_109/module_data_in[0] scanchain_109/module_data_in[1]
+ scanchain_109/module_data_in[2] scanchain_109/module_data_in[3] scanchain_109/module_data_in[4]
+ scanchain_109/module_data_in[5] scanchain_109/module_data_in[6] scanchain_109/module_data_in[7]
+ scanchain_109/module_data_out[0] scanchain_109/module_data_out[1] scanchain_109/module_data_out[2]
+ scanchain_109/module_data_out[3] scanchain_109/module_data_out[4] scanchain_109/module_data_out[5]
+ scanchain_109/module_data_out[6] scanchain_109/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_462 scanchain_462/module_data_in[0] scanchain_462/module_data_in[1]
+ scanchain_462/module_data_in[2] scanchain_462/module_data_in[3] scanchain_462/module_data_in[4]
+ scanchain_462/module_data_in[5] scanchain_462/module_data_in[6] scanchain_462/module_data_in[7]
+ scanchain_462/module_data_out[0] scanchain_462/module_data_out[1] scanchain_462/module_data_out[2]
+ scanchain_462/module_data_out[3] scanchain_462/module_data_out[4] scanchain_462/module_data_out[5]
+ scanchain_462/module_data_out[6] scanchain_462/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_459 scanchain_459/clk_in scanchain_460/clk_in scanchain_459/data_in scanchain_460/data_in
+ scanchain_459/latch_enable_in scanchain_460/latch_enable_in scanchain_459/module_data_in[0]
+ scanchain_459/module_data_in[1] scanchain_459/module_data_in[2] scanchain_459/module_data_in[3]
+ scanchain_459/module_data_in[4] scanchain_459/module_data_in[5] scanchain_459/module_data_in[6]
+ scanchain_459/module_data_in[7] scanchain_459/module_data_out[0] scanchain_459/module_data_out[1]
+ scanchain_459/module_data_out[2] scanchain_459/module_data_out[3] scanchain_459/module_data_out[4]
+ scanchain_459/module_data_out[5] scanchain_459/module_data_out[6] scanchain_459/module_data_out[7]
+ scanchain_459/scan_select_in scanchain_460/scan_select_in vccd1 vssd1 scanchain
Xscanchain_437 scanchain_437/clk_in scanchain_438/clk_in scanchain_437/data_in scanchain_438/data_in
+ scanchain_437/latch_enable_in scanchain_438/latch_enable_in scanchain_437/module_data_in[0]
+ scanchain_437/module_data_in[1] scanchain_437/module_data_in[2] scanchain_437/module_data_in[3]
+ scanchain_437/module_data_in[4] scanchain_437/module_data_in[5] scanchain_437/module_data_in[6]
+ scanchain_437/module_data_in[7] scanchain_437/module_data_out[0] scanchain_437/module_data_out[1]
+ scanchain_437/module_data_out[2] scanchain_437/module_data_out[3] scanchain_437/module_data_out[4]
+ scanchain_437/module_data_out[5] scanchain_437/module_data_out[6] scanchain_437/module_data_out[7]
+ scanchain_437/scan_select_in scanchain_438/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_440 scanchain_440/module_data_in[0] scanchain_440/module_data_in[1]
+ scanchain_440/module_data_in[2] scanchain_440/module_data_in[3] scanchain_440/module_data_in[4]
+ scanchain_440/module_data_in[5] scanchain_440/module_data_in[6] scanchain_440/module_data_in[7]
+ scanchain_440/module_data_out[0] scanchain_440/module_data_out[1] scanchain_440/module_data_out[2]
+ scanchain_440/module_data_out[3] scanchain_440/module_data_out[4] scanchain_440/module_data_out[5]
+ scanchain_440/module_data_out[6] scanchain_440/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_448 scanchain_448/clk_in scanchain_449/clk_in scanchain_448/data_in scanchain_449/data_in
+ scanchain_448/latch_enable_in scanchain_449/latch_enable_in scanchain_448/module_data_in[0]
+ scanchain_448/module_data_in[1] scanchain_448/module_data_in[2] scanchain_448/module_data_in[3]
+ scanchain_448/module_data_in[4] scanchain_448/module_data_in[5] scanchain_448/module_data_in[6]
+ scanchain_448/module_data_in[7] scanchain_448/module_data_out[0] scanchain_448/module_data_out[1]
+ scanchain_448/module_data_out[2] scanchain_448/module_data_out[3] scanchain_448/module_data_out[4]
+ scanchain_448/module_data_out[5] scanchain_448/module_data_out[6] scanchain_448/module_data_out[7]
+ scanchain_448/scan_select_in scanchain_449/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_451 scanchain_451/module_data_in[0] scanchain_451/module_data_in[1]
+ scanchain_451/module_data_in[2] scanchain_451/module_data_in[3] scanchain_451/module_data_in[4]
+ scanchain_451/module_data_in[5] scanchain_451/module_data_in[6] scanchain_451/module_data_in[7]
+ scanchain_451/module_data_out[0] scanchain_451/module_data_out[1] scanchain_451/module_data_out[2]
+ scanchain_451/module_data_out[3] scanchain_451/module_data_out[4] scanchain_451/module_data_out[5]
+ scanchain_451/module_data_out[6] scanchain_451/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_426 scanchain_426/clk_in scanchain_427/clk_in scanchain_426/data_in scanchain_427/data_in
+ scanchain_426/latch_enable_in scanchain_427/latch_enable_in scanchain_426/module_data_in[0]
+ scanchain_426/module_data_in[1] scanchain_426/module_data_in[2] scanchain_426/module_data_in[3]
+ scanchain_426/module_data_in[4] scanchain_426/module_data_in[5] scanchain_426/module_data_in[6]
+ scanchain_426/module_data_in[7] scanchain_426/module_data_out[0] scanchain_426/module_data_out[1]
+ scanchain_426/module_data_out[2] scanchain_426/module_data_out[3] scanchain_426/module_data_out[4]
+ scanchain_426/module_data_out[5] scanchain_426/module_data_out[6] scanchain_426/module_data_out[7]
+ scanchain_426/scan_select_in scanchain_427/scan_select_in vccd1 vssd1 scanchain
Xscanchain_404 scanchain_404/clk_in scanchain_405/clk_in scanchain_404/data_in scanchain_405/data_in
+ scanchain_404/latch_enable_in scanchain_405/latch_enable_in scanchain_404/module_data_in[0]
+ scanchain_404/module_data_in[1] scanchain_404/module_data_in[2] scanchain_404/module_data_in[3]
+ scanchain_404/module_data_in[4] scanchain_404/module_data_in[5] scanchain_404/module_data_in[6]
+ scanchain_404/module_data_in[7] scanchain_404/module_data_out[0] scanchain_404/module_data_out[1]
+ scanchain_404/module_data_out[2] scanchain_404/module_data_out[3] scanchain_404/module_data_out[4]
+ scanchain_404/module_data_out[5] scanchain_404/module_data_out[6] scanchain_404/module_data_out[7]
+ scanchain_404/scan_select_in scanchain_405/scan_select_in vccd1 vssd1 scanchain
Xscanchain_415 scanchain_415/clk_in scanchain_416/clk_in scanchain_415/data_in scanchain_416/data_in
+ scanchain_415/latch_enable_in scanchain_416/latch_enable_in scanchain_415/module_data_in[0]
+ scanchain_415/module_data_in[1] scanchain_415/module_data_in[2] scanchain_415/module_data_in[3]
+ scanchain_415/module_data_in[4] scanchain_415/module_data_in[5] scanchain_415/module_data_in[6]
+ scanchain_415/module_data_in[7] scanchain_415/module_data_out[0] scanchain_415/module_data_out[1]
+ scanchain_415/module_data_out[2] scanchain_415/module_data_out[3] scanchain_415/module_data_out[4]
+ scanchain_415/module_data_out[5] scanchain_415/module_data_out[6] scanchain_415/module_data_out[7]
+ scanchain_415/scan_select_in scanchain_416/scan_select_in vccd1 vssd1 scanchain
Xasic_multiplier_wrapper_23 scanchain_23/module_data_in[0] scanchain_23/module_data_in[1]
+ scanchain_23/module_data_in[2] scanchain_23/module_data_in[3] scanchain_23/module_data_in[4]
+ scanchain_23/module_data_in[5] scanchain_23/module_data_in[6] scanchain_23/module_data_in[7]
+ scanchain_23/module_data_out[0] scanchain_23/module_data_out[1] scanchain_23/module_data_out[2]
+ scanchain_23/module_data_out[3] scanchain_23/module_data_out[4] scanchain_23/module_data_out[5]
+ scanchain_23/module_data_out[6] scanchain_23/module_data_out[7] vccd1 vssd1 asic_multiplier_wrapper
Xscanchain_289 scanchain_289/clk_in scanchain_290/clk_in scanchain_289/data_in scanchain_290/data_in
+ scanchain_289/latch_enable_in scanchain_290/latch_enable_in scanchain_289/module_data_in[0]
+ scanchain_289/module_data_in[1] scanchain_289/module_data_in[2] scanchain_289/module_data_in[3]
+ scanchain_289/module_data_in[4] scanchain_289/module_data_in[5] scanchain_289/module_data_in[6]
+ scanchain_289/module_data_in[7] scanchain_289/module_data_out[0] scanchain_289/module_data_out[1]
+ scanchain_289/module_data_out[2] scanchain_289/module_data_out[3] scanchain_289/module_data_out[4]
+ scanchain_289/module_data_out[5] scanchain_289/module_data_out[6] scanchain_289/module_data_out[7]
+ scanchain_289/scan_select_in scanchain_290/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_292 scanchain_292/module_data_in[0] scanchain_292/module_data_in[1]
+ scanchain_292/module_data_in[2] scanchain_292/module_data_in[3] scanchain_292/module_data_in[4]
+ scanchain_292/module_data_in[5] scanchain_292/module_data_in[6] scanchain_292/module_data_in[7]
+ scanchain_292/module_data_out[0] scanchain_292/module_data_out[1] scanchain_292/module_data_out[2]
+ scanchain_292/module_data_out[3] scanchain_292/module_data_out[4] scanchain_292/module_data_out[5]
+ scanchain_292/module_data_out[6] scanchain_292/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_281 scanchain_281/module_data_in[0] scanchain_281/module_data_in[1]
+ scanchain_281/module_data_in[2] scanchain_281/module_data_in[3] scanchain_281/module_data_in[4]
+ scanchain_281/module_data_in[5] scanchain_281/module_data_in[6] scanchain_281/module_data_in[7]
+ scanchain_281/module_data_out[0] scanchain_281/module_data_out[1] scanchain_281/module_data_out[2]
+ scanchain_281/module_data_out[3] scanchain_281/module_data_out[4] scanchain_281/module_data_out[5]
+ scanchain_281/module_data_out[6] scanchain_281/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_278 scanchain_278/clk_in scanchain_279/clk_in scanchain_278/data_in scanchain_279/data_in
+ scanchain_278/latch_enable_in scanchain_279/latch_enable_in scanchain_278/module_data_in[0]
+ scanchain_278/module_data_in[1] scanchain_278/module_data_in[2] scanchain_278/module_data_in[3]
+ scanchain_278/module_data_in[4] scanchain_278/module_data_in[5] scanchain_278/module_data_in[6]
+ scanchain_278/module_data_in[7] scanchain_278/module_data_out[0] scanchain_278/module_data_out[1]
+ scanchain_278/module_data_out[2] scanchain_278/module_data_out[3] scanchain_278/module_data_out[4]
+ scanchain_278/module_data_out[5] scanchain_278/module_data_out[6] scanchain_278/module_data_out[7]
+ scanchain_278/scan_select_in scanchain_279/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_270 scanchain_270/module_data_in[0] scanchain_270/module_data_in[1]
+ scanchain_270/module_data_in[2] scanchain_270/module_data_in[3] scanchain_270/module_data_in[4]
+ scanchain_270/module_data_in[5] scanchain_270/module_data_in[6] scanchain_270/module_data_in[7]
+ scanchain_270/module_data_out[0] scanchain_270/module_data_out[1] scanchain_270/module_data_out[2]
+ scanchain_270/module_data_out[3] scanchain_270/module_data_out[4] scanchain_270/module_data_out[5]
+ scanchain_270/module_data_out[6] scanchain_270/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_267 scanchain_267/clk_in scanchain_268/clk_in scanchain_267/data_in scanchain_268/data_in
+ scanchain_267/latch_enable_in scanchain_268/latch_enable_in scanchain_267/module_data_in[0]
+ scanchain_267/module_data_in[1] scanchain_267/module_data_in[2] scanchain_267/module_data_in[3]
+ scanchain_267/module_data_in[4] scanchain_267/module_data_in[5] scanchain_267/module_data_in[6]
+ scanchain_267/module_data_in[7] scanchain_267/module_data_out[0] scanchain_267/module_data_out[1]
+ scanchain_267/module_data_out[2] scanchain_267/module_data_out[3] scanchain_267/module_data_out[4]
+ scanchain_267/module_data_out[5] scanchain_267/module_data_out[6] scanchain_267/module_data_out[7]
+ scanchain_267/scan_select_in scanchain_268/scan_select_in vccd1 vssd1 scanchain
Xscanchain_245 scanchain_245/clk_in scanchain_246/clk_in scanchain_245/data_in scanchain_246/data_in
+ scanchain_245/latch_enable_in scanchain_246/latch_enable_in scanchain_245/module_data_in[0]
+ scanchain_245/module_data_in[1] scanchain_245/module_data_in[2] scanchain_245/module_data_in[3]
+ scanchain_245/module_data_in[4] scanchain_245/module_data_in[5] scanchain_245/module_data_in[6]
+ scanchain_245/module_data_in[7] scanchain_245/module_data_out[0] scanchain_245/module_data_out[1]
+ scanchain_245/module_data_out[2] scanchain_245/module_data_out[3] scanchain_245/module_data_out[4]
+ scanchain_245/module_data_out[5] scanchain_245/module_data_out[6] scanchain_245/module_data_out[7]
+ scanchain_245/scan_select_in scanchain_246/scan_select_in vccd1 vssd1 scanchain
Xscanchain_256 scanchain_256/clk_in scanchain_257/clk_in scanchain_256/data_in scanchain_257/data_in
+ scanchain_256/latch_enable_in scanchain_257/latch_enable_in scanchain_256/module_data_in[0]
+ scanchain_256/module_data_in[1] scanchain_256/module_data_in[2] scanchain_256/module_data_in[3]
+ scanchain_256/module_data_in[4] scanchain_256/module_data_in[5] scanchain_256/module_data_in[6]
+ scanchain_256/module_data_in[7] scanchain_256/module_data_out[0] scanchain_256/module_data_out[1]
+ scanchain_256/module_data_out[2] scanchain_256/module_data_out[3] scanchain_256/module_data_out[4]
+ scanchain_256/module_data_out[5] scanchain_256/module_data_out[6] scanchain_256/module_data_out[7]
+ scanchain_256/scan_select_in scanchain_257/scan_select_in vccd1 vssd1 scanchain
Xscanchain_234 scanchain_234/clk_in scanchain_235/clk_in scanchain_234/data_in scanchain_235/data_in
+ scanchain_234/latch_enable_in scanchain_235/latch_enable_in scanchain_234/module_data_in[0]
+ scanchain_234/module_data_in[1] scanchain_234/module_data_in[2] scanchain_234/module_data_in[3]
+ scanchain_234/module_data_in[4] scanchain_234/module_data_in[5] scanchain_234/module_data_in[6]
+ scanchain_234/module_data_in[7] scanchain_234/module_data_out[0] scanchain_234/module_data_out[1]
+ scanchain_234/module_data_out[2] scanchain_234/module_data_out[3] scanchain_234/module_data_out[4]
+ scanchain_234/module_data_out[5] scanchain_234/module_data_out[6] scanchain_234/module_data_out[7]
+ scanchain_234/scan_select_in scanchain_235/scan_select_in vccd1 vssd1 scanchain
Xscanchain_212 scanchain_212/clk_in scanchain_213/clk_in scanchain_212/data_in scanchain_213/data_in
+ scanchain_212/latch_enable_in scanchain_213/latch_enable_in scanchain_212/module_data_in[0]
+ scanchain_212/module_data_in[1] scanchain_212/module_data_in[2] scanchain_212/module_data_in[3]
+ scanchain_212/module_data_in[4] scanchain_212/module_data_in[5] scanchain_212/module_data_in[6]
+ scanchain_212/module_data_in[7] scanchain_212/module_data_out[0] scanchain_212/module_data_out[1]
+ scanchain_212/module_data_out[2] scanchain_212/module_data_out[3] scanchain_212/module_data_out[4]
+ scanchain_212/module_data_out[5] scanchain_212/module_data_out[6] scanchain_212/module_data_out[7]
+ scanchain_212/scan_select_in scanchain_213/scan_select_in vccd1 vssd1 scanchain
Xscanchain_223 scanchain_223/clk_in scanchain_224/clk_in scanchain_223/data_in scanchain_224/data_in
+ scanchain_223/latch_enable_in scanchain_224/latch_enable_in scanchain_223/module_data_in[0]
+ scanchain_223/module_data_in[1] scanchain_223/module_data_in[2] scanchain_223/module_data_in[3]
+ scanchain_223/module_data_in[4] scanchain_223/module_data_in[5] scanchain_223/module_data_in[6]
+ scanchain_223/module_data_in[7] scanchain_223/module_data_out[0] scanchain_223/module_data_out[1]
+ scanchain_223/module_data_out[2] scanchain_223/module_data_out[3] scanchain_223/module_data_out[4]
+ scanchain_223/module_data_out[5] scanchain_223/module_data_out[6] scanchain_223/module_data_out[7]
+ scanchain_223/scan_select_in scanchain_224/scan_select_in vccd1 vssd1 scanchain
Xscanchain_201 scanchain_201/clk_in scanchain_202/clk_in scanchain_201/data_in scanchain_202/data_in
+ scanchain_201/latch_enable_in scanchain_202/latch_enable_in scanchain_201/module_data_in[0]
+ scanchain_201/module_data_in[1] scanchain_201/module_data_in[2] scanchain_201/module_data_in[3]
+ scanchain_201/module_data_in[4] scanchain_201/module_data_in[5] scanchain_201/module_data_in[6]
+ scanchain_201/module_data_in[7] scanchain_201/module_data_out[0] scanchain_201/module_data_out[1]
+ scanchain_201/module_data_out[2] scanchain_201/module_data_out[3] scanchain_201/module_data_out[4]
+ scanchain_201/module_data_out[5] scanchain_201/module_data_out[6] scanchain_201/module_data_out[7]
+ scanchain_201/scan_select_in scanchain_202/scan_select_in vccd1 vssd1 scanchain
Xloxodes_sequencer_4 loxodes_sequencer_4/io_in[0] loxodes_sequencer_4/io_in[1] loxodes_sequencer_4/io_in[2]
+ loxodes_sequencer_4/io_in[3] loxodes_sequencer_4/io_in[4] loxodes_sequencer_4/io_in[5]
+ loxodes_sequencer_4/io_in[6] loxodes_sequencer_4/io_in[7] loxodes_sequencer_4/io_out[0]
+ loxodes_sequencer_4/io_out[1] loxodes_sequencer_4/io_out[2] loxodes_sequencer_4/io_out[3]
+ loxodes_sequencer_4/io_out[4] loxodes_sequencer_4/io_out[5] loxodes_sequencer_4/io_out[6]
+ loxodes_sequencer_4/io_out[7] vccd1 vssd1 loxodes_sequencer
Xuser_module_339501025136214612_90 scanchain_90/module_data_in[0] scanchain_90/module_data_in[1]
+ scanchain_90/module_data_in[2] scanchain_90/module_data_in[3] scanchain_90/module_data_in[4]
+ scanchain_90/module_data_in[5] scanchain_90/module_data_in[6] scanchain_90/module_data_in[7]
+ scanchain_90/module_data_out[0] scanchain_90/module_data_out[1] scanchain_90/module_data_out[2]
+ scanchain_90/module_data_out[3] scanchain_90/module_data_out[4] scanchain_90/module_data_out[5]
+ scanchain_90/module_data_out[6] scanchain_90/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_50 scanchain_50/clk_in scanchain_51/clk_in scanchain_50/data_in scanchain_51/data_in
+ scanchain_50/latch_enable_in scanchain_51/latch_enable_in scanchain_50/module_data_in[0]
+ scanchain_50/module_data_in[1] scanchain_50/module_data_in[2] scanchain_50/module_data_in[3]
+ scanchain_50/module_data_in[4] scanchain_50/module_data_in[5] scanchain_50/module_data_in[6]
+ scanchain_50/module_data_in[7] scanchain_50/module_data_out[0] scanchain_50/module_data_out[1]
+ scanchain_50/module_data_out[2] scanchain_50/module_data_out[3] scanchain_50/module_data_out[4]
+ scanchain_50/module_data_out[5] scanchain_50/module_data_out[6] scanchain_50/module_data_out[7]
+ scanchain_50/scan_select_in scanchain_51/scan_select_in vccd1 vssd1 scanchain
Xscanchain_72 scanchain_72/clk_in scanchain_73/clk_in scanchain_72/data_in scanchain_73/data_in
+ scanchain_72/latch_enable_in scanchain_73/latch_enable_in scanchain_72/module_data_in[0]
+ scanchain_72/module_data_in[1] scanchain_72/module_data_in[2] scanchain_72/module_data_in[3]
+ scanchain_72/module_data_in[4] scanchain_72/module_data_in[5] scanchain_72/module_data_in[6]
+ scanchain_72/module_data_in[7] scanchain_72/module_data_out[0] scanchain_72/module_data_out[1]
+ scanchain_72/module_data_out[2] scanchain_72/module_data_out[3] scanchain_72/module_data_out[4]
+ scanchain_72/module_data_out[5] scanchain_72/module_data_out[6] scanchain_72/module_data_out[7]
+ scanchain_72/scan_select_in scanchain_73/scan_select_in vccd1 vssd1 scanchain
Xscanchain_61 scanchain_61/clk_in scanchain_62/clk_in scanchain_61/data_in scanchain_62/data_in
+ scanchain_61/latch_enable_in scanchain_62/latch_enable_in scanchain_61/module_data_in[0]
+ scanchain_61/module_data_in[1] scanchain_61/module_data_in[2] scanchain_61/module_data_in[3]
+ scanchain_61/module_data_in[4] scanchain_61/module_data_in[5] scanchain_61/module_data_in[6]
+ scanchain_61/module_data_in[7] scanchain_61/module_data_out[0] scanchain_61/module_data_out[1]
+ scanchain_61/module_data_out[2] scanchain_61/module_data_out[3] scanchain_61/module_data_out[4]
+ scanchain_61/module_data_out[5] scanchain_61/module_data_out[6] scanchain_61/module_data_out[7]
+ scanchain_61/scan_select_in scanchain_62/scan_select_in vccd1 vssd1 scanchain
Xscanchain_83 scanchain_83/clk_in scanchain_84/clk_in scanchain_83/data_in scanchain_84/data_in
+ scanchain_83/latch_enable_in scanchain_84/latch_enable_in scanchain_83/module_data_in[0]
+ scanchain_83/module_data_in[1] scanchain_83/module_data_in[2] scanchain_83/module_data_in[3]
+ scanchain_83/module_data_in[4] scanchain_83/module_data_in[5] scanchain_83/module_data_in[6]
+ scanchain_83/module_data_in[7] scanchain_83/module_data_out[0] scanchain_83/module_data_out[1]
+ scanchain_83/module_data_out[2] scanchain_83/module_data_out[3] scanchain_83/module_data_out[4]
+ scanchain_83/module_data_out[5] scanchain_83/module_data_out[6] scanchain_83/module_data_out[7]
+ scanchain_83/scan_select_in scanchain_84/scan_select_in vccd1 vssd1 scanchain
Xscanchain_94 scanchain_94/clk_in scanchain_95/clk_in scanchain_94/data_in scanchain_95/data_in
+ scanchain_94/latch_enable_in scanchain_95/latch_enable_in scanchain_94/module_data_in[0]
+ scanchain_94/module_data_in[1] scanchain_94/module_data_in[2] scanchain_94/module_data_in[3]
+ scanchain_94/module_data_in[4] scanchain_94/module_data_in[5] scanchain_94/module_data_in[6]
+ scanchain_94/module_data_in[7] scanchain_94/module_data_out[0] scanchain_94/module_data_out[1]
+ scanchain_94/module_data_out[2] scanchain_94/module_data_out[3] scanchain_94/module_data_out[4]
+ scanchain_94/module_data_out[5] scanchain_94/module_data_out[6] scanchain_94/module_data_out[7]
+ scanchain_94/scan_select_in scanchain_95/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_463 scanchain_463/module_data_in[0] scanchain_463/module_data_in[1]
+ scanchain_463/module_data_in[2] scanchain_463/module_data_in[3] scanchain_463/module_data_in[4]
+ scanchain_463/module_data_in[5] scanchain_463/module_data_in[6] scanchain_463/module_data_in[7]
+ scanchain_463/module_data_out[0] scanchain_463/module_data_out[1] scanchain_463/module_data_out[2]
+ scanchain_463/module_data_out[3] scanchain_463/module_data_out[4] scanchain_463/module_data_out[5]
+ scanchain_463/module_data_out[6] scanchain_463/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_441 scanchain_441/module_data_in[0] scanchain_441/module_data_in[1]
+ scanchain_441/module_data_in[2] scanchain_441/module_data_in[3] scanchain_441/module_data_in[4]
+ scanchain_441/module_data_in[5] scanchain_441/module_data_in[6] scanchain_441/module_data_in[7]
+ scanchain_441/module_data_out[0] scanchain_441/module_data_out[1] scanchain_441/module_data_out[2]
+ scanchain_441/module_data_out[3] scanchain_441/module_data_out[4] scanchain_441/module_data_out[5]
+ scanchain_441/module_data_out[6] scanchain_441/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_452 scanchain_452/module_data_in[0] scanchain_452/module_data_in[1]
+ scanchain_452/module_data_in[2] scanchain_452/module_data_in[3] scanchain_452/module_data_in[4]
+ scanchain_452/module_data_in[5] scanchain_452/module_data_in[6] scanchain_452/module_data_in[7]
+ scanchain_452/module_data_out[0] scanchain_452/module_data_out[1] scanchain_452/module_data_out[2]
+ scanchain_452/module_data_out[3] scanchain_452/module_data_out[4] scanchain_452/module_data_out[5]
+ scanchain_452/module_data_out[6] scanchain_452/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_430 scanchain_430/module_data_in[0] scanchain_430/module_data_in[1]
+ scanchain_430/module_data_in[2] scanchain_430/module_data_in[3] scanchain_430/module_data_in[4]
+ scanchain_430/module_data_in[5] scanchain_430/module_data_in[6] scanchain_430/module_data_in[7]
+ scanchain_430/module_data_out[0] scanchain_430/module_data_out[1] scanchain_430/module_data_out[2]
+ scanchain_430/module_data_out[3] scanchain_430/module_data_out[4] scanchain_430/module_data_out[5]
+ scanchain_430/module_data_out[6] scanchain_430/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_416 scanchain_416/clk_in scanchain_417/clk_in scanchain_416/data_in scanchain_417/data_in
+ scanchain_416/latch_enable_in scanchain_417/latch_enable_in scanchain_416/module_data_in[0]
+ scanchain_416/module_data_in[1] scanchain_416/module_data_in[2] scanchain_416/module_data_in[3]
+ scanchain_416/module_data_in[4] scanchain_416/module_data_in[5] scanchain_416/module_data_in[6]
+ scanchain_416/module_data_in[7] scanchain_416/module_data_out[0] scanchain_416/module_data_out[1]
+ scanchain_416/module_data_out[2] scanchain_416/module_data_out[3] scanchain_416/module_data_out[4]
+ scanchain_416/module_data_out[5] scanchain_416/module_data_out[6] scanchain_416/module_data_out[7]
+ scanchain_416/scan_select_in scanchain_417/scan_select_in vccd1 vssd1 scanchain
Xscanchain_405 scanchain_405/clk_in scanchain_406/clk_in scanchain_405/data_in scanchain_406/data_in
+ scanchain_405/latch_enable_in scanchain_406/latch_enable_in scanchain_405/module_data_in[0]
+ scanchain_405/module_data_in[1] scanchain_405/module_data_in[2] scanchain_405/module_data_in[3]
+ scanchain_405/module_data_in[4] scanchain_405/module_data_in[5] scanchain_405/module_data_in[6]
+ scanchain_405/module_data_in[7] scanchain_405/module_data_out[0] scanchain_405/module_data_out[1]
+ scanchain_405/module_data_out[2] scanchain_405/module_data_out[3] scanchain_405/module_data_out[4]
+ scanchain_405/module_data_out[5] scanchain_405/module_data_out[6] scanchain_405/module_data_out[7]
+ scanchain_405/scan_select_in scanchain_406/scan_select_in vccd1 vssd1 scanchain
Xscanchain_438 scanchain_438/clk_in scanchain_439/clk_in scanchain_438/data_in scanchain_439/data_in
+ scanchain_438/latch_enable_in scanchain_439/latch_enable_in scanchain_438/module_data_in[0]
+ scanchain_438/module_data_in[1] scanchain_438/module_data_in[2] scanchain_438/module_data_in[3]
+ scanchain_438/module_data_in[4] scanchain_438/module_data_in[5] scanchain_438/module_data_in[6]
+ scanchain_438/module_data_in[7] scanchain_438/module_data_out[0] scanchain_438/module_data_out[1]
+ scanchain_438/module_data_out[2] scanchain_438/module_data_out[3] scanchain_438/module_data_out[4]
+ scanchain_438/module_data_out[5] scanchain_438/module_data_out[6] scanchain_438/module_data_out[7]
+ scanchain_438/scan_select_in scanchain_439/scan_select_in vccd1 vssd1 scanchain
Xscanchain_449 scanchain_449/clk_in scanchain_450/clk_in scanchain_449/data_in scanchain_450/data_in
+ scanchain_449/latch_enable_in scanchain_450/latch_enable_in scanchain_449/module_data_in[0]
+ scanchain_449/module_data_in[1] scanchain_449/module_data_in[2] scanchain_449/module_data_in[3]
+ scanchain_449/module_data_in[4] scanchain_449/module_data_in[5] scanchain_449/module_data_in[6]
+ scanchain_449/module_data_in[7] scanchain_449/module_data_out[0] scanchain_449/module_data_out[1]
+ scanchain_449/module_data_out[2] scanchain_449/module_data_out[3] scanchain_449/module_data_out[4]
+ scanchain_449/module_data_out[5] scanchain_449/module_data_out[6] scanchain_449/module_data_out[7]
+ scanchain_449/scan_select_in scanchain_450/scan_select_in vccd1 vssd1 scanchain
Xscanchain_427 scanchain_427/clk_in scanchain_428/clk_in scanchain_427/data_in scanchain_428/data_in
+ scanchain_427/latch_enable_in scanchain_428/latch_enable_in scanchain_427/module_data_in[0]
+ scanchain_427/module_data_in[1] scanchain_427/module_data_in[2] scanchain_427/module_data_in[3]
+ scanchain_427/module_data_in[4] scanchain_427/module_data_in[5] scanchain_427/module_data_in[6]
+ scanchain_427/module_data_in[7] scanchain_427/module_data_out[0] scanchain_427/module_data_out[1]
+ scanchain_427/module_data_out[2] scanchain_427/module_data_out[3] scanchain_427/module_data_out[4]
+ scanchain_427/module_data_out[5] scanchain_427/module_data_out[6] scanchain_427/module_data_out[7]
+ scanchain_427/scan_select_in scanchain_428/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_293 scanchain_293/module_data_in[0] scanchain_293/module_data_in[1]
+ scanchain_293/module_data_in[2] scanchain_293/module_data_in[3] scanchain_293/module_data_in[4]
+ scanchain_293/module_data_in[5] scanchain_293/module_data_in[6] scanchain_293/module_data_in[7]
+ scanchain_293/module_data_out[0] scanchain_293/module_data_out[1] scanchain_293/module_data_out[2]
+ scanchain_293/module_data_out[3] scanchain_293/module_data_out[4] scanchain_293/module_data_out[5]
+ scanchain_293/module_data_out[6] scanchain_293/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_282 scanchain_282/module_data_in[0] scanchain_282/module_data_in[1]
+ scanchain_282/module_data_in[2] scanchain_282/module_data_in[3] scanchain_282/module_data_in[4]
+ scanchain_282/module_data_in[5] scanchain_282/module_data_in[6] scanchain_282/module_data_in[7]
+ scanchain_282/module_data_out[0] scanchain_282/module_data_out[1] scanchain_282/module_data_out[2]
+ scanchain_282/module_data_out[3] scanchain_282/module_data_out[4] scanchain_282/module_data_out[5]
+ scanchain_282/module_data_out[6] scanchain_282/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_279 scanchain_279/clk_in scanchain_280/clk_in scanchain_279/data_in scanchain_280/data_in
+ scanchain_279/latch_enable_in scanchain_280/latch_enable_in scanchain_279/module_data_in[0]
+ scanchain_279/module_data_in[1] scanchain_279/module_data_in[2] scanchain_279/module_data_in[3]
+ scanchain_279/module_data_in[4] scanchain_279/module_data_in[5] scanchain_279/module_data_in[6]
+ scanchain_279/module_data_in[7] scanchain_279/module_data_out[0] scanchain_279/module_data_out[1]
+ scanchain_279/module_data_out[2] scanchain_279/module_data_out[3] scanchain_279/module_data_out[4]
+ scanchain_279/module_data_out[5] scanchain_279/module_data_out[6] scanchain_279/module_data_out[7]
+ scanchain_279/scan_select_in scanchain_280/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_271 scanchain_271/module_data_in[0] scanchain_271/module_data_in[1]
+ scanchain_271/module_data_in[2] scanchain_271/module_data_in[3] scanchain_271/module_data_in[4]
+ scanchain_271/module_data_in[5] scanchain_271/module_data_in[6] scanchain_271/module_data_in[7]
+ scanchain_271/module_data_out[0] scanchain_271/module_data_out[1] scanchain_271/module_data_out[2]
+ scanchain_271/module_data_out[3] scanchain_271/module_data_out[4] scanchain_271/module_data_out[5]
+ scanchain_271/module_data_out[6] scanchain_271/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_268 scanchain_268/clk_in scanchain_269/clk_in scanchain_268/data_in scanchain_269/data_in
+ scanchain_268/latch_enable_in scanchain_269/latch_enable_in scanchain_268/module_data_in[0]
+ scanchain_268/module_data_in[1] scanchain_268/module_data_in[2] scanchain_268/module_data_in[3]
+ scanchain_268/module_data_in[4] scanchain_268/module_data_in[5] scanchain_268/module_data_in[6]
+ scanchain_268/module_data_in[7] scanchain_268/module_data_out[0] scanchain_268/module_data_out[1]
+ scanchain_268/module_data_out[2] scanchain_268/module_data_out[3] scanchain_268/module_data_out[4]
+ scanchain_268/module_data_out[5] scanchain_268/module_data_out[6] scanchain_268/module_data_out[7]
+ scanchain_268/scan_select_in scanchain_269/scan_select_in vccd1 vssd1 scanchain
Xscanchain_246 scanchain_246/clk_in scanchain_247/clk_in scanchain_246/data_in scanchain_247/data_in
+ scanchain_246/latch_enable_in scanchain_247/latch_enable_in scanchain_246/module_data_in[0]
+ scanchain_246/module_data_in[1] scanchain_246/module_data_in[2] scanchain_246/module_data_in[3]
+ scanchain_246/module_data_in[4] scanchain_246/module_data_in[5] scanchain_246/module_data_in[6]
+ scanchain_246/module_data_in[7] scanchain_246/module_data_out[0] scanchain_246/module_data_out[1]
+ scanchain_246/module_data_out[2] scanchain_246/module_data_out[3] scanchain_246/module_data_out[4]
+ scanchain_246/module_data_out[5] scanchain_246/module_data_out[6] scanchain_246/module_data_out[7]
+ scanchain_246/scan_select_in scanchain_247/scan_select_in vccd1 vssd1 scanchain
Xscanchain_257 scanchain_257/clk_in scanchain_258/clk_in scanchain_257/data_in scanchain_258/data_in
+ scanchain_257/latch_enable_in scanchain_258/latch_enable_in scanchain_257/module_data_in[0]
+ scanchain_257/module_data_in[1] scanchain_257/module_data_in[2] scanchain_257/module_data_in[3]
+ scanchain_257/module_data_in[4] scanchain_257/module_data_in[5] scanchain_257/module_data_in[6]
+ scanchain_257/module_data_in[7] scanchain_257/module_data_out[0] scanchain_257/module_data_out[1]
+ scanchain_257/module_data_out[2] scanchain_257/module_data_out[3] scanchain_257/module_data_out[4]
+ scanchain_257/module_data_out[5] scanchain_257/module_data_out[6] scanchain_257/module_data_out[7]
+ scanchain_257/scan_select_in scanchain_258/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_260 scanchain_260/module_data_in[0] scanchain_260/module_data_in[1]
+ scanchain_260/module_data_in[2] scanchain_260/module_data_in[3] scanchain_260/module_data_in[4]
+ scanchain_260/module_data_in[5] scanchain_260/module_data_in[6] scanchain_260/module_data_in[7]
+ scanchain_260/module_data_out[0] scanchain_260/module_data_out[1] scanchain_260/module_data_out[2]
+ scanchain_260/module_data_out[3] scanchain_260/module_data_out[4] scanchain_260/module_data_out[5]
+ scanchain_260/module_data_out[6] scanchain_260/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_235 scanchain_235/clk_in scanchain_236/clk_in scanchain_235/data_in scanchain_236/data_in
+ scanchain_235/latch_enable_in scanchain_236/latch_enable_in scanchain_235/module_data_in[0]
+ scanchain_235/module_data_in[1] scanchain_235/module_data_in[2] scanchain_235/module_data_in[3]
+ scanchain_235/module_data_in[4] scanchain_235/module_data_in[5] scanchain_235/module_data_in[6]
+ scanchain_235/module_data_in[7] scanchain_235/module_data_out[0] scanchain_235/module_data_out[1]
+ scanchain_235/module_data_out[2] scanchain_235/module_data_out[3] scanchain_235/module_data_out[4]
+ scanchain_235/module_data_out[5] scanchain_235/module_data_out[6] scanchain_235/module_data_out[7]
+ scanchain_235/scan_select_in scanchain_236/scan_select_in vccd1 vssd1 scanchain
Xscanchain_213 scanchain_213/clk_in scanchain_214/clk_in scanchain_213/data_in scanchain_214/data_in
+ scanchain_213/latch_enable_in scanchain_214/latch_enable_in scanchain_213/module_data_in[0]
+ scanchain_213/module_data_in[1] scanchain_213/module_data_in[2] scanchain_213/module_data_in[3]
+ scanchain_213/module_data_in[4] scanchain_213/module_data_in[5] scanchain_213/module_data_in[6]
+ scanchain_213/module_data_in[7] scanchain_213/module_data_out[0] scanchain_213/module_data_out[1]
+ scanchain_213/module_data_out[2] scanchain_213/module_data_out[3] scanchain_213/module_data_out[4]
+ scanchain_213/module_data_out[5] scanchain_213/module_data_out[6] scanchain_213/module_data_out[7]
+ scanchain_213/scan_select_in scanchain_214/scan_select_in vccd1 vssd1 scanchain
Xscanchain_224 scanchain_224/clk_in scanchain_225/clk_in scanchain_224/data_in scanchain_225/data_in
+ scanchain_224/latch_enable_in scanchain_225/latch_enable_in scanchain_224/module_data_in[0]
+ scanchain_224/module_data_in[1] scanchain_224/module_data_in[2] scanchain_224/module_data_in[3]
+ scanchain_224/module_data_in[4] scanchain_224/module_data_in[5] scanchain_224/module_data_in[6]
+ scanchain_224/module_data_in[7] scanchain_224/module_data_out[0] scanchain_224/module_data_out[1]
+ scanchain_224/module_data_out[2] scanchain_224/module_data_out[3] scanchain_224/module_data_out[4]
+ scanchain_224/module_data_out[5] scanchain_224/module_data_out[6] scanchain_224/module_data_out[7]
+ scanchain_224/scan_select_in scanchain_225/scan_select_in vccd1 vssd1 scanchain
Xscanchain_202 scanchain_202/clk_in scanchain_203/clk_in scanchain_202/data_in scanchain_203/data_in
+ scanchain_202/latch_enable_in scanchain_203/latch_enable_in scanchain_202/module_data_in[0]
+ scanchain_202/module_data_in[1] scanchain_202/module_data_in[2] scanchain_202/module_data_in[3]
+ scanchain_202/module_data_in[4] scanchain_202/module_data_in[5] scanchain_202/module_data_in[6]
+ scanchain_202/module_data_in[7] scanchain_202/module_data_out[0] scanchain_202/module_data_out[1]
+ scanchain_202/module_data_out[2] scanchain_202/module_data_out[3] scanchain_202/module_data_out[4]
+ scanchain_202/module_data_out[5] scanchain_202/module_data_out[6] scanchain_202/module_data_out[7]
+ scanchain_202/scan_select_in scanchain_203/scan_select_in vccd1 vssd1 scanchain
Xscanchain_40 scanchain_40/clk_in scanchain_41/clk_in scanchain_40/data_in scanchain_41/data_in
+ scanchain_40/latch_enable_in scanchain_41/latch_enable_in yupferris_bitslam_40/io_in[0]
+ yupferris_bitslam_40/io_in[1] yupferris_bitslam_40/io_in[2] yupferris_bitslam_40/io_in[3]
+ yupferris_bitslam_40/io_in[4] yupferris_bitslam_40/io_in[5] yupferris_bitslam_40/io_in[6]
+ yupferris_bitslam_40/io_in[7] yupferris_bitslam_40/io_out[0] yupferris_bitslam_40/io_out[1]
+ yupferris_bitslam_40/io_out[2] yupferris_bitslam_40/io_out[3] yupferris_bitslam_40/io_out[4]
+ yupferris_bitslam_40/io_out[5] yupferris_bitslam_40/io_out[6] yupferris_bitslam_40/io_out[7]
+ scanchain_40/scan_select_in scanchain_41/scan_select_in vccd1 vssd1 scanchain
Xscanchain_51 scanchain_51/clk_in scanchain_52/clk_in scanchain_51/data_in scanchain_52/data_in
+ scanchain_51/latch_enable_in scanchain_52/latch_enable_in scanchain_51/module_data_in[0]
+ scanchain_51/module_data_in[1] scanchain_51/module_data_in[2] scanchain_51/module_data_in[3]
+ scanchain_51/module_data_in[4] scanchain_51/module_data_in[5] scanchain_51/module_data_in[6]
+ scanchain_51/module_data_in[7] scanchain_51/module_data_out[0] scanchain_51/module_data_out[1]
+ scanchain_51/module_data_out[2] scanchain_51/module_data_out[3] scanchain_51/module_data_out[4]
+ scanchain_51/module_data_out[5] scanchain_51/module_data_out[6] scanchain_51/module_data_out[7]
+ scanchain_51/scan_select_in scanchain_52/scan_select_in vccd1 vssd1 scanchain
Xscanchain_73 scanchain_73/clk_in scanchain_74/clk_in scanchain_73/data_in scanchain_74/data_in
+ scanchain_73/latch_enable_in scanchain_74/latch_enable_in scanchain_73/module_data_in[0]
+ scanchain_73/module_data_in[1] scanchain_73/module_data_in[2] scanchain_73/module_data_in[3]
+ scanchain_73/module_data_in[4] scanchain_73/module_data_in[5] scanchain_73/module_data_in[6]
+ scanchain_73/module_data_in[7] scanchain_73/module_data_out[0] scanchain_73/module_data_out[1]
+ scanchain_73/module_data_out[2] scanchain_73/module_data_out[3] scanchain_73/module_data_out[4]
+ scanchain_73/module_data_out[5] scanchain_73/module_data_out[6] scanchain_73/module_data_out[7]
+ scanchain_73/scan_select_in scanchain_74/scan_select_in vccd1 vssd1 scanchain
Xscanchain_62 scanchain_62/clk_in scanchain_63/clk_in scanchain_62/data_in scanchain_63/data_in
+ scanchain_62/latch_enable_in scanchain_63/latch_enable_in scanchain_62/module_data_in[0]
+ scanchain_62/module_data_in[1] scanchain_62/module_data_in[2] scanchain_62/module_data_in[3]
+ scanchain_62/module_data_in[4] scanchain_62/module_data_in[5] scanchain_62/module_data_in[6]
+ scanchain_62/module_data_in[7] scanchain_62/module_data_out[0] scanchain_62/module_data_out[1]
+ scanchain_62/module_data_out[2] scanchain_62/module_data_out[3] scanchain_62/module_data_out[4]
+ scanchain_62/module_data_out[5] scanchain_62/module_data_out[6] scanchain_62/module_data_out[7]
+ scanchain_62/scan_select_in scanchain_63/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_80 scanchain_80/module_data_in[0] scanchain_80/module_data_in[1]
+ scanchain_80/module_data_in[2] scanchain_80/module_data_in[3] scanchain_80/module_data_in[4]
+ scanchain_80/module_data_in[5] scanchain_80/module_data_in[6] scanchain_80/module_data_in[7]
+ scanchain_80/module_data_out[0] scanchain_80/module_data_out[1] scanchain_80/module_data_out[2]
+ scanchain_80/module_data_out[3] scanchain_80/module_data_out[4] scanchain_80/module_data_out[5]
+ scanchain_80/module_data_out[6] scanchain_80/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_84 scanchain_84/clk_in scanchain_85/clk_in scanchain_84/data_in scanchain_85/data_in
+ scanchain_84/latch_enable_in scanchain_85/latch_enable_in scanchain_84/module_data_in[0]
+ scanchain_84/module_data_in[1] scanchain_84/module_data_in[2] scanchain_84/module_data_in[3]
+ scanchain_84/module_data_in[4] scanchain_84/module_data_in[5] scanchain_84/module_data_in[6]
+ scanchain_84/module_data_in[7] scanchain_84/module_data_out[0] scanchain_84/module_data_out[1]
+ scanchain_84/module_data_out[2] scanchain_84/module_data_out[3] scanchain_84/module_data_out[4]
+ scanchain_84/module_data_out[5] scanchain_84/module_data_out[6] scanchain_84/module_data_out[7]
+ scanchain_84/scan_select_in scanchain_85/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_91 scanchain_91/module_data_in[0] scanchain_91/module_data_in[1]
+ scanchain_91/module_data_in[2] scanchain_91/module_data_in[3] scanchain_91/module_data_in[4]
+ scanchain_91/module_data_in[5] scanchain_91/module_data_in[6] scanchain_91/module_data_in[7]
+ scanchain_91/module_data_out[0] scanchain_91/module_data_out[1] scanchain_91/module_data_out[2]
+ scanchain_91/module_data_out[3] scanchain_91/module_data_out[4] scanchain_91/module_data_out[5]
+ scanchain_91/module_data_out[6] scanchain_91/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_95 scanchain_95/clk_in scanchain_96/clk_in scanchain_95/data_in scanchain_96/data_in
+ scanchain_95/latch_enable_in scanchain_96/latch_enable_in scanchain_95/module_data_in[0]
+ scanchain_95/module_data_in[1] scanchain_95/module_data_in[2] scanchain_95/module_data_in[3]
+ scanchain_95/module_data_in[4] scanchain_95/module_data_in[5] scanchain_95/module_data_in[6]
+ scanchain_95/module_data_in[7] scanchain_95/module_data_out[0] scanchain_95/module_data_out[1]
+ scanchain_95/module_data_out[2] scanchain_95/module_data_out[3] scanchain_95/module_data_out[4]
+ scanchain_95/module_data_out[5] scanchain_95/module_data_out[6] scanchain_95/module_data_out[7]
+ scanchain_95/scan_select_in scanchain_96/scan_select_in vccd1 vssd1 scanchain
Xjar_illegal_logic_36 jar_illegal_logic_36/io_in[0] jar_illegal_logic_36/io_in[1]
+ jar_illegal_logic_36/io_in[2] jar_illegal_logic_36/io_in[3] jar_illegal_logic_36/io_in[4]
+ jar_illegal_logic_36/io_in[5] jar_illegal_logic_36/io_in[6] jar_illegal_logic_36/io_in[7]
+ jar_illegal_logic_36/io_out[0] jar_illegal_logic_36/io_out[1] jar_illegal_logic_36/io_out[2]
+ jar_illegal_logic_36/io_out[3] jar_illegal_logic_36/io_out[4] jar_illegal_logic_36/io_out[5]
+ jar_illegal_logic_36/io_out[6] jar_illegal_logic_36/io_out[7] vccd1 vssd1 jar_illegal_logic
Xaidan_McCoy_8 aidan_McCoy_8/io_in[0] aidan_McCoy_8/io_in[1] aidan_McCoy_8/io_in[2]
+ aidan_McCoy_8/io_in[3] aidan_McCoy_8/io_in[4] aidan_McCoy_8/io_in[5] aidan_McCoy_8/io_in[6]
+ aidan_McCoy_8/io_in[7] aidan_McCoy_8/io_out[0] aidan_McCoy_8/io_out[1] aidan_McCoy_8/io_out[2]
+ aidan_McCoy_8/io_out[3] aidan_McCoy_8/io_out[4] aidan_McCoy_8/io_out[5] aidan_McCoy_8/io_out[6]
+ aidan_McCoy_8/io_out[7] vccd1 vssd1 aidan_McCoy
Xuser_module_339501025136214612_464 scanchain_464/module_data_in[0] scanchain_464/module_data_in[1]
+ scanchain_464/module_data_in[2] scanchain_464/module_data_in[3] scanchain_464/module_data_in[4]
+ scanchain_464/module_data_in[5] scanchain_464/module_data_in[6] scanchain_464/module_data_in[7]
+ scanchain_464/module_data_out[0] scanchain_464/module_data_out[1] scanchain_464/module_data_out[2]
+ scanchain_464/module_data_out[3] scanchain_464/module_data_out[4] scanchain_464/module_data_out[5]
+ scanchain_464/module_data_out[6] scanchain_464/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_442 scanchain_442/module_data_in[0] scanchain_442/module_data_in[1]
+ scanchain_442/module_data_in[2] scanchain_442/module_data_in[3] scanchain_442/module_data_in[4]
+ scanchain_442/module_data_in[5] scanchain_442/module_data_in[6] scanchain_442/module_data_in[7]
+ scanchain_442/module_data_out[0] scanchain_442/module_data_out[1] scanchain_442/module_data_out[2]
+ scanchain_442/module_data_out[3] scanchain_442/module_data_out[4] scanchain_442/module_data_out[5]
+ scanchain_442/module_data_out[6] scanchain_442/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_453 scanchain_453/module_data_in[0] scanchain_453/module_data_in[1]
+ scanchain_453/module_data_in[2] scanchain_453/module_data_in[3] scanchain_453/module_data_in[4]
+ scanchain_453/module_data_in[5] scanchain_453/module_data_in[6] scanchain_453/module_data_in[7]
+ scanchain_453/module_data_out[0] scanchain_453/module_data_out[1] scanchain_453/module_data_out[2]
+ scanchain_453/module_data_out[3] scanchain_453/module_data_out[4] scanchain_453/module_data_out[5]
+ scanchain_453/module_data_out[6] scanchain_453/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_431 scanchain_431/module_data_in[0] scanchain_431/module_data_in[1]
+ scanchain_431/module_data_in[2] scanchain_431/module_data_in[3] scanchain_431/module_data_in[4]
+ scanchain_431/module_data_in[5] scanchain_431/module_data_in[6] scanchain_431/module_data_in[7]
+ scanchain_431/module_data_out[0] scanchain_431/module_data_out[1] scanchain_431/module_data_out[2]
+ scanchain_431/module_data_out[3] scanchain_431/module_data_out[4] scanchain_431/module_data_out[5]
+ scanchain_431/module_data_out[6] scanchain_431/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_420 scanchain_420/module_data_in[0] scanchain_420/module_data_in[1]
+ scanchain_420/module_data_in[2] scanchain_420/module_data_in[3] scanchain_420/module_data_in[4]
+ scanchain_420/module_data_in[5] scanchain_420/module_data_in[6] scanchain_420/module_data_in[7]
+ scanchain_420/module_data_out[0] scanchain_420/module_data_out[1] scanchain_420/module_data_out[2]
+ scanchain_420/module_data_out[3] scanchain_420/module_data_out[4] scanchain_420/module_data_out[5]
+ scanchain_420/module_data_out[6] scanchain_420/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_439 scanchain_439/clk_in scanchain_440/clk_in scanchain_439/data_in scanchain_440/data_in
+ scanchain_439/latch_enable_in scanchain_440/latch_enable_in scanchain_439/module_data_in[0]
+ scanchain_439/module_data_in[1] scanchain_439/module_data_in[2] scanchain_439/module_data_in[3]
+ scanchain_439/module_data_in[4] scanchain_439/module_data_in[5] scanchain_439/module_data_in[6]
+ scanchain_439/module_data_in[7] scanchain_439/module_data_out[0] scanchain_439/module_data_out[1]
+ scanchain_439/module_data_out[2] scanchain_439/module_data_out[3] scanchain_439/module_data_out[4]
+ scanchain_439/module_data_out[5] scanchain_439/module_data_out[6] scanchain_439/module_data_out[7]
+ scanchain_439/scan_select_in scanchain_440/scan_select_in vccd1 vssd1 scanchain
Xscanchain_428 scanchain_428/clk_in scanchain_429/clk_in scanchain_428/data_in scanchain_429/data_in
+ scanchain_428/latch_enable_in scanchain_429/latch_enable_in scanchain_428/module_data_in[0]
+ scanchain_428/module_data_in[1] scanchain_428/module_data_in[2] scanchain_428/module_data_in[3]
+ scanchain_428/module_data_in[4] scanchain_428/module_data_in[5] scanchain_428/module_data_in[6]
+ scanchain_428/module_data_in[7] scanchain_428/module_data_out[0] scanchain_428/module_data_out[1]
+ scanchain_428/module_data_out[2] scanchain_428/module_data_out[3] scanchain_428/module_data_out[4]
+ scanchain_428/module_data_out[5] scanchain_428/module_data_out[6] scanchain_428/module_data_out[7]
+ scanchain_428/scan_select_in scanchain_429/scan_select_in vccd1 vssd1 scanchain
Xscanchain_417 scanchain_417/clk_in scanchain_418/clk_in scanchain_417/data_in scanchain_418/data_in
+ scanchain_417/latch_enable_in scanchain_418/latch_enable_in scanchain_417/module_data_in[0]
+ scanchain_417/module_data_in[1] scanchain_417/module_data_in[2] scanchain_417/module_data_in[3]
+ scanchain_417/module_data_in[4] scanchain_417/module_data_in[5] scanchain_417/module_data_in[6]
+ scanchain_417/module_data_in[7] scanchain_417/module_data_out[0] scanchain_417/module_data_out[1]
+ scanchain_417/module_data_out[2] scanchain_417/module_data_out[3] scanchain_417/module_data_out[4]
+ scanchain_417/module_data_out[5] scanchain_417/module_data_out[6] scanchain_417/module_data_out[7]
+ scanchain_417/scan_select_in scanchain_418/scan_select_in vccd1 vssd1 scanchain
Xscanchain_406 scanchain_406/clk_in scanchain_407/clk_in scanchain_406/data_in scanchain_407/data_in
+ scanchain_406/latch_enable_in scanchain_407/latch_enable_in scanchain_406/module_data_in[0]
+ scanchain_406/module_data_in[1] scanchain_406/module_data_in[2] scanchain_406/module_data_in[3]
+ scanchain_406/module_data_in[4] scanchain_406/module_data_in[5] scanchain_406/module_data_in[6]
+ scanchain_406/module_data_in[7] scanchain_406/module_data_out[0] scanchain_406/module_data_out[1]
+ scanchain_406/module_data_out[2] scanchain_406/module_data_out[3] scanchain_406/module_data_out[4]
+ scanchain_406/module_data_out[5] scanchain_406/module_data_out[6] scanchain_406/module_data_out[7]
+ scanchain_406/scan_select_in scanchain_407/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_283 scanchain_283/module_data_in[0] scanchain_283/module_data_in[1]
+ scanchain_283/module_data_in[2] scanchain_283/module_data_in[3] scanchain_283/module_data_in[4]
+ scanchain_283/module_data_in[5] scanchain_283/module_data_in[6] scanchain_283/module_data_in[7]
+ scanchain_283/module_data_out[0] scanchain_283/module_data_out[1] scanchain_283/module_data_out[2]
+ scanchain_283/module_data_out[3] scanchain_283/module_data_out[4] scanchain_283/module_data_out[5]
+ scanchain_283/module_data_out[6] scanchain_283/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_294 scanchain_294/module_data_in[0] scanchain_294/module_data_in[1]
+ scanchain_294/module_data_in[2] scanchain_294/module_data_in[3] scanchain_294/module_data_in[4]
+ scanchain_294/module_data_in[5] scanchain_294/module_data_in[6] scanchain_294/module_data_in[7]
+ scanchain_294/module_data_out[0] scanchain_294/module_data_out[1] scanchain_294/module_data_out[2]
+ scanchain_294/module_data_out[3] scanchain_294/module_data_out[4] scanchain_294/module_data_out[5]
+ scanchain_294/module_data_out[6] scanchain_294/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_272 scanchain_272/module_data_in[0] scanchain_272/module_data_in[1]
+ scanchain_272/module_data_in[2] scanchain_272/module_data_in[3] scanchain_272/module_data_in[4]
+ scanchain_272/module_data_in[5] scanchain_272/module_data_in[6] scanchain_272/module_data_in[7]
+ scanchain_272/module_data_out[0] scanchain_272/module_data_out[1] scanchain_272/module_data_out[2]
+ scanchain_272/module_data_out[3] scanchain_272/module_data_out[4] scanchain_272/module_data_out[5]
+ scanchain_272/module_data_out[6] scanchain_272/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_269 scanchain_269/clk_in scanchain_270/clk_in scanchain_269/data_in scanchain_270/data_in
+ scanchain_269/latch_enable_in scanchain_270/latch_enable_in scanchain_269/module_data_in[0]
+ scanchain_269/module_data_in[1] scanchain_269/module_data_in[2] scanchain_269/module_data_in[3]
+ scanchain_269/module_data_in[4] scanchain_269/module_data_in[5] scanchain_269/module_data_in[6]
+ scanchain_269/module_data_in[7] scanchain_269/module_data_out[0] scanchain_269/module_data_out[1]
+ scanchain_269/module_data_out[2] scanchain_269/module_data_out[3] scanchain_269/module_data_out[4]
+ scanchain_269/module_data_out[5] scanchain_269/module_data_out[6] scanchain_269/module_data_out[7]
+ scanchain_269/scan_select_in scanchain_270/scan_select_in vccd1 vssd1 scanchain
Xscanchain_247 scanchain_247/clk_in scanchain_248/clk_in scanchain_247/data_in scanchain_248/data_in
+ scanchain_247/latch_enable_in scanchain_248/latch_enable_in scanchain_247/module_data_in[0]
+ scanchain_247/module_data_in[1] scanchain_247/module_data_in[2] scanchain_247/module_data_in[3]
+ scanchain_247/module_data_in[4] scanchain_247/module_data_in[5] scanchain_247/module_data_in[6]
+ scanchain_247/module_data_in[7] scanchain_247/module_data_out[0] scanchain_247/module_data_out[1]
+ scanchain_247/module_data_out[2] scanchain_247/module_data_out[3] scanchain_247/module_data_out[4]
+ scanchain_247/module_data_out[5] scanchain_247/module_data_out[6] scanchain_247/module_data_out[7]
+ scanchain_247/scan_select_in scanchain_248/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_250 scanchain_250/module_data_in[0] scanchain_250/module_data_in[1]
+ scanchain_250/module_data_in[2] scanchain_250/module_data_in[3] scanchain_250/module_data_in[4]
+ scanchain_250/module_data_in[5] scanchain_250/module_data_in[6] scanchain_250/module_data_in[7]
+ scanchain_250/module_data_out[0] scanchain_250/module_data_out[1] scanchain_250/module_data_out[2]
+ scanchain_250/module_data_out[3] scanchain_250/module_data_out[4] scanchain_250/module_data_out[5]
+ scanchain_250/module_data_out[6] scanchain_250/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_258 scanchain_258/clk_in scanchain_259/clk_in scanchain_258/data_in scanchain_259/data_in
+ scanchain_258/latch_enable_in scanchain_259/latch_enable_in scanchain_258/module_data_in[0]
+ scanchain_258/module_data_in[1] scanchain_258/module_data_in[2] scanchain_258/module_data_in[3]
+ scanchain_258/module_data_in[4] scanchain_258/module_data_in[5] scanchain_258/module_data_in[6]
+ scanchain_258/module_data_in[7] scanchain_258/module_data_out[0] scanchain_258/module_data_out[1]
+ scanchain_258/module_data_out[2] scanchain_258/module_data_out[3] scanchain_258/module_data_out[4]
+ scanchain_258/module_data_out[5] scanchain_258/module_data_out[6] scanchain_258/module_data_out[7]
+ scanchain_258/scan_select_in scanchain_259/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_261 scanchain_261/module_data_in[0] scanchain_261/module_data_in[1]
+ scanchain_261/module_data_in[2] scanchain_261/module_data_in[3] scanchain_261/module_data_in[4]
+ scanchain_261/module_data_in[5] scanchain_261/module_data_in[6] scanchain_261/module_data_in[7]
+ scanchain_261/module_data_out[0] scanchain_261/module_data_out[1] scanchain_261/module_data_out[2]
+ scanchain_261/module_data_out[3] scanchain_261/module_data_out[4] scanchain_261/module_data_out[5]
+ scanchain_261/module_data_out[6] scanchain_261/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_236 scanchain_236/clk_in scanchain_237/clk_in scanchain_236/data_in scanchain_237/data_in
+ scanchain_236/latch_enable_in scanchain_237/latch_enable_in scanchain_236/module_data_in[0]
+ scanchain_236/module_data_in[1] scanchain_236/module_data_in[2] scanchain_236/module_data_in[3]
+ scanchain_236/module_data_in[4] scanchain_236/module_data_in[5] scanchain_236/module_data_in[6]
+ scanchain_236/module_data_in[7] scanchain_236/module_data_out[0] scanchain_236/module_data_out[1]
+ scanchain_236/module_data_out[2] scanchain_236/module_data_out[3] scanchain_236/module_data_out[4]
+ scanchain_236/module_data_out[5] scanchain_236/module_data_out[6] scanchain_236/module_data_out[7]
+ scanchain_236/scan_select_in scanchain_237/scan_select_in vccd1 vssd1 scanchain
Xscanchain_214 scanchain_214/clk_in scanchain_215/clk_in scanchain_214/data_in scanchain_215/data_in
+ scanchain_214/latch_enable_in scanchain_215/latch_enable_in scanchain_214/module_data_in[0]
+ scanchain_214/module_data_in[1] scanchain_214/module_data_in[2] scanchain_214/module_data_in[3]
+ scanchain_214/module_data_in[4] scanchain_214/module_data_in[5] scanchain_214/module_data_in[6]
+ scanchain_214/module_data_in[7] scanchain_214/module_data_out[0] scanchain_214/module_data_out[1]
+ scanchain_214/module_data_out[2] scanchain_214/module_data_out[3] scanchain_214/module_data_out[4]
+ scanchain_214/module_data_out[5] scanchain_214/module_data_out[6] scanchain_214/module_data_out[7]
+ scanchain_214/scan_select_in scanchain_215/scan_select_in vccd1 vssd1 scanchain
Xscanchain_225 scanchain_225/clk_in scanchain_226/clk_in scanchain_225/data_in scanchain_226/data_in
+ scanchain_225/latch_enable_in scanchain_226/latch_enable_in scanchain_225/module_data_in[0]
+ scanchain_225/module_data_in[1] scanchain_225/module_data_in[2] scanchain_225/module_data_in[3]
+ scanchain_225/module_data_in[4] scanchain_225/module_data_in[5] scanchain_225/module_data_in[6]
+ scanchain_225/module_data_in[7] scanchain_225/module_data_out[0] scanchain_225/module_data_out[1]
+ scanchain_225/module_data_out[2] scanchain_225/module_data_out[3] scanchain_225/module_data_out[4]
+ scanchain_225/module_data_out[5] scanchain_225/module_data_out[6] scanchain_225/module_data_out[7]
+ scanchain_225/scan_select_in scanchain_226/scan_select_in vccd1 vssd1 scanchain
Xscanchain_203 scanchain_203/clk_in scanchain_204/clk_in scanchain_203/data_in scanchain_204/data_in
+ scanchain_203/latch_enable_in scanchain_204/latch_enable_in scanchain_203/module_data_in[0]
+ scanchain_203/module_data_in[1] scanchain_203/module_data_in[2] scanchain_203/module_data_in[3]
+ scanchain_203/module_data_in[4] scanchain_203/module_data_in[5] scanchain_203/module_data_in[6]
+ scanchain_203/module_data_in[7] scanchain_203/module_data_out[0] scanchain_203/module_data_out[1]
+ scanchain_203/module_data_out[2] scanchain_203/module_data_out[3] scanchain_203/module_data_out[4]
+ scanchain_203/module_data_out[5] scanchain_203/module_data_out[6] scanchain_203/module_data_out[7]
+ scanchain_203/scan_select_in scanchain_204/scan_select_in vccd1 vssd1 scanchain
Xscanchain_41 scanchain_41/clk_in scanchain_42/clk_in scanchain_41/data_in scanchain_42/data_in
+ scanchain_41/latch_enable_in scanchain_42/latch_enable_in scanchain_41/module_data_in[0]
+ scanchain_41/module_data_in[1] scanchain_41/module_data_in[2] scanchain_41/module_data_in[3]
+ scanchain_41/module_data_in[4] scanchain_41/module_data_in[5] scanchain_41/module_data_in[6]
+ scanchain_41/module_data_in[7] scanchain_41/module_data_out[0] scanchain_41/module_data_out[1]
+ scanchain_41/module_data_out[2] scanchain_41/module_data_out[3] scanchain_41/module_data_out[4]
+ scanchain_41/module_data_out[5] scanchain_41/module_data_out[6] scanchain_41/module_data_out[7]
+ scanchain_41/scan_select_in scanchain_42/scan_select_in vccd1 vssd1 scanchain
Xscanchain_30 scanchain_30/clk_in scanchain_31/clk_in scanchain_30/data_in scanchain_31/data_in
+ scanchain_30/latch_enable_in scanchain_31/latch_enable_in scanchain_30/module_data_in[0]
+ scanchain_30/module_data_in[1] scanchain_30/module_data_in[2] scanchain_30/module_data_in[3]
+ scanchain_30/module_data_in[4] scanchain_30/module_data_in[5] scanchain_30/module_data_in[6]
+ scanchain_30/module_data_in[7] scanchain_30/module_data_out[0] scanchain_30/module_data_out[1]
+ scanchain_30/module_data_out[2] scanchain_30/module_data_out[3] scanchain_30/module_data_out[4]
+ scanchain_30/module_data_out[5] scanchain_30/module_data_out[6] scanchain_30/module_data_out[7]
+ scanchain_30/scan_select_in scanchain_31/scan_select_in vccd1 vssd1 scanchain
Xscanchain_52 scanchain_52/clk_in scanchain_53/clk_in scanchain_52/data_in scanchain_53/data_in
+ scanchain_52/latch_enable_in scanchain_53/latch_enable_in xor_shift32_evango_52/io_in[0]
+ xor_shift32_evango_52/io_in[1] xor_shift32_evango_52/io_in[2] xor_shift32_evango_52/io_in[3]
+ xor_shift32_evango_52/io_in[4] xor_shift32_evango_52/io_in[5] xor_shift32_evango_52/io_in[6]
+ xor_shift32_evango_52/io_in[7] xor_shift32_evango_52/io_out[0] xor_shift32_evango_52/io_out[1]
+ xor_shift32_evango_52/io_out[2] xor_shift32_evango_52/io_out[3] xor_shift32_evango_52/io_out[4]
+ xor_shift32_evango_52/io_out[5] xor_shift32_evango_52/io_out[6] xor_shift32_evango_52/io_out[7]
+ scanchain_52/scan_select_in scanchain_53/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_70 scanchain_70/module_data_in[0] scanchain_70/module_data_in[1]
+ scanchain_70/module_data_in[2] scanchain_70/module_data_in[3] scanchain_70/module_data_in[4]
+ scanchain_70/module_data_in[5] scanchain_70/module_data_in[6] scanchain_70/module_data_in[7]
+ scanchain_70/module_data_out[0] scanchain_70/module_data_out[1] scanchain_70/module_data_out[2]
+ scanchain_70/module_data_out[3] scanchain_70/module_data_out[4] scanchain_70/module_data_out[5]
+ scanchain_70/module_data_out[6] scanchain_70/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_81 scanchain_81/module_data_in[0] scanchain_81/module_data_in[1]
+ scanchain_81/module_data_in[2] scanchain_81/module_data_in[3] scanchain_81/module_data_in[4]
+ scanchain_81/module_data_in[5] scanchain_81/module_data_in[6] scanchain_81/module_data_in[7]
+ scanchain_81/module_data_out[0] scanchain_81/module_data_out[1] scanchain_81/module_data_out[2]
+ scanchain_81/module_data_out[3] scanchain_81/module_data_out[4] scanchain_81/module_data_out[5]
+ scanchain_81/module_data_out[6] scanchain_81/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_92 scanchain_92/module_data_in[0] scanchain_92/module_data_in[1]
+ scanchain_92/module_data_in[2] scanchain_92/module_data_in[3] scanchain_92/module_data_in[4]
+ scanchain_92/module_data_in[5] scanchain_92/module_data_in[6] scanchain_92/module_data_in[7]
+ scanchain_92/module_data_out[0] scanchain_92/module_data_out[1] scanchain_92/module_data_out[2]
+ scanchain_92/module_data_out[3] scanchain_92/module_data_out[4] scanchain_92/module_data_out[5]
+ scanchain_92/module_data_out[6] scanchain_92/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_63 scanchain_63/clk_in scanchain_64/clk_in scanchain_63/data_in scanchain_64/data_in
+ scanchain_63/latch_enable_in scanchain_64/latch_enable_in scanchain_63/module_data_in[0]
+ scanchain_63/module_data_in[1] scanchain_63/module_data_in[2] scanchain_63/module_data_in[3]
+ scanchain_63/module_data_in[4] scanchain_63/module_data_in[5] scanchain_63/module_data_in[6]
+ scanchain_63/module_data_in[7] scanchain_63/module_data_out[0] scanchain_63/module_data_out[1]
+ scanchain_63/module_data_out[2] scanchain_63/module_data_out[3] scanchain_63/module_data_out[4]
+ scanchain_63/module_data_out[5] scanchain_63/module_data_out[6] scanchain_63/module_data_out[7]
+ scanchain_63/scan_select_in scanchain_64/scan_select_in vccd1 vssd1 scanchain
Xscanchain_74 scanchain_74/clk_in scanchain_75/clk_in scanchain_74/data_in scanchain_75/data_in
+ scanchain_74/latch_enable_in scanchain_75/latch_enable_in scanchain_74/module_data_in[0]
+ scanchain_74/module_data_in[1] scanchain_74/module_data_in[2] scanchain_74/module_data_in[3]
+ scanchain_74/module_data_in[4] scanchain_74/module_data_in[5] scanchain_74/module_data_in[6]
+ scanchain_74/module_data_in[7] scanchain_74/module_data_out[0] scanchain_74/module_data_out[1]
+ scanchain_74/module_data_out[2] scanchain_74/module_data_out[3] scanchain_74/module_data_out[4]
+ scanchain_74/module_data_out[5] scanchain_74/module_data_out[6] scanchain_74/module_data_out[7]
+ scanchain_74/scan_select_in scanchain_75/scan_select_in vccd1 vssd1 scanchain
Xscanchain_85 scanchain_85/clk_in scanchain_86/clk_in scanchain_85/data_in scanchain_86/data_in
+ scanchain_85/latch_enable_in scanchain_86/latch_enable_in scanchain_85/module_data_in[0]
+ scanchain_85/module_data_in[1] scanchain_85/module_data_in[2] scanchain_85/module_data_in[3]
+ scanchain_85/module_data_in[4] scanchain_85/module_data_in[5] scanchain_85/module_data_in[6]
+ scanchain_85/module_data_in[7] scanchain_85/module_data_out[0] scanchain_85/module_data_out[1]
+ scanchain_85/module_data_out[2] scanchain_85/module_data_out[3] scanchain_85/module_data_out[4]
+ scanchain_85/module_data_out[5] scanchain_85/module_data_out[6] scanchain_85/module_data_out[7]
+ scanchain_85/scan_select_in scanchain_86/scan_select_in vccd1 vssd1 scanchain
Xscanchain_96 scanchain_96/clk_in scanchain_97/clk_in scanchain_96/data_in scanchain_97/data_in
+ scanchain_96/latch_enable_in scanchain_97/latch_enable_in scanchain_96/module_data_in[0]
+ scanchain_96/module_data_in[1] scanchain_96/module_data_in[2] scanchain_96/module_data_in[3]
+ scanchain_96/module_data_in[4] scanchain_96/module_data_in[5] scanchain_96/module_data_in[6]
+ scanchain_96/module_data_in[7] scanchain_96/module_data_out[0] scanchain_96/module_data_out[1]
+ scanchain_96/module_data_out[2] scanchain_96/module_data_out[3] scanchain_96/module_data_out[4]
+ scanchain_96/module_data_out[5] scanchain_96/module_data_out[6] scanchain_96/module_data_out[7]
+ scanchain_96/scan_select_in scanchain_97/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_454 scanchain_454/module_data_in[0] scanchain_454/module_data_in[1]
+ scanchain_454/module_data_in[2] scanchain_454/module_data_in[3] scanchain_454/module_data_in[4]
+ scanchain_454/module_data_in[5] scanchain_454/module_data_in[6] scanchain_454/module_data_in[7]
+ scanchain_454/module_data_out[0] scanchain_454/module_data_out[1] scanchain_454/module_data_out[2]
+ scanchain_454/module_data_out[3] scanchain_454/module_data_out[4] scanchain_454/module_data_out[5]
+ scanchain_454/module_data_out[6] scanchain_454/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_443 scanchain_443/module_data_in[0] scanchain_443/module_data_in[1]
+ scanchain_443/module_data_in[2] scanchain_443/module_data_in[3] scanchain_443/module_data_in[4]
+ scanchain_443/module_data_in[5] scanchain_443/module_data_in[6] scanchain_443/module_data_in[7]
+ scanchain_443/module_data_out[0] scanchain_443/module_data_out[1] scanchain_443/module_data_out[2]
+ scanchain_443/module_data_out[3] scanchain_443/module_data_out[4] scanchain_443/module_data_out[5]
+ scanchain_443/module_data_out[6] scanchain_443/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_432 scanchain_432/module_data_in[0] scanchain_432/module_data_in[1]
+ scanchain_432/module_data_in[2] scanchain_432/module_data_in[3] scanchain_432/module_data_in[4]
+ scanchain_432/module_data_in[5] scanchain_432/module_data_in[6] scanchain_432/module_data_in[7]
+ scanchain_432/module_data_out[0] scanchain_432/module_data_out[1] scanchain_432/module_data_out[2]
+ scanchain_432/module_data_out[3] scanchain_432/module_data_out[4] scanchain_432/module_data_out[5]
+ scanchain_432/module_data_out[6] scanchain_432/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_421 scanchain_421/module_data_in[0] scanchain_421/module_data_in[1]
+ scanchain_421/module_data_in[2] scanchain_421/module_data_in[3] scanchain_421/module_data_in[4]
+ scanchain_421/module_data_in[5] scanchain_421/module_data_in[6] scanchain_421/module_data_in[7]
+ scanchain_421/module_data_out[0] scanchain_421/module_data_out[1] scanchain_421/module_data_out[2]
+ scanchain_421/module_data_out[3] scanchain_421/module_data_out[4] scanchain_421/module_data_out[5]
+ scanchain_421/module_data_out[6] scanchain_421/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_410 scanchain_410/module_data_in[0] scanchain_410/module_data_in[1]
+ scanchain_410/module_data_in[2] scanchain_410/module_data_in[3] scanchain_410/module_data_in[4]
+ scanchain_410/module_data_in[5] scanchain_410/module_data_in[6] scanchain_410/module_data_in[7]
+ scanchain_410/module_data_out[0] scanchain_410/module_data_out[1] scanchain_410/module_data_out[2]
+ scanchain_410/module_data_out[3] scanchain_410/module_data_out[4] scanchain_410/module_data_out[5]
+ scanchain_410/module_data_out[6] scanchain_410/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_465 scanchain_465/module_data_in[0] scanchain_465/module_data_in[1]
+ scanchain_465/module_data_in[2] scanchain_465/module_data_in[3] scanchain_465/module_data_in[4]
+ scanchain_465/module_data_in[5] scanchain_465/module_data_in[6] scanchain_465/module_data_in[7]
+ scanchain_465/module_data_out[0] scanchain_465/module_data_out[1] scanchain_465/module_data_out[2]
+ scanchain_465/module_data_out[3] scanchain_465/module_data_out[4] scanchain_465/module_data_out[5]
+ scanchain_465/module_data_out[6] scanchain_465/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_429 scanchain_429/clk_in scanchain_430/clk_in scanchain_429/data_in scanchain_430/data_in
+ scanchain_429/latch_enable_in scanchain_430/latch_enable_in scanchain_429/module_data_in[0]
+ scanchain_429/module_data_in[1] scanchain_429/module_data_in[2] scanchain_429/module_data_in[3]
+ scanchain_429/module_data_in[4] scanchain_429/module_data_in[5] scanchain_429/module_data_in[6]
+ scanchain_429/module_data_in[7] scanchain_429/module_data_out[0] scanchain_429/module_data_out[1]
+ scanchain_429/module_data_out[2] scanchain_429/module_data_out[3] scanchain_429/module_data_out[4]
+ scanchain_429/module_data_out[5] scanchain_429/module_data_out[6] scanchain_429/module_data_out[7]
+ scanchain_429/scan_select_in scanchain_430/scan_select_in vccd1 vssd1 scanchain
Xscanchain_418 scanchain_418/clk_in scanchain_419/clk_in scanchain_418/data_in scanchain_419/data_in
+ scanchain_418/latch_enable_in scanchain_419/latch_enable_in scanchain_418/module_data_in[0]
+ scanchain_418/module_data_in[1] scanchain_418/module_data_in[2] scanchain_418/module_data_in[3]
+ scanchain_418/module_data_in[4] scanchain_418/module_data_in[5] scanchain_418/module_data_in[6]
+ scanchain_418/module_data_in[7] scanchain_418/module_data_out[0] scanchain_418/module_data_out[1]
+ scanchain_418/module_data_out[2] scanchain_418/module_data_out[3] scanchain_418/module_data_out[4]
+ scanchain_418/module_data_out[5] scanchain_418/module_data_out[6] scanchain_418/module_data_out[7]
+ scanchain_418/scan_select_in scanchain_419/scan_select_in vccd1 vssd1 scanchain
Xscanchain_407 scanchain_407/clk_in scanchain_408/clk_in scanchain_407/data_in scanchain_408/data_in
+ scanchain_407/latch_enable_in scanchain_408/latch_enable_in scanchain_407/module_data_in[0]
+ scanchain_407/module_data_in[1] scanchain_407/module_data_in[2] scanchain_407/module_data_in[3]
+ scanchain_407/module_data_in[4] scanchain_407/module_data_in[5] scanchain_407/module_data_in[6]
+ scanchain_407/module_data_in[7] scanchain_407/module_data_out[0] scanchain_407/module_data_out[1]
+ scanchain_407/module_data_out[2] scanchain_407/module_data_out[3] scanchain_407/module_data_out[4]
+ scanchain_407/module_data_out[5] scanchain_407/module_data_out[6] scanchain_407/module_data_out[7]
+ scanchain_407/scan_select_in scanchain_408/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_284 scanchain_284/module_data_in[0] scanchain_284/module_data_in[1]
+ scanchain_284/module_data_in[2] scanchain_284/module_data_in[3] scanchain_284/module_data_in[4]
+ scanchain_284/module_data_in[5] scanchain_284/module_data_in[6] scanchain_284/module_data_in[7]
+ scanchain_284/module_data_out[0] scanchain_284/module_data_out[1] scanchain_284/module_data_out[2]
+ scanchain_284/module_data_out[3] scanchain_284/module_data_out[4] scanchain_284/module_data_out[5]
+ scanchain_284/module_data_out[6] scanchain_284/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_295 scanchain_295/module_data_in[0] scanchain_295/module_data_in[1]
+ scanchain_295/module_data_in[2] scanchain_295/module_data_in[3] scanchain_295/module_data_in[4]
+ scanchain_295/module_data_in[5] scanchain_295/module_data_in[6] scanchain_295/module_data_in[7]
+ scanchain_295/module_data_out[0] scanchain_295/module_data_out[1] scanchain_295/module_data_out[2]
+ scanchain_295/module_data_out[3] scanchain_295/module_data_out[4] scanchain_295/module_data_out[5]
+ scanchain_295/module_data_out[6] scanchain_295/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_273 scanchain_273/module_data_in[0] scanchain_273/module_data_in[1]
+ scanchain_273/module_data_in[2] scanchain_273/module_data_in[3] scanchain_273/module_data_in[4]
+ scanchain_273/module_data_in[5] scanchain_273/module_data_in[6] scanchain_273/module_data_in[7]
+ scanchain_273/module_data_out[0] scanchain_273/module_data_out[1] scanchain_273/module_data_out[2]
+ scanchain_273/module_data_out[3] scanchain_273/module_data_out[4] scanchain_273/module_data_out[5]
+ scanchain_273/module_data_out[6] scanchain_273/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_251 scanchain_251/module_data_in[0] scanchain_251/module_data_in[1]
+ scanchain_251/module_data_in[2] scanchain_251/module_data_in[3] scanchain_251/module_data_in[4]
+ scanchain_251/module_data_in[5] scanchain_251/module_data_in[6] scanchain_251/module_data_in[7]
+ scanchain_251/module_data_out[0] scanchain_251/module_data_out[1] scanchain_251/module_data_out[2]
+ scanchain_251/module_data_out[3] scanchain_251/module_data_out[4] scanchain_251/module_data_out[5]
+ scanchain_251/module_data_out[6] scanchain_251/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_262 scanchain_262/module_data_in[0] scanchain_262/module_data_in[1]
+ scanchain_262/module_data_in[2] scanchain_262/module_data_in[3] scanchain_262/module_data_in[4]
+ scanchain_262/module_data_in[5] scanchain_262/module_data_in[6] scanchain_262/module_data_in[7]
+ scanchain_262/module_data_out[0] scanchain_262/module_data_out[1] scanchain_262/module_data_out[2]
+ scanchain_262/module_data_out[3] scanchain_262/module_data_out[4] scanchain_262/module_data_out[5]
+ scanchain_262/module_data_out[6] scanchain_262/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_240 scanchain_240/module_data_in[0] scanchain_240/module_data_in[1]
+ scanchain_240/module_data_in[2] scanchain_240/module_data_in[3] scanchain_240/module_data_in[4]
+ scanchain_240/module_data_in[5] scanchain_240/module_data_in[6] scanchain_240/module_data_in[7]
+ scanchain_240/module_data_out[0] scanchain_240/module_data_out[1] scanchain_240/module_data_out[2]
+ scanchain_240/module_data_out[3] scanchain_240/module_data_out[4] scanchain_240/module_data_out[5]
+ scanchain_240/module_data_out[6] scanchain_240/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_248 scanchain_248/clk_in scanchain_249/clk_in scanchain_248/data_in scanchain_249/data_in
+ scanchain_248/latch_enable_in scanchain_249/latch_enable_in scanchain_248/module_data_in[0]
+ scanchain_248/module_data_in[1] scanchain_248/module_data_in[2] scanchain_248/module_data_in[3]
+ scanchain_248/module_data_in[4] scanchain_248/module_data_in[5] scanchain_248/module_data_in[6]
+ scanchain_248/module_data_in[7] scanchain_248/module_data_out[0] scanchain_248/module_data_out[1]
+ scanchain_248/module_data_out[2] scanchain_248/module_data_out[3] scanchain_248/module_data_out[4]
+ scanchain_248/module_data_out[5] scanchain_248/module_data_out[6] scanchain_248/module_data_out[7]
+ scanchain_248/scan_select_in scanchain_249/scan_select_in vccd1 vssd1 scanchain
Xscanchain_259 scanchain_259/clk_in scanchain_260/clk_in scanchain_259/data_in scanchain_260/data_in
+ scanchain_259/latch_enable_in scanchain_260/latch_enable_in scanchain_259/module_data_in[0]
+ scanchain_259/module_data_in[1] scanchain_259/module_data_in[2] scanchain_259/module_data_in[3]
+ scanchain_259/module_data_in[4] scanchain_259/module_data_in[5] scanchain_259/module_data_in[6]
+ scanchain_259/module_data_in[7] scanchain_259/module_data_out[0] scanchain_259/module_data_out[1]
+ scanchain_259/module_data_out[2] scanchain_259/module_data_out[3] scanchain_259/module_data_out[4]
+ scanchain_259/module_data_out[5] scanchain_259/module_data_out[6] scanchain_259/module_data_out[7]
+ scanchain_259/scan_select_in scanchain_260/scan_select_in vccd1 vssd1 scanchain
Xscanchain_237 scanchain_237/clk_in scanchain_238/clk_in scanchain_237/data_in scanchain_238/data_in
+ scanchain_237/latch_enable_in scanchain_238/latch_enable_in scanchain_237/module_data_in[0]
+ scanchain_237/module_data_in[1] scanchain_237/module_data_in[2] scanchain_237/module_data_in[3]
+ scanchain_237/module_data_in[4] scanchain_237/module_data_in[5] scanchain_237/module_data_in[6]
+ scanchain_237/module_data_in[7] scanchain_237/module_data_out[0] scanchain_237/module_data_out[1]
+ scanchain_237/module_data_out[2] scanchain_237/module_data_out[3] scanchain_237/module_data_out[4]
+ scanchain_237/module_data_out[5] scanchain_237/module_data_out[6] scanchain_237/module_data_out[7]
+ scanchain_237/scan_select_in scanchain_238/scan_select_in vccd1 vssd1 scanchain
Xscanchain_226 scanchain_226/clk_in scanchain_227/clk_in scanchain_226/data_in scanchain_227/data_in
+ scanchain_226/latch_enable_in scanchain_227/latch_enable_in scanchain_226/module_data_in[0]
+ scanchain_226/module_data_in[1] scanchain_226/module_data_in[2] scanchain_226/module_data_in[3]
+ scanchain_226/module_data_in[4] scanchain_226/module_data_in[5] scanchain_226/module_data_in[6]
+ scanchain_226/module_data_in[7] scanchain_226/module_data_out[0] scanchain_226/module_data_out[1]
+ scanchain_226/module_data_out[2] scanchain_226/module_data_out[3] scanchain_226/module_data_out[4]
+ scanchain_226/module_data_out[5] scanchain_226/module_data_out[6] scanchain_226/module_data_out[7]
+ scanchain_226/scan_select_in scanchain_227/scan_select_in vccd1 vssd1 scanchain
Xscanchain_215 scanchain_215/clk_in scanchain_216/clk_in scanchain_215/data_in scanchain_216/data_in
+ scanchain_215/latch_enable_in scanchain_216/latch_enable_in scanchain_215/module_data_in[0]
+ scanchain_215/module_data_in[1] scanchain_215/module_data_in[2] scanchain_215/module_data_in[3]
+ scanchain_215/module_data_in[4] scanchain_215/module_data_in[5] scanchain_215/module_data_in[6]
+ scanchain_215/module_data_in[7] scanchain_215/module_data_out[0] scanchain_215/module_data_out[1]
+ scanchain_215/module_data_out[2] scanchain_215/module_data_out[3] scanchain_215/module_data_out[4]
+ scanchain_215/module_data_out[5] scanchain_215/module_data_out[6] scanchain_215/module_data_out[7]
+ scanchain_215/scan_select_in scanchain_216/scan_select_in vccd1 vssd1 scanchain
Xscanchain_204 scanchain_204/clk_in scanchain_205/clk_in scanchain_204/data_in scanchain_205/data_in
+ scanchain_204/latch_enable_in scanchain_205/latch_enable_in scanchain_204/module_data_in[0]
+ scanchain_204/module_data_in[1] scanchain_204/module_data_in[2] scanchain_204/module_data_in[3]
+ scanchain_204/module_data_in[4] scanchain_204/module_data_in[5] scanchain_204/module_data_in[6]
+ scanchain_204/module_data_in[7] scanchain_204/module_data_out[0] scanchain_204/module_data_out[1]
+ scanchain_204/module_data_out[2] scanchain_204/module_data_out[3] scanchain_204/module_data_out[4]
+ scanchain_204/module_data_out[5] scanchain_204/module_data_out[6] scanchain_204/module_data_out[7]
+ scanchain_204/scan_select_in scanchain_205/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_71 scanchain_71/module_data_in[0] scanchain_71/module_data_in[1]
+ scanchain_71/module_data_in[2] scanchain_71/module_data_in[3] scanchain_71/module_data_in[4]
+ scanchain_71/module_data_in[5] scanchain_71/module_data_in[6] scanchain_71/module_data_in[7]
+ scanchain_71/module_data_out[0] scanchain_71/module_data_out[1] scanchain_71/module_data_out[2]
+ scanchain_71/module_data_out[3] scanchain_71/module_data_out[4] scanchain_71/module_data_out[5]
+ scanchain_71/module_data_out[6] scanchain_71/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_60 scanchain_60/module_data_in[0] scanchain_60/module_data_in[1]
+ scanchain_60/module_data_in[2] scanchain_60/module_data_in[3] scanchain_60/module_data_in[4]
+ scanchain_60/module_data_in[5] scanchain_60/module_data_in[6] scanchain_60/module_data_in[7]
+ scanchain_60/module_data_out[0] scanchain_60/module_data_out[1] scanchain_60/module_data_out[2]
+ scanchain_60/module_data_out[3] scanchain_60/module_data_out[4] scanchain_60/module_data_out[5]
+ scanchain_60/module_data_out[6] scanchain_60/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_82 scanchain_82/module_data_in[0] scanchain_82/module_data_in[1]
+ scanchain_82/module_data_in[2] scanchain_82/module_data_in[3] scanchain_82/module_data_in[4]
+ scanchain_82/module_data_in[5] scanchain_82/module_data_in[6] scanchain_82/module_data_in[7]
+ scanchain_82/module_data_out[0] scanchain_82/module_data_out[1] scanchain_82/module_data_out[2]
+ scanchain_82/module_data_out[3] scanchain_82/module_data_out[4] scanchain_82/module_data_out[5]
+ scanchain_82/module_data_out[6] scanchain_82/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_93 scanchain_93/module_data_in[0] scanchain_93/module_data_in[1]
+ scanchain_93/module_data_in[2] scanchain_93/module_data_in[3] scanchain_93/module_data_in[4]
+ scanchain_93/module_data_in[5] scanchain_93/module_data_in[6] scanchain_93/module_data_in[7]
+ scanchain_93/module_data_out[0] scanchain_93/module_data_out[1] scanchain_93/module_data_out[2]
+ scanchain_93/module_data_out[3] scanchain_93/module_data_out[4] scanchain_93/module_data_out[5]
+ scanchain_93/module_data_out[6] scanchain_93/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_42 scanchain_42/clk_in scanchain_43/clk_in scanchain_42/data_in scanchain_43/data_in
+ scanchain_42/latch_enable_in scanchain_43/latch_enable_in top_42/io_in[0] top_42/io_in[1]
+ top_42/io_in[2] top_42/io_in[3] top_42/io_in[4] top_42/io_in[5] top_42/io_in[6]
+ top_42/io_in[7] top_42/io_out[0] top_42/io_out[1] top_42/io_out[2] top_42/io_out[3]
+ top_42/io_out[4] top_42/io_out[5] top_42/io_out[6] top_42/io_out[7] scanchain_42/scan_select_in
+ scanchain_43/scan_select_in vccd1 vssd1 scanchain
Xscanchain_20 scanchain_20/clk_in scanchain_21/clk_in scanchain_20/data_in scanchain_21/data_in
+ scanchain_20/latch_enable_in scanchain_21/latch_enable_in chase_the_beat_20/io_in[0]
+ chase_the_beat_20/io_in[1] chase_the_beat_20/io_in[2] chase_the_beat_20/io_in[3]
+ chase_the_beat_20/io_in[4] chase_the_beat_20/io_in[5] chase_the_beat_20/io_in[6]
+ chase_the_beat_20/io_in[7] chase_the_beat_20/io_out[0] chase_the_beat_20/io_out[1]
+ chase_the_beat_20/io_out[2] chase_the_beat_20/io_out[3] chase_the_beat_20/io_out[4]
+ chase_the_beat_20/io_out[5] chase_the_beat_20/io_out[6] chase_the_beat_20/io_out[7]
+ scanchain_20/scan_select_in scanchain_21/scan_select_in vccd1 vssd1 scanchain
Xscanchain_31 scanchain_31/clk_in scanchain_32/clk_in scanchain_31/data_in scanchain_32/data_in
+ scanchain_31/latch_enable_in scanchain_32/latch_enable_in zoechip_31/io_in[0] zoechip_31/io_in[1]
+ zoechip_31/io_in[2] zoechip_31/io_in[3] zoechip_31/io_in[4] zoechip_31/io_in[5]
+ zoechip_31/io_in[6] zoechip_31/io_in[7] zoechip_31/io_out[0] zoechip_31/io_out[1]
+ zoechip_31/io_out[2] zoechip_31/io_out[3] zoechip_31/io_out[4] zoechip_31/io_out[5]
+ zoechip_31/io_out[6] zoechip_31/io_out[7] scanchain_31/scan_select_in scanchain_32/scan_select_in
+ vccd1 vssd1 scanchain
Xscanchain_53 scanchain_53/clk_in scanchain_54/clk_in scanchain_53/data_in scanchain_54/data_in
+ scanchain_53/latch_enable_in scanchain_54/latch_enable_in scanchain_53/module_data_in[0]
+ scanchain_53/module_data_in[1] scanchain_53/module_data_in[2] scanchain_53/module_data_in[3]
+ scanchain_53/module_data_in[4] scanchain_53/module_data_in[5] scanchain_53/module_data_in[6]
+ scanchain_53/module_data_in[7] scanchain_53/module_data_out[0] scanchain_53/module_data_out[1]
+ scanchain_53/module_data_out[2] scanchain_53/module_data_out[3] scanchain_53/module_data_out[4]
+ scanchain_53/module_data_out[5] scanchain_53/module_data_out[6] scanchain_53/module_data_out[7]
+ scanchain_53/scan_select_in scanchain_54/scan_select_in vccd1 vssd1 scanchain
Xscanchain_64 scanchain_64/clk_in scanchain_65/clk_in scanchain_64/data_in scanchain_65/data_in
+ scanchain_64/latch_enable_in scanchain_65/latch_enable_in scanchain_64/module_data_in[0]
+ scanchain_64/module_data_in[1] scanchain_64/module_data_in[2] scanchain_64/module_data_in[3]
+ scanchain_64/module_data_in[4] scanchain_64/module_data_in[5] scanchain_64/module_data_in[6]
+ scanchain_64/module_data_in[7] scanchain_64/module_data_out[0] scanchain_64/module_data_out[1]
+ scanchain_64/module_data_out[2] scanchain_64/module_data_out[3] scanchain_64/module_data_out[4]
+ scanchain_64/module_data_out[5] scanchain_64/module_data_out[6] scanchain_64/module_data_out[7]
+ scanchain_64/scan_select_in scanchain_65/scan_select_in vccd1 vssd1 scanchain
Xscanchain_75 scanchain_75/clk_in scanchain_76/clk_in scanchain_75/data_in scanchain_76/data_in
+ scanchain_75/latch_enable_in scanchain_76/latch_enable_in scanchain_75/module_data_in[0]
+ scanchain_75/module_data_in[1] scanchain_75/module_data_in[2] scanchain_75/module_data_in[3]
+ scanchain_75/module_data_in[4] scanchain_75/module_data_in[5] scanchain_75/module_data_in[6]
+ scanchain_75/module_data_in[7] scanchain_75/module_data_out[0] scanchain_75/module_data_out[1]
+ scanchain_75/module_data_out[2] scanchain_75/module_data_out[3] scanchain_75/module_data_out[4]
+ scanchain_75/module_data_out[5] scanchain_75/module_data_out[6] scanchain_75/module_data_out[7]
+ scanchain_75/scan_select_in scanchain_76/scan_select_in vccd1 vssd1 scanchain
Xscanchain_86 scanchain_86/clk_in scanchain_87/clk_in scanchain_86/data_in scanchain_87/data_in
+ scanchain_86/latch_enable_in scanchain_87/latch_enable_in scanchain_86/module_data_in[0]
+ scanchain_86/module_data_in[1] scanchain_86/module_data_in[2] scanchain_86/module_data_in[3]
+ scanchain_86/module_data_in[4] scanchain_86/module_data_in[5] scanchain_86/module_data_in[6]
+ scanchain_86/module_data_in[7] scanchain_86/module_data_out[0] scanchain_86/module_data_out[1]
+ scanchain_86/module_data_out[2] scanchain_86/module_data_out[3] scanchain_86/module_data_out[4]
+ scanchain_86/module_data_out[5] scanchain_86/module_data_out[6] scanchain_86/module_data_out[7]
+ scanchain_86/scan_select_in scanchain_87/scan_select_in vccd1 vssd1 scanchain
Xscanchain_97 scanchain_97/clk_in scanchain_98/clk_in scanchain_97/data_in scanchain_98/data_in
+ scanchain_97/latch_enable_in scanchain_98/latch_enable_in scanchain_97/module_data_in[0]
+ scanchain_97/module_data_in[1] scanchain_97/module_data_in[2] scanchain_97/module_data_in[3]
+ scanchain_97/module_data_in[4] scanchain_97/module_data_in[5] scanchain_97/module_data_in[6]
+ scanchain_97/module_data_in[7] scanchain_97/module_data_out[0] scanchain_97/module_data_out[1]
+ scanchain_97/module_data_out[2] scanchain_97/module_data_out[3] scanchain_97/module_data_out[4]
+ scanchain_97/module_data_out[5] scanchain_97/module_data_out[6] scanchain_97/module_data_out[7]
+ scanchain_97/scan_select_in scanchain_98/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_466 scanchain_466/module_data_in[0] scanchain_466/module_data_in[1]
+ scanchain_466/module_data_in[2] scanchain_466/module_data_in[3] scanchain_466/module_data_in[4]
+ scanchain_466/module_data_in[5] scanchain_466/module_data_in[6] scanchain_466/module_data_in[7]
+ scanchain_466/module_data_out[0] scanchain_466/module_data_out[1] scanchain_466/module_data_out[2]
+ scanchain_466/module_data_out[3] scanchain_466/module_data_out[4] scanchain_466/module_data_out[5]
+ scanchain_466/module_data_out[6] scanchain_466/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_455 scanchain_455/module_data_in[0] scanchain_455/module_data_in[1]
+ scanchain_455/module_data_in[2] scanchain_455/module_data_in[3] scanchain_455/module_data_in[4]
+ scanchain_455/module_data_in[5] scanchain_455/module_data_in[6] scanchain_455/module_data_in[7]
+ scanchain_455/module_data_out[0] scanchain_455/module_data_out[1] scanchain_455/module_data_out[2]
+ scanchain_455/module_data_out[3] scanchain_455/module_data_out[4] scanchain_455/module_data_out[5]
+ scanchain_455/module_data_out[6] scanchain_455/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_444 scanchain_444/module_data_in[0] scanchain_444/module_data_in[1]
+ scanchain_444/module_data_in[2] scanchain_444/module_data_in[3] scanchain_444/module_data_in[4]
+ scanchain_444/module_data_in[5] scanchain_444/module_data_in[6] scanchain_444/module_data_in[7]
+ scanchain_444/module_data_out[0] scanchain_444/module_data_out[1] scanchain_444/module_data_out[2]
+ scanchain_444/module_data_out[3] scanchain_444/module_data_out[4] scanchain_444/module_data_out[5]
+ scanchain_444/module_data_out[6] scanchain_444/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_433 scanchain_433/module_data_in[0] scanchain_433/module_data_in[1]
+ scanchain_433/module_data_in[2] scanchain_433/module_data_in[3] scanchain_433/module_data_in[4]
+ scanchain_433/module_data_in[5] scanchain_433/module_data_in[6] scanchain_433/module_data_in[7]
+ scanchain_433/module_data_out[0] scanchain_433/module_data_out[1] scanchain_433/module_data_out[2]
+ scanchain_433/module_data_out[3] scanchain_433/module_data_out[4] scanchain_433/module_data_out[5]
+ scanchain_433/module_data_out[6] scanchain_433/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_422 scanchain_422/module_data_in[0] scanchain_422/module_data_in[1]
+ scanchain_422/module_data_in[2] scanchain_422/module_data_in[3] scanchain_422/module_data_in[4]
+ scanchain_422/module_data_in[5] scanchain_422/module_data_in[6] scanchain_422/module_data_in[7]
+ scanchain_422/module_data_out[0] scanchain_422/module_data_out[1] scanchain_422/module_data_out[2]
+ scanchain_422/module_data_out[3] scanchain_422/module_data_out[4] scanchain_422/module_data_out[5]
+ scanchain_422/module_data_out[6] scanchain_422/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_419 scanchain_419/clk_in scanchain_420/clk_in scanchain_419/data_in scanchain_420/data_in
+ scanchain_419/latch_enable_in scanchain_420/latch_enable_in scanchain_419/module_data_in[0]
+ scanchain_419/module_data_in[1] scanchain_419/module_data_in[2] scanchain_419/module_data_in[3]
+ scanchain_419/module_data_in[4] scanchain_419/module_data_in[5] scanchain_419/module_data_in[6]
+ scanchain_419/module_data_in[7] scanchain_419/module_data_out[0] scanchain_419/module_data_out[1]
+ scanchain_419/module_data_out[2] scanchain_419/module_data_out[3] scanchain_419/module_data_out[4]
+ scanchain_419/module_data_out[5] scanchain_419/module_data_out[6] scanchain_419/module_data_out[7]
+ scanchain_419/scan_select_in scanchain_420/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_400 scanchain_400/module_data_in[0] scanchain_400/module_data_in[1]
+ scanchain_400/module_data_in[2] scanchain_400/module_data_in[3] scanchain_400/module_data_in[4]
+ scanchain_400/module_data_in[5] scanchain_400/module_data_in[6] scanchain_400/module_data_in[7]
+ scanchain_400/module_data_out[0] scanchain_400/module_data_out[1] scanchain_400/module_data_out[2]
+ scanchain_400/module_data_out[3] scanchain_400/module_data_out[4] scanchain_400/module_data_out[5]
+ scanchain_400/module_data_out[6] scanchain_400/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_408 scanchain_408/clk_in scanchain_409/clk_in scanchain_408/data_in scanchain_409/data_in
+ scanchain_408/latch_enable_in scanchain_409/latch_enable_in scanchain_408/module_data_in[0]
+ scanchain_408/module_data_in[1] scanchain_408/module_data_in[2] scanchain_408/module_data_in[3]
+ scanchain_408/module_data_in[4] scanchain_408/module_data_in[5] scanchain_408/module_data_in[6]
+ scanchain_408/module_data_in[7] scanchain_408/module_data_out[0] scanchain_408/module_data_out[1]
+ scanchain_408/module_data_out[2] scanchain_408/module_data_out[3] scanchain_408/module_data_out[4]
+ scanchain_408/module_data_out[5] scanchain_408/module_data_out[6] scanchain_408/module_data_out[7]
+ scanchain_408/scan_select_in scanchain_409/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_411 scanchain_411/module_data_in[0] scanchain_411/module_data_in[1]
+ scanchain_411/module_data_in[2] scanchain_411/module_data_in[3] scanchain_411/module_data_in[4]
+ scanchain_411/module_data_in[5] scanchain_411/module_data_in[6] scanchain_411/module_data_in[7]
+ scanchain_411/module_data_out[0] scanchain_411/module_data_out[1] scanchain_411/module_data_out[2]
+ scanchain_411/module_data_out[3] scanchain_411/module_data_out[4] scanchain_411/module_data_out[5]
+ scanchain_411/module_data_out[6] scanchain_411/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_285 scanchain_285/module_data_in[0] scanchain_285/module_data_in[1]
+ scanchain_285/module_data_in[2] scanchain_285/module_data_in[3] scanchain_285/module_data_in[4]
+ scanchain_285/module_data_in[5] scanchain_285/module_data_in[6] scanchain_285/module_data_in[7]
+ scanchain_285/module_data_out[0] scanchain_285/module_data_out[1] scanchain_285/module_data_out[2]
+ scanchain_285/module_data_out[3] scanchain_285/module_data_out[4] scanchain_285/module_data_out[5]
+ scanchain_285/module_data_out[6] scanchain_285/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_296 scanchain_296/module_data_in[0] scanchain_296/module_data_in[1]
+ scanchain_296/module_data_in[2] scanchain_296/module_data_in[3] scanchain_296/module_data_in[4]
+ scanchain_296/module_data_in[5] scanchain_296/module_data_in[6] scanchain_296/module_data_in[7]
+ scanchain_296/module_data_out[0] scanchain_296/module_data_out[1] scanchain_296/module_data_out[2]
+ scanchain_296/module_data_out[3] scanchain_296/module_data_out[4] scanchain_296/module_data_out[5]
+ scanchain_296/module_data_out[6] scanchain_296/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_274 scanchain_274/module_data_in[0] scanchain_274/module_data_in[1]
+ scanchain_274/module_data_in[2] scanchain_274/module_data_in[3] scanchain_274/module_data_in[4]
+ scanchain_274/module_data_in[5] scanchain_274/module_data_in[6] scanchain_274/module_data_in[7]
+ scanchain_274/module_data_out[0] scanchain_274/module_data_out[1] scanchain_274/module_data_out[2]
+ scanchain_274/module_data_out[3] scanchain_274/module_data_out[4] scanchain_274/module_data_out[5]
+ scanchain_274/module_data_out[6] scanchain_274/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_252 scanchain_252/module_data_in[0] scanchain_252/module_data_in[1]
+ scanchain_252/module_data_in[2] scanchain_252/module_data_in[3] scanchain_252/module_data_in[4]
+ scanchain_252/module_data_in[5] scanchain_252/module_data_in[6] scanchain_252/module_data_in[7]
+ scanchain_252/module_data_out[0] scanchain_252/module_data_out[1] scanchain_252/module_data_out[2]
+ scanchain_252/module_data_out[3] scanchain_252/module_data_out[4] scanchain_252/module_data_out[5]
+ scanchain_252/module_data_out[6] scanchain_252/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_263 scanchain_263/module_data_in[0] scanchain_263/module_data_in[1]
+ scanchain_263/module_data_in[2] scanchain_263/module_data_in[3] scanchain_263/module_data_in[4]
+ scanchain_263/module_data_in[5] scanchain_263/module_data_in[6] scanchain_263/module_data_in[7]
+ scanchain_263/module_data_out[0] scanchain_263/module_data_out[1] scanchain_263/module_data_out[2]
+ scanchain_263/module_data_out[3] scanchain_263/module_data_out[4] scanchain_263/module_data_out[5]
+ scanchain_263/module_data_out[6] scanchain_263/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_241 scanchain_241/module_data_in[0] scanchain_241/module_data_in[1]
+ scanchain_241/module_data_in[2] scanchain_241/module_data_in[3] scanchain_241/module_data_in[4]
+ scanchain_241/module_data_in[5] scanchain_241/module_data_in[6] scanchain_241/module_data_in[7]
+ scanchain_241/module_data_out[0] scanchain_241/module_data_out[1] scanchain_241/module_data_out[2]
+ scanchain_241/module_data_out[3] scanchain_241/module_data_out[4] scanchain_241/module_data_out[5]
+ scanchain_241/module_data_out[6] scanchain_241/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_230 scanchain_230/module_data_in[0] scanchain_230/module_data_in[1]
+ scanchain_230/module_data_in[2] scanchain_230/module_data_in[3] scanchain_230/module_data_in[4]
+ scanchain_230/module_data_in[5] scanchain_230/module_data_in[6] scanchain_230/module_data_in[7]
+ scanchain_230/module_data_out[0] scanchain_230/module_data_out[1] scanchain_230/module_data_out[2]
+ scanchain_230/module_data_out[3] scanchain_230/module_data_out[4] scanchain_230/module_data_out[5]
+ scanchain_230/module_data_out[6] scanchain_230/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_249 scanchain_249/clk_in scanchain_250/clk_in scanchain_249/data_in scanchain_250/data_in
+ scanchain_249/latch_enable_in scanchain_250/latch_enable_in scanchain_249/module_data_in[0]
+ scanchain_249/module_data_in[1] scanchain_249/module_data_in[2] scanchain_249/module_data_in[3]
+ scanchain_249/module_data_in[4] scanchain_249/module_data_in[5] scanchain_249/module_data_in[6]
+ scanchain_249/module_data_in[7] scanchain_249/module_data_out[0] scanchain_249/module_data_out[1]
+ scanchain_249/module_data_out[2] scanchain_249/module_data_out[3] scanchain_249/module_data_out[4]
+ scanchain_249/module_data_out[5] scanchain_249/module_data_out[6] scanchain_249/module_data_out[7]
+ scanchain_249/scan_select_in scanchain_250/scan_select_in vccd1 vssd1 scanchain
Xscanchain_238 scanchain_238/clk_in scanchain_239/clk_in scanchain_238/data_in scanchain_239/data_in
+ scanchain_238/latch_enable_in scanchain_239/latch_enable_in scanchain_238/module_data_in[0]
+ scanchain_238/module_data_in[1] scanchain_238/module_data_in[2] scanchain_238/module_data_in[3]
+ scanchain_238/module_data_in[4] scanchain_238/module_data_in[5] scanchain_238/module_data_in[6]
+ scanchain_238/module_data_in[7] scanchain_238/module_data_out[0] scanchain_238/module_data_out[1]
+ scanchain_238/module_data_out[2] scanchain_238/module_data_out[3] scanchain_238/module_data_out[4]
+ scanchain_238/module_data_out[5] scanchain_238/module_data_out[6] scanchain_238/module_data_out[7]
+ scanchain_238/scan_select_in scanchain_239/scan_select_in vccd1 vssd1 scanchain
Xscanchain_227 scanchain_227/clk_in scanchain_228/clk_in scanchain_227/data_in scanchain_228/data_in
+ scanchain_227/latch_enable_in scanchain_228/latch_enable_in scanchain_227/module_data_in[0]
+ scanchain_227/module_data_in[1] scanchain_227/module_data_in[2] scanchain_227/module_data_in[3]
+ scanchain_227/module_data_in[4] scanchain_227/module_data_in[5] scanchain_227/module_data_in[6]
+ scanchain_227/module_data_in[7] scanchain_227/module_data_out[0] scanchain_227/module_data_out[1]
+ scanchain_227/module_data_out[2] scanchain_227/module_data_out[3] scanchain_227/module_data_out[4]
+ scanchain_227/module_data_out[5] scanchain_227/module_data_out[6] scanchain_227/module_data_out[7]
+ scanchain_227/scan_select_in scanchain_228/scan_select_in vccd1 vssd1 scanchain
Xscanchain_216 scanchain_216/clk_in scanchain_217/clk_in scanchain_216/data_in scanchain_217/data_in
+ scanchain_216/latch_enable_in scanchain_217/latch_enable_in scanchain_216/module_data_in[0]
+ scanchain_216/module_data_in[1] scanchain_216/module_data_in[2] scanchain_216/module_data_in[3]
+ scanchain_216/module_data_in[4] scanchain_216/module_data_in[5] scanchain_216/module_data_in[6]
+ scanchain_216/module_data_in[7] scanchain_216/module_data_out[0] scanchain_216/module_data_out[1]
+ scanchain_216/module_data_out[2] scanchain_216/module_data_out[3] scanchain_216/module_data_out[4]
+ scanchain_216/module_data_out[5] scanchain_216/module_data_out[6] scanchain_216/module_data_out[7]
+ scanchain_216/scan_select_in scanchain_217/scan_select_in vccd1 vssd1 scanchain
Xscanchain_205 scanchain_205/clk_in scanchain_206/clk_in scanchain_205/data_in scanchain_206/data_in
+ scanchain_205/latch_enable_in scanchain_206/latch_enable_in scanchain_205/module_data_in[0]
+ scanchain_205/module_data_in[1] scanchain_205/module_data_in[2] scanchain_205/module_data_in[3]
+ scanchain_205/module_data_in[4] scanchain_205/module_data_in[5] scanchain_205/module_data_in[6]
+ scanchain_205/module_data_in[7] scanchain_205/module_data_out[0] scanchain_205/module_data_out[1]
+ scanchain_205/module_data_out[2] scanchain_205/module_data_out[3] scanchain_205/module_data_out[4]
+ scanchain_205/module_data_out[5] scanchain_205/module_data_out[6] scanchain_205/module_data_out[7]
+ scanchain_205/scan_select_in scanchain_206/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_72 scanchain_72/module_data_in[0] scanchain_72/module_data_in[1]
+ scanchain_72/module_data_in[2] scanchain_72/module_data_in[3] scanchain_72/module_data_in[4]
+ scanchain_72/module_data_in[5] scanchain_72/module_data_in[6] scanchain_72/module_data_in[7]
+ scanchain_72/module_data_out[0] scanchain_72/module_data_out[1] scanchain_72/module_data_out[2]
+ scanchain_72/module_data_out[3] scanchain_72/module_data_out[4] scanchain_72/module_data_out[5]
+ scanchain_72/module_data_out[6] scanchain_72/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_61 scanchain_61/module_data_in[0] scanchain_61/module_data_in[1]
+ scanchain_61/module_data_in[2] scanchain_61/module_data_in[3] scanchain_61/module_data_in[4]
+ scanchain_61/module_data_in[5] scanchain_61/module_data_in[6] scanchain_61/module_data_in[7]
+ scanchain_61/module_data_out[0] scanchain_61/module_data_out[1] scanchain_61/module_data_out[2]
+ scanchain_61/module_data_out[3] scanchain_61/module_data_out[4] scanchain_61/module_data_out[5]
+ scanchain_61/module_data_out[6] scanchain_61/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_83 scanchain_83/module_data_in[0] scanchain_83/module_data_in[1]
+ scanchain_83/module_data_in[2] scanchain_83/module_data_in[3] scanchain_83/module_data_in[4]
+ scanchain_83/module_data_in[5] scanchain_83/module_data_in[6] scanchain_83/module_data_in[7]
+ scanchain_83/module_data_out[0] scanchain_83/module_data_out[1] scanchain_83/module_data_out[2]
+ scanchain_83/module_data_out[3] scanchain_83/module_data_out[4] scanchain_83/module_data_out[5]
+ scanchain_83/module_data_out[6] scanchain_83/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_94 scanchain_94/module_data_in[0] scanchain_94/module_data_in[1]
+ scanchain_94/module_data_in[2] scanchain_94/module_data_in[3] scanchain_94/module_data_in[4]
+ scanchain_94/module_data_in[5] scanchain_94/module_data_in[6] scanchain_94/module_data_in[7]
+ scanchain_94/module_data_out[0] scanchain_94/module_data_out[1] scanchain_94/module_data_out[2]
+ scanchain_94/module_data_out[3] scanchain_94/module_data_out[4] scanchain_94/module_data_out[5]
+ scanchain_94/module_data_out[6] scanchain_94/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_43 scanchain_43/clk_in scanchain_44/clk_in scanchain_43/data_in scanchain_44/data_in
+ scanchain_43/latch_enable_in scanchain_44/latch_enable_in rc5_top_43/io_in[0] rc5_top_43/io_in[1]
+ rc5_top_43/io_in[2] rc5_top_43/io_in[3] rc5_top_43/io_in[4] rc5_top_43/io_in[5]
+ rc5_top_43/io_in[6] rc5_top_43/io_in[7] rc5_top_43/io_out[0] rc5_top_43/io_out[1]
+ rc5_top_43/io_out[2] rc5_top_43/io_out[3] rc5_top_43/io_out[4] rc5_top_43/io_out[5]
+ rc5_top_43/io_out[6] rc5_top_43/io_out[7] scanchain_43/scan_select_in scanchain_44/scan_select_in
+ vccd1 vssd1 scanchain
Xscanchain_21 scanchain_21/clk_in scanchain_22/clk_in scanchain_21/data_in scanchain_22/data_in
+ scanchain_21/latch_enable_in scanchain_22/latch_enable_in scanchain_21/module_data_in[0]
+ scanchain_21/module_data_in[1] scanchain_21/module_data_in[2] scanchain_21/module_data_in[3]
+ scanchain_21/module_data_in[4] scanchain_21/module_data_in[5] scanchain_21/module_data_in[6]
+ scanchain_21/module_data_in[7] scanchain_21/module_data_out[0] scanchain_21/module_data_out[1]
+ scanchain_21/module_data_out[2] scanchain_21/module_data_out[3] scanchain_21/module_data_out[4]
+ scanchain_21/module_data_out[5] scanchain_21/module_data_out[6] scanchain_21/module_data_out[7]
+ scanchain_21/scan_select_in scanchain_22/scan_select_in vccd1 vssd1 scanchain
Xscanchain_32 scanchain_32/clk_in scanchain_33/clk_in scanchain_32/data_in scanchain_33/data_in
+ scanchain_32/latch_enable_in scanchain_33/latch_enable_in scanchain_32/module_data_in[0]
+ scanchain_32/module_data_in[1] scanchain_32/module_data_in[2] scanchain_32/module_data_in[3]
+ scanchain_32/module_data_in[4] scanchain_32/module_data_in[5] scanchain_32/module_data_in[6]
+ scanchain_32/module_data_in[7] scanchain_32/module_data_out[0] scanchain_32/module_data_out[1]
+ scanchain_32/module_data_out[2] scanchain_32/module_data_out[3] scanchain_32/module_data_out[4]
+ scanchain_32/module_data_out[5] scanchain_32/module_data_out[6] scanchain_32/module_data_out[7]
+ scanchain_32/scan_select_in scanchain_33/scan_select_in vccd1 vssd1 scanchain
Xscanchain_10 scanchain_9/clk_out scanchain_11/clk_in scanchain_9/data_out scanchain_11/data_in
+ scanchain_9/latch_enable_out scanchain_11/latch_enable_in scanchain_10/module_data_in[0]
+ scanchain_10/module_data_in[1] scanchain_10/module_data_in[2] scanchain_10/module_data_in[3]
+ scanchain_10/module_data_in[4] scanchain_10/module_data_in[5] scanchain_10/module_data_in[6]
+ scanchain_10/module_data_in[7] scanchain_10/module_data_out[0] scanchain_10/module_data_out[1]
+ scanchain_10/module_data_out[2] scanchain_10/module_data_out[3] scanchain_10/module_data_out[4]
+ scanchain_10/module_data_out[5] scanchain_10/module_data_out[6] scanchain_10/module_data_out[7]
+ scanchain_9/scan_select_out scanchain_11/scan_select_in vccd1 vssd1 scanchain
Xscanchain_54 scanchain_54/clk_in scanchain_55/clk_in scanchain_54/data_in scanchain_55/data_in
+ scanchain_54/latch_enable_in scanchain_55/latch_enable_in jleightcap_top_54/io_in[0]
+ jleightcap_top_54/io_in[1] jleightcap_top_54/io_in[2] jleightcap_top_54/io_in[3]
+ jleightcap_top_54/io_in[4] jleightcap_top_54/io_in[5] jleightcap_top_54/io_in[6]
+ jleightcap_top_54/io_in[7] jleightcap_top_54/io_out[0] jleightcap_top_54/io_out[1]
+ jleightcap_top_54/io_out[2] jleightcap_top_54/io_out[3] jleightcap_top_54/io_out[4]
+ jleightcap_top_54/io_out[5] jleightcap_top_54/io_out[6] jleightcap_top_54/io_out[7]
+ scanchain_54/scan_select_in scanchain_55/scan_select_in vccd1 vssd1 scanchain
Xscanchain_65 scanchain_65/clk_in scanchain_66/clk_in scanchain_65/data_in scanchain_66/data_in
+ scanchain_65/latch_enable_in scanchain_66/latch_enable_in scanchain_65/module_data_in[0]
+ scanchain_65/module_data_in[1] scanchain_65/module_data_in[2] scanchain_65/module_data_in[3]
+ scanchain_65/module_data_in[4] scanchain_65/module_data_in[5] scanchain_65/module_data_in[6]
+ scanchain_65/module_data_in[7] scanchain_65/module_data_out[0] scanchain_65/module_data_out[1]
+ scanchain_65/module_data_out[2] scanchain_65/module_data_out[3] scanchain_65/module_data_out[4]
+ scanchain_65/module_data_out[5] scanchain_65/module_data_out[6] scanchain_65/module_data_out[7]
+ scanchain_65/scan_select_in scanchain_66/scan_select_in vccd1 vssd1 scanchain
Xscanchain_76 scanchain_76/clk_in scanchain_77/clk_in scanchain_76/data_in scanchain_77/data_in
+ scanchain_76/latch_enable_in scanchain_77/latch_enable_in scanchain_76/module_data_in[0]
+ scanchain_76/module_data_in[1] scanchain_76/module_data_in[2] scanchain_76/module_data_in[3]
+ scanchain_76/module_data_in[4] scanchain_76/module_data_in[5] scanchain_76/module_data_in[6]
+ scanchain_76/module_data_in[7] scanchain_76/module_data_out[0] scanchain_76/module_data_out[1]
+ scanchain_76/module_data_out[2] scanchain_76/module_data_out[3] scanchain_76/module_data_out[4]
+ scanchain_76/module_data_out[5] scanchain_76/module_data_out[6] scanchain_76/module_data_out[7]
+ scanchain_76/scan_select_in scanchain_77/scan_select_in vccd1 vssd1 scanchain
Xscanchain_87 scanchain_87/clk_in scanchain_88/clk_in scanchain_87/data_in scanchain_88/data_in
+ scanchain_87/latch_enable_in scanchain_88/latch_enable_in scanchain_87/module_data_in[0]
+ scanchain_87/module_data_in[1] scanchain_87/module_data_in[2] scanchain_87/module_data_in[3]
+ scanchain_87/module_data_in[4] scanchain_87/module_data_in[5] scanchain_87/module_data_in[6]
+ scanchain_87/module_data_in[7] scanchain_87/module_data_out[0] scanchain_87/module_data_out[1]
+ scanchain_87/module_data_out[2] scanchain_87/module_data_out[3] scanchain_87/module_data_out[4]
+ scanchain_87/module_data_out[5] scanchain_87/module_data_out[6] scanchain_87/module_data_out[7]
+ scanchain_87/scan_select_in scanchain_88/scan_select_in vccd1 vssd1 scanchain
Xscanchain_98 scanchain_98/clk_in scanchain_99/clk_in scanchain_98/data_in scanchain_99/data_in
+ scanchain_98/latch_enable_in scanchain_99/latch_enable_in scanchain_98/module_data_in[0]
+ scanchain_98/module_data_in[1] scanchain_98/module_data_in[2] scanchain_98/module_data_in[3]
+ scanchain_98/module_data_in[4] scanchain_98/module_data_in[5] scanchain_98/module_data_in[6]
+ scanchain_98/module_data_in[7] scanchain_98/module_data_out[0] scanchain_98/module_data_out[1]
+ scanchain_98/module_data_out[2] scanchain_98/module_data_out[3] scanchain_98/module_data_out[4]
+ scanchain_98/module_data_out[5] scanchain_98/module_data_out[6] scanchain_98/module_data_out[7]
+ scanchain_98/scan_select_in scanchain_99/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_467 scanchain_467/module_data_in[0] scanchain_467/module_data_in[1]
+ scanchain_467/module_data_in[2] scanchain_467/module_data_in[3] scanchain_467/module_data_in[4]
+ scanchain_467/module_data_in[5] scanchain_467/module_data_in[6] scanchain_467/module_data_in[7]
+ scanchain_467/module_data_out[0] scanchain_467/module_data_out[1] scanchain_467/module_data_out[2]
+ scanchain_467/module_data_out[3] scanchain_467/module_data_out[4] scanchain_467/module_data_out[5]
+ scanchain_467/module_data_out[6] scanchain_467/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_456 scanchain_456/module_data_in[0] scanchain_456/module_data_in[1]
+ scanchain_456/module_data_in[2] scanchain_456/module_data_in[3] scanchain_456/module_data_in[4]
+ scanchain_456/module_data_in[5] scanchain_456/module_data_in[6] scanchain_456/module_data_in[7]
+ scanchain_456/module_data_out[0] scanchain_456/module_data_out[1] scanchain_456/module_data_out[2]
+ scanchain_456/module_data_out[3] scanchain_456/module_data_out[4] scanchain_456/module_data_out[5]
+ scanchain_456/module_data_out[6] scanchain_456/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_445 scanchain_445/module_data_in[0] scanchain_445/module_data_in[1]
+ scanchain_445/module_data_in[2] scanchain_445/module_data_in[3] scanchain_445/module_data_in[4]
+ scanchain_445/module_data_in[5] scanchain_445/module_data_in[6] scanchain_445/module_data_in[7]
+ scanchain_445/module_data_out[0] scanchain_445/module_data_out[1] scanchain_445/module_data_out[2]
+ scanchain_445/module_data_out[3] scanchain_445/module_data_out[4] scanchain_445/module_data_out[5]
+ scanchain_445/module_data_out[6] scanchain_445/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_434 scanchain_434/module_data_in[0] scanchain_434/module_data_in[1]
+ scanchain_434/module_data_in[2] scanchain_434/module_data_in[3] scanchain_434/module_data_in[4]
+ scanchain_434/module_data_in[5] scanchain_434/module_data_in[6] scanchain_434/module_data_in[7]
+ scanchain_434/module_data_out[0] scanchain_434/module_data_out[1] scanchain_434/module_data_out[2]
+ scanchain_434/module_data_out[3] scanchain_434/module_data_out[4] scanchain_434/module_data_out[5]
+ scanchain_434/module_data_out[6] scanchain_434/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_423 scanchain_423/module_data_in[0] scanchain_423/module_data_in[1]
+ scanchain_423/module_data_in[2] scanchain_423/module_data_in[3] scanchain_423/module_data_in[4]
+ scanchain_423/module_data_in[5] scanchain_423/module_data_in[6] scanchain_423/module_data_in[7]
+ scanchain_423/module_data_out[0] scanchain_423/module_data_out[1] scanchain_423/module_data_out[2]
+ scanchain_423/module_data_out[3] scanchain_423/module_data_out[4] scanchain_423/module_data_out[5]
+ scanchain_423/module_data_out[6] scanchain_423/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_401 scanchain_401/module_data_in[0] scanchain_401/module_data_in[1]
+ scanchain_401/module_data_in[2] scanchain_401/module_data_in[3] scanchain_401/module_data_in[4]
+ scanchain_401/module_data_in[5] scanchain_401/module_data_in[6] scanchain_401/module_data_in[7]
+ scanchain_401/module_data_out[0] scanchain_401/module_data_out[1] scanchain_401/module_data_out[2]
+ scanchain_401/module_data_out[3] scanchain_401/module_data_out[4] scanchain_401/module_data_out[5]
+ scanchain_401/module_data_out[6] scanchain_401/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_409 scanchain_409/clk_in scanchain_410/clk_in scanchain_409/data_in scanchain_410/data_in
+ scanchain_409/latch_enable_in scanchain_410/latch_enable_in scanchain_409/module_data_in[0]
+ scanchain_409/module_data_in[1] scanchain_409/module_data_in[2] scanchain_409/module_data_in[3]
+ scanchain_409/module_data_in[4] scanchain_409/module_data_in[5] scanchain_409/module_data_in[6]
+ scanchain_409/module_data_in[7] scanchain_409/module_data_out[0] scanchain_409/module_data_out[1]
+ scanchain_409/module_data_out[2] scanchain_409/module_data_out[3] scanchain_409/module_data_out[4]
+ scanchain_409/module_data_out[5] scanchain_409/module_data_out[6] scanchain_409/module_data_out[7]
+ scanchain_409/scan_select_in scanchain_410/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_412 scanchain_412/module_data_in[0] scanchain_412/module_data_in[1]
+ scanchain_412/module_data_in[2] scanchain_412/module_data_in[3] scanchain_412/module_data_in[4]
+ scanchain_412/module_data_in[5] scanchain_412/module_data_in[6] scanchain_412/module_data_in[7]
+ scanchain_412/module_data_out[0] scanchain_412/module_data_out[1] scanchain_412/module_data_out[2]
+ scanchain_412/module_data_out[3] scanchain_412/module_data_out[4] scanchain_412/module_data_out[5]
+ scanchain_412/module_data_out[6] scanchain_412/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_220 scanchain_220/module_data_in[0] scanchain_220/module_data_in[1]
+ scanchain_220/module_data_in[2] scanchain_220/module_data_in[3] scanchain_220/module_data_in[4]
+ scanchain_220/module_data_in[5] scanchain_220/module_data_in[6] scanchain_220/module_data_in[7]
+ scanchain_220/module_data_out[0] scanchain_220/module_data_out[1] scanchain_220/module_data_out[2]
+ scanchain_220/module_data_out[3] scanchain_220/module_data_out[4] scanchain_220/module_data_out[5]
+ scanchain_220/module_data_out[6] scanchain_220/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_286 scanchain_286/module_data_in[0] scanchain_286/module_data_in[1]
+ scanchain_286/module_data_in[2] scanchain_286/module_data_in[3] scanchain_286/module_data_in[4]
+ scanchain_286/module_data_in[5] scanchain_286/module_data_in[6] scanchain_286/module_data_in[7]
+ scanchain_286/module_data_out[0] scanchain_286/module_data_out[1] scanchain_286/module_data_out[2]
+ scanchain_286/module_data_out[3] scanchain_286/module_data_out[4] scanchain_286/module_data_out[5]
+ scanchain_286/module_data_out[6] scanchain_286/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_297 scanchain_297/module_data_in[0] scanchain_297/module_data_in[1]
+ scanchain_297/module_data_in[2] scanchain_297/module_data_in[3] scanchain_297/module_data_in[4]
+ scanchain_297/module_data_in[5] scanchain_297/module_data_in[6] scanchain_297/module_data_in[7]
+ scanchain_297/module_data_out[0] scanchain_297/module_data_out[1] scanchain_297/module_data_out[2]
+ scanchain_297/module_data_out[3] scanchain_297/module_data_out[4] scanchain_297/module_data_out[5]
+ scanchain_297/module_data_out[6] scanchain_297/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_275 scanchain_275/module_data_in[0] scanchain_275/module_data_in[1]
+ scanchain_275/module_data_in[2] scanchain_275/module_data_in[3] scanchain_275/module_data_in[4]
+ scanchain_275/module_data_in[5] scanchain_275/module_data_in[6] scanchain_275/module_data_in[7]
+ scanchain_275/module_data_out[0] scanchain_275/module_data_out[1] scanchain_275/module_data_out[2]
+ scanchain_275/module_data_out[3] scanchain_275/module_data_out[4] scanchain_275/module_data_out[5]
+ scanchain_275/module_data_out[6] scanchain_275/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_264 scanchain_264/module_data_in[0] scanchain_264/module_data_in[1]
+ scanchain_264/module_data_in[2] scanchain_264/module_data_in[3] scanchain_264/module_data_in[4]
+ scanchain_264/module_data_in[5] scanchain_264/module_data_in[6] scanchain_264/module_data_in[7]
+ scanchain_264/module_data_out[0] scanchain_264/module_data_out[1] scanchain_264/module_data_out[2]
+ scanchain_264/module_data_out[3] scanchain_264/module_data_out[4] scanchain_264/module_data_out[5]
+ scanchain_264/module_data_out[6] scanchain_264/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_253 scanchain_253/module_data_in[0] scanchain_253/module_data_in[1]
+ scanchain_253/module_data_in[2] scanchain_253/module_data_in[3] scanchain_253/module_data_in[4]
+ scanchain_253/module_data_in[5] scanchain_253/module_data_in[6] scanchain_253/module_data_in[7]
+ scanchain_253/module_data_out[0] scanchain_253/module_data_out[1] scanchain_253/module_data_out[2]
+ scanchain_253/module_data_out[3] scanchain_253/module_data_out[4] scanchain_253/module_data_out[5]
+ scanchain_253/module_data_out[6] scanchain_253/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_242 scanchain_242/module_data_in[0] scanchain_242/module_data_in[1]
+ scanchain_242/module_data_in[2] scanchain_242/module_data_in[3] scanchain_242/module_data_in[4]
+ scanchain_242/module_data_in[5] scanchain_242/module_data_in[6] scanchain_242/module_data_in[7]
+ scanchain_242/module_data_out[0] scanchain_242/module_data_out[1] scanchain_242/module_data_out[2]
+ scanchain_242/module_data_out[3] scanchain_242/module_data_out[4] scanchain_242/module_data_out[5]
+ scanchain_242/module_data_out[6] scanchain_242/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_239 scanchain_239/clk_in scanchain_240/clk_in scanchain_239/data_in scanchain_240/data_in
+ scanchain_239/latch_enable_in scanchain_240/latch_enable_in scanchain_239/module_data_in[0]
+ scanchain_239/module_data_in[1] scanchain_239/module_data_in[2] scanchain_239/module_data_in[3]
+ scanchain_239/module_data_in[4] scanchain_239/module_data_in[5] scanchain_239/module_data_in[6]
+ scanchain_239/module_data_in[7] scanchain_239/module_data_out[0] scanchain_239/module_data_out[1]
+ scanchain_239/module_data_out[2] scanchain_239/module_data_out[3] scanchain_239/module_data_out[4]
+ scanchain_239/module_data_out[5] scanchain_239/module_data_out[6] scanchain_239/module_data_out[7]
+ scanchain_239/scan_select_in scanchain_240/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_231 scanchain_231/module_data_in[0] scanchain_231/module_data_in[1]
+ scanchain_231/module_data_in[2] scanchain_231/module_data_in[3] scanchain_231/module_data_in[4]
+ scanchain_231/module_data_in[5] scanchain_231/module_data_in[6] scanchain_231/module_data_in[7]
+ scanchain_231/module_data_out[0] scanchain_231/module_data_out[1] scanchain_231/module_data_out[2]
+ scanchain_231/module_data_out[3] scanchain_231/module_data_out[4] scanchain_231/module_data_out[5]
+ scanchain_231/module_data_out[6] scanchain_231/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_228 scanchain_228/clk_in scanchain_229/clk_in scanchain_228/data_in scanchain_229/data_in
+ scanchain_228/latch_enable_in scanchain_229/latch_enable_in scanchain_228/module_data_in[0]
+ scanchain_228/module_data_in[1] scanchain_228/module_data_in[2] scanchain_228/module_data_in[3]
+ scanchain_228/module_data_in[4] scanchain_228/module_data_in[5] scanchain_228/module_data_in[6]
+ scanchain_228/module_data_in[7] scanchain_228/module_data_out[0] scanchain_228/module_data_out[1]
+ scanchain_228/module_data_out[2] scanchain_228/module_data_out[3] scanchain_228/module_data_out[4]
+ scanchain_228/module_data_out[5] scanchain_228/module_data_out[6] scanchain_228/module_data_out[7]
+ scanchain_228/scan_select_in scanchain_229/scan_select_in vccd1 vssd1 scanchain
Xscanchain_217 scanchain_217/clk_in scanchain_218/clk_in scanchain_217/data_in scanchain_218/data_in
+ scanchain_217/latch_enable_in scanchain_218/latch_enable_in scanchain_217/module_data_in[0]
+ scanchain_217/module_data_in[1] scanchain_217/module_data_in[2] scanchain_217/module_data_in[3]
+ scanchain_217/module_data_in[4] scanchain_217/module_data_in[5] scanchain_217/module_data_in[6]
+ scanchain_217/module_data_in[7] scanchain_217/module_data_out[0] scanchain_217/module_data_out[1]
+ scanchain_217/module_data_out[2] scanchain_217/module_data_out[3] scanchain_217/module_data_out[4]
+ scanchain_217/module_data_out[5] scanchain_217/module_data_out[6] scanchain_217/module_data_out[7]
+ scanchain_217/scan_select_in scanchain_218/scan_select_in vccd1 vssd1 scanchain
Xscanchain_206 scanchain_206/clk_in scanchain_207/clk_in scanchain_206/data_in scanchain_207/data_in
+ scanchain_206/latch_enable_in scanchain_207/latch_enable_in scanchain_206/module_data_in[0]
+ scanchain_206/module_data_in[1] scanchain_206/module_data_in[2] scanchain_206/module_data_in[3]
+ scanchain_206/module_data_in[4] scanchain_206/module_data_in[5] scanchain_206/module_data_in[6]
+ scanchain_206/module_data_in[7] scanchain_206/module_data_out[0] scanchain_206/module_data_out[1]
+ scanchain_206/module_data_out[2] scanchain_206/module_data_out[3] scanchain_206/module_data_out[4]
+ scanchain_206/module_data_out[5] scanchain_206/module_data_out[6] scanchain_206/module_data_out[7]
+ scanchain_206/scan_select_in scanchain_207/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_73 scanchain_73/module_data_in[0] scanchain_73/module_data_in[1]
+ scanchain_73/module_data_in[2] scanchain_73/module_data_in[3] scanchain_73/module_data_in[4]
+ scanchain_73/module_data_in[5] scanchain_73/module_data_in[6] scanchain_73/module_data_in[7]
+ scanchain_73/module_data_out[0] scanchain_73/module_data_out[1] scanchain_73/module_data_out[2]
+ scanchain_73/module_data_out[3] scanchain_73/module_data_out[4] scanchain_73/module_data_out[5]
+ scanchain_73/module_data_out[6] scanchain_73/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_62 scanchain_62/module_data_in[0] scanchain_62/module_data_in[1]
+ scanchain_62/module_data_in[2] scanchain_62/module_data_in[3] scanchain_62/module_data_in[4]
+ scanchain_62/module_data_in[5] scanchain_62/module_data_in[6] scanchain_62/module_data_in[7]
+ scanchain_62/module_data_out[0] scanchain_62/module_data_out[1] scanchain_62/module_data_out[2]
+ scanchain_62/module_data_out[3] scanchain_62/module_data_out[4] scanchain_62/module_data_out[5]
+ scanchain_62/module_data_out[6] scanchain_62/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_84 scanchain_84/module_data_in[0] scanchain_84/module_data_in[1]
+ scanchain_84/module_data_in[2] scanchain_84/module_data_in[3] scanchain_84/module_data_in[4]
+ scanchain_84/module_data_in[5] scanchain_84/module_data_in[6] scanchain_84/module_data_in[7]
+ scanchain_84/module_data_out[0] scanchain_84/module_data_out[1] scanchain_84/module_data_out[2]
+ scanchain_84/module_data_out[3] scanchain_84/module_data_out[4] scanchain_84/module_data_out[5]
+ scanchain_84/module_data_out[6] scanchain_84/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_95 scanchain_95/module_data_in[0] scanchain_95/module_data_in[1]
+ scanchain_95/module_data_in[2] scanchain_95/module_data_in[3] scanchain_95/module_data_in[4]
+ scanchain_95/module_data_in[5] scanchain_95/module_data_in[6] scanchain_95/module_data_in[7]
+ scanchain_95/module_data_out[0] scanchain_95/module_data_out[1] scanchain_95/module_data_out[2]
+ scanchain_95/module_data_out[3] scanchain_95/module_data_out[4] scanchain_95/module_data_out[5]
+ scanchain_95/module_data_out[6] scanchain_95/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_44 scanchain_44/clk_in scanchain_45/clk_in scanchain_44/data_in scanchain_45/data_in
+ scanchain_44/latch_enable_in scanchain_45/latch_enable_in scanchain_44/module_data_in[0]
+ scanchain_44/module_data_in[1] scanchain_44/module_data_in[2] scanchain_44/module_data_in[3]
+ scanchain_44/module_data_in[4] scanchain_44/module_data_in[5] scanchain_44/module_data_in[6]
+ scanchain_44/module_data_in[7] scanchain_44/module_data_out[0] scanchain_44/module_data_out[1]
+ scanchain_44/module_data_out[2] scanchain_44/module_data_out[3] scanchain_44/module_data_out[4]
+ scanchain_44/module_data_out[5] scanchain_44/module_data_out[6] scanchain_44/module_data_out[7]
+ scanchain_44/scan_select_in scanchain_45/scan_select_in vccd1 vssd1 scanchain
Xscanchain_22 scanchain_22/clk_in scanchain_23/clk_in scanchain_22/data_in scanchain_23/data_in
+ scanchain_22/latch_enable_in scanchain_23/latch_enable_in scanchain_22/module_data_in[0]
+ scanchain_22/module_data_in[1] scanchain_22/module_data_in[2] scanchain_22/module_data_in[3]
+ scanchain_22/module_data_in[4] scanchain_22/module_data_in[5] scanchain_22/module_data_in[6]
+ scanchain_22/module_data_in[7] scanchain_22/module_data_out[0] scanchain_22/module_data_out[1]
+ scanchain_22/module_data_out[2] scanchain_22/module_data_out[3] scanchain_22/module_data_out[4]
+ scanchain_22/module_data_out[5] scanchain_22/module_data_out[6] scanchain_22/module_data_out[7]
+ scanchain_22/scan_select_in scanchain_23/scan_select_in vccd1 vssd1 scanchain
Xscanchain_33 scanchain_33/clk_in scanchain_34/clk_in scanchain_33/data_in scanchain_34/data_in
+ scanchain_33/latch_enable_in scanchain_34/latch_enable_in mbikovitsky_top_33/io_in[0]
+ mbikovitsky_top_33/io_in[1] mbikovitsky_top_33/io_in[2] mbikovitsky_top_33/io_in[3]
+ mbikovitsky_top_33/io_in[4] mbikovitsky_top_33/io_in[5] mbikovitsky_top_33/io_in[6]
+ mbikovitsky_top_33/io_in[7] mbikovitsky_top_33/io_out[0] mbikovitsky_top_33/io_out[1]
+ mbikovitsky_top_33/io_out[2] mbikovitsky_top_33/io_out[3] mbikovitsky_top_33/io_out[4]
+ mbikovitsky_top_33/io_out[5] mbikovitsky_top_33/io_out[6] mbikovitsky_top_33/io_out[7]
+ scanchain_33/scan_select_in scanchain_34/scan_select_in vccd1 vssd1 scanchain
Xscanchain_11 scanchain_11/clk_in scanchain_12/clk_in scanchain_11/data_in scanchain_12/data_in
+ scanchain_11/latch_enable_in scanchain_12/latch_enable_in jar_sram_top_11/io_in[0]
+ jar_sram_top_11/io_in[1] jar_sram_top_11/io_in[2] jar_sram_top_11/io_in[3] jar_sram_top_11/io_in[4]
+ jar_sram_top_11/io_in[5] jar_sram_top_11/io_in[6] jar_sram_top_11/io_in[7] jar_sram_top_11/io_out[0]
+ jar_sram_top_11/io_out[1] jar_sram_top_11/io_out[2] jar_sram_top_11/io_out[3] jar_sram_top_11/io_out[4]
+ jar_sram_top_11/io_out[5] jar_sram_top_11/io_out[6] jar_sram_top_11/io_out[7] scanchain_11/scan_select_in
+ scanchain_12/scan_select_in vccd1 vssd1 scanchain
Xscanchain_66 scanchain_66/clk_in scanchain_67/clk_in scanchain_66/data_in scanchain_67/data_in
+ scanchain_66/latch_enable_in scanchain_67/latch_enable_in scanchain_66/module_data_in[0]
+ scanchain_66/module_data_in[1] scanchain_66/module_data_in[2] scanchain_66/module_data_in[3]
+ scanchain_66/module_data_in[4] scanchain_66/module_data_in[5] scanchain_66/module_data_in[6]
+ scanchain_66/module_data_in[7] scanchain_66/module_data_out[0] scanchain_66/module_data_out[1]
+ scanchain_66/module_data_out[2] scanchain_66/module_data_out[3] scanchain_66/module_data_out[4]
+ scanchain_66/module_data_out[5] scanchain_66/module_data_out[6] scanchain_66/module_data_out[7]
+ scanchain_66/scan_select_in scanchain_67/scan_select_in vccd1 vssd1 scanchain
Xscanchain_55 scanchain_55/clk_in scanchain_56/clk_in scanchain_55/data_in scanchain_56/data_in
+ scanchain_55/latch_enable_in scanchain_56/latch_enable_in scanchain_55/module_data_in[0]
+ scanchain_55/module_data_in[1] scanchain_55/module_data_in[2] scanchain_55/module_data_in[3]
+ scanchain_55/module_data_in[4] scanchain_55/module_data_in[5] scanchain_55/module_data_in[6]
+ scanchain_55/module_data_in[7] scanchain_55/module_data_out[0] scanchain_55/module_data_out[1]
+ scanchain_55/module_data_out[2] scanchain_55/module_data_out[3] scanchain_55/module_data_out[4]
+ scanchain_55/module_data_out[5] scanchain_55/module_data_out[6] scanchain_55/module_data_out[7]
+ scanchain_55/scan_select_in scanchain_56/scan_select_in vccd1 vssd1 scanchain
Xscanchain_77 scanchain_77/clk_in scanchain_78/clk_in scanchain_77/data_in scanchain_78/data_in
+ scanchain_77/latch_enable_in scanchain_78/latch_enable_in scanchain_77/module_data_in[0]
+ scanchain_77/module_data_in[1] scanchain_77/module_data_in[2] scanchain_77/module_data_in[3]
+ scanchain_77/module_data_in[4] scanchain_77/module_data_in[5] scanchain_77/module_data_in[6]
+ scanchain_77/module_data_in[7] scanchain_77/module_data_out[0] scanchain_77/module_data_out[1]
+ scanchain_77/module_data_out[2] scanchain_77/module_data_out[3] scanchain_77/module_data_out[4]
+ scanchain_77/module_data_out[5] scanchain_77/module_data_out[6] scanchain_77/module_data_out[7]
+ scanchain_77/scan_select_in scanchain_78/scan_select_in vccd1 vssd1 scanchain
Xscanchain_88 scanchain_88/clk_in scanchain_89/clk_in scanchain_88/data_in scanchain_89/data_in
+ scanchain_88/latch_enable_in scanchain_89/latch_enable_in scanchain_88/module_data_in[0]
+ scanchain_88/module_data_in[1] scanchain_88/module_data_in[2] scanchain_88/module_data_in[3]
+ scanchain_88/module_data_in[4] scanchain_88/module_data_in[5] scanchain_88/module_data_in[6]
+ scanchain_88/module_data_in[7] scanchain_88/module_data_out[0] scanchain_88/module_data_out[1]
+ scanchain_88/module_data_out[2] scanchain_88/module_data_out[3] scanchain_88/module_data_out[4]
+ scanchain_88/module_data_out[5] scanchain_88/module_data_out[6] scanchain_88/module_data_out[7]
+ scanchain_88/scan_select_in scanchain_89/scan_select_in vccd1 vssd1 scanchain
Xscanchain_99 scanchain_99/clk_in scanchain_99/clk_out scanchain_99/data_in scanchain_99/data_out
+ scanchain_99/latch_enable_in scanchain_99/latch_enable_out scanchain_99/module_data_in[0]
+ scanchain_99/module_data_in[1] scanchain_99/module_data_in[2] scanchain_99/module_data_in[3]
+ scanchain_99/module_data_in[4] scanchain_99/module_data_in[5] scanchain_99/module_data_in[6]
+ scanchain_99/module_data_in[7] scanchain_99/module_data_out[0] scanchain_99/module_data_out[1]
+ scanchain_99/module_data_out[2] scanchain_99/module_data_out[3] scanchain_99/module_data_out[4]
+ scanchain_99/module_data_out[5] scanchain_99/module_data_out[6] scanchain_99/module_data_out[7]
+ scanchain_99/scan_select_in scanchain_99/scan_select_out vccd1 vssd1 scanchain
Xuser_module_339501025136214612_468 scanchain_468/module_data_in[0] scanchain_468/module_data_in[1]
+ scanchain_468/module_data_in[2] scanchain_468/module_data_in[3] scanchain_468/module_data_in[4]
+ scanchain_468/module_data_in[5] scanchain_468/module_data_in[6] scanchain_468/module_data_in[7]
+ scanchain_468/module_data_out[0] scanchain_468/module_data_out[1] scanchain_468/module_data_out[2]
+ scanchain_468/module_data_out[3] scanchain_468/module_data_out[4] scanchain_468/module_data_out[5]
+ scanchain_468/module_data_out[6] scanchain_468/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_457 scanchain_457/module_data_in[0] scanchain_457/module_data_in[1]
+ scanchain_457/module_data_in[2] scanchain_457/module_data_in[3] scanchain_457/module_data_in[4]
+ scanchain_457/module_data_in[5] scanchain_457/module_data_in[6] scanchain_457/module_data_in[7]
+ scanchain_457/module_data_out[0] scanchain_457/module_data_out[1] scanchain_457/module_data_out[2]
+ scanchain_457/module_data_out[3] scanchain_457/module_data_out[4] scanchain_457/module_data_out[5]
+ scanchain_457/module_data_out[6] scanchain_457/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_435 scanchain_435/module_data_in[0] scanchain_435/module_data_in[1]
+ scanchain_435/module_data_in[2] scanchain_435/module_data_in[3] scanchain_435/module_data_in[4]
+ scanchain_435/module_data_in[5] scanchain_435/module_data_in[6] scanchain_435/module_data_in[7]
+ scanchain_435/module_data_out[0] scanchain_435/module_data_out[1] scanchain_435/module_data_out[2]
+ scanchain_435/module_data_out[3] scanchain_435/module_data_out[4] scanchain_435/module_data_out[5]
+ scanchain_435/module_data_out[6] scanchain_435/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_446 scanchain_446/module_data_in[0] scanchain_446/module_data_in[1]
+ scanchain_446/module_data_in[2] scanchain_446/module_data_in[3] scanchain_446/module_data_in[4]
+ scanchain_446/module_data_in[5] scanchain_446/module_data_in[6] scanchain_446/module_data_in[7]
+ scanchain_446/module_data_out[0] scanchain_446/module_data_out[1] scanchain_446/module_data_out[2]
+ scanchain_446/module_data_out[3] scanchain_446/module_data_out[4] scanchain_446/module_data_out[5]
+ scanchain_446/module_data_out[6] scanchain_446/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_424 scanchain_424/module_data_in[0] scanchain_424/module_data_in[1]
+ scanchain_424/module_data_in[2] scanchain_424/module_data_in[3] scanchain_424/module_data_in[4]
+ scanchain_424/module_data_in[5] scanchain_424/module_data_in[6] scanchain_424/module_data_in[7]
+ scanchain_424/module_data_out[0] scanchain_424/module_data_out[1] scanchain_424/module_data_out[2]
+ scanchain_424/module_data_out[3] scanchain_424/module_data_out[4] scanchain_424/module_data_out[5]
+ scanchain_424/module_data_out[6] scanchain_424/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_402 scanchain_402/module_data_in[0] scanchain_402/module_data_in[1]
+ scanchain_402/module_data_in[2] scanchain_402/module_data_in[3] scanchain_402/module_data_in[4]
+ scanchain_402/module_data_in[5] scanchain_402/module_data_in[6] scanchain_402/module_data_in[7]
+ scanchain_402/module_data_out[0] scanchain_402/module_data_out[1] scanchain_402/module_data_out[2]
+ scanchain_402/module_data_out[3] scanchain_402/module_data_out[4] scanchain_402/module_data_out[5]
+ scanchain_402/module_data_out[6] scanchain_402/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_413 scanchain_413/module_data_in[0] scanchain_413/module_data_in[1]
+ scanchain_413/module_data_in[2] scanchain_413/module_data_in[3] scanchain_413/module_data_in[4]
+ scanchain_413/module_data_in[5] scanchain_413/module_data_in[6] scanchain_413/module_data_in[7]
+ scanchain_413/module_data_out[0] scanchain_413/module_data_out[1] scanchain_413/module_data_out[2]
+ scanchain_413/module_data_out[3] scanchain_413/module_data_out[4] scanchain_413/module_data_out[5]
+ scanchain_413/module_data_out[6] scanchain_413/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_287 scanchain_287/module_data_in[0] scanchain_287/module_data_in[1]
+ scanchain_287/module_data_in[2] scanchain_287/module_data_in[3] scanchain_287/module_data_in[4]
+ scanchain_287/module_data_in[5] scanchain_287/module_data_in[6] scanchain_287/module_data_in[7]
+ scanchain_287/module_data_out[0] scanchain_287/module_data_out[1] scanchain_287/module_data_out[2]
+ scanchain_287/module_data_out[3] scanchain_287/module_data_out[4] scanchain_287/module_data_out[5]
+ scanchain_287/module_data_out[6] scanchain_287/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_298 scanchain_298/module_data_in[0] scanchain_298/module_data_in[1]
+ scanchain_298/module_data_in[2] scanchain_298/module_data_in[3] scanchain_298/module_data_in[4]
+ scanchain_298/module_data_in[5] scanchain_298/module_data_in[6] scanchain_298/module_data_in[7]
+ scanchain_298/module_data_out[0] scanchain_298/module_data_out[1] scanchain_298/module_data_out[2]
+ scanchain_298/module_data_out[3] scanchain_298/module_data_out[4] scanchain_298/module_data_out[5]
+ scanchain_298/module_data_out[6] scanchain_298/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_276 scanchain_276/module_data_in[0] scanchain_276/module_data_in[1]
+ scanchain_276/module_data_in[2] scanchain_276/module_data_in[3] scanchain_276/module_data_in[4]
+ scanchain_276/module_data_in[5] scanchain_276/module_data_in[6] scanchain_276/module_data_in[7]
+ scanchain_276/module_data_out[0] scanchain_276/module_data_out[1] scanchain_276/module_data_out[2]
+ scanchain_276/module_data_out[3] scanchain_276/module_data_out[4] scanchain_276/module_data_out[5]
+ scanchain_276/module_data_out[6] scanchain_276/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_265 scanchain_265/module_data_in[0] scanchain_265/module_data_in[1]
+ scanchain_265/module_data_in[2] scanchain_265/module_data_in[3] scanchain_265/module_data_in[4]
+ scanchain_265/module_data_in[5] scanchain_265/module_data_in[6] scanchain_265/module_data_in[7]
+ scanchain_265/module_data_out[0] scanchain_265/module_data_out[1] scanchain_265/module_data_out[2]
+ scanchain_265/module_data_out[3] scanchain_265/module_data_out[4] scanchain_265/module_data_out[5]
+ scanchain_265/module_data_out[6] scanchain_265/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_254 scanchain_254/module_data_in[0] scanchain_254/module_data_in[1]
+ scanchain_254/module_data_in[2] scanchain_254/module_data_in[3] scanchain_254/module_data_in[4]
+ scanchain_254/module_data_in[5] scanchain_254/module_data_in[6] scanchain_254/module_data_in[7]
+ scanchain_254/module_data_out[0] scanchain_254/module_data_out[1] scanchain_254/module_data_out[2]
+ scanchain_254/module_data_out[3] scanchain_254/module_data_out[4] scanchain_254/module_data_out[5]
+ scanchain_254/module_data_out[6] scanchain_254/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_243 scanchain_243/module_data_in[0] scanchain_243/module_data_in[1]
+ scanchain_243/module_data_in[2] scanchain_243/module_data_in[3] scanchain_243/module_data_in[4]
+ scanchain_243/module_data_in[5] scanchain_243/module_data_in[6] scanchain_243/module_data_in[7]
+ scanchain_243/module_data_out[0] scanchain_243/module_data_out[1] scanchain_243/module_data_out[2]
+ scanchain_243/module_data_out[3] scanchain_243/module_data_out[4] scanchain_243/module_data_out[5]
+ scanchain_243/module_data_out[6] scanchain_243/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_232 scanchain_232/module_data_in[0] scanchain_232/module_data_in[1]
+ scanchain_232/module_data_in[2] scanchain_232/module_data_in[3] scanchain_232/module_data_in[4]
+ scanchain_232/module_data_in[5] scanchain_232/module_data_in[6] scanchain_232/module_data_in[7]
+ scanchain_232/module_data_out[0] scanchain_232/module_data_out[1] scanchain_232/module_data_out[2]
+ scanchain_232/module_data_out[3] scanchain_232/module_data_out[4] scanchain_232/module_data_out[5]
+ scanchain_232/module_data_out[6] scanchain_232/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_229 scanchain_229/clk_in scanchain_230/clk_in scanchain_229/data_in scanchain_230/data_in
+ scanchain_229/latch_enable_in scanchain_230/latch_enable_in scanchain_229/module_data_in[0]
+ scanchain_229/module_data_in[1] scanchain_229/module_data_in[2] scanchain_229/module_data_in[3]
+ scanchain_229/module_data_in[4] scanchain_229/module_data_in[5] scanchain_229/module_data_in[6]
+ scanchain_229/module_data_in[7] scanchain_229/module_data_out[0] scanchain_229/module_data_out[1]
+ scanchain_229/module_data_out[2] scanchain_229/module_data_out[3] scanchain_229/module_data_out[4]
+ scanchain_229/module_data_out[5] scanchain_229/module_data_out[6] scanchain_229/module_data_out[7]
+ scanchain_229/scan_select_in scanchain_230/scan_select_in vccd1 vssd1 scanchain
Xscanchain_207 scanchain_207/clk_in scanchain_208/clk_in scanchain_207/data_in scanchain_208/data_in
+ scanchain_207/latch_enable_in scanchain_208/latch_enable_in scanchain_207/module_data_in[0]
+ scanchain_207/module_data_in[1] scanchain_207/module_data_in[2] scanchain_207/module_data_in[3]
+ scanchain_207/module_data_in[4] scanchain_207/module_data_in[5] scanchain_207/module_data_in[6]
+ scanchain_207/module_data_in[7] scanchain_207/module_data_out[0] scanchain_207/module_data_out[1]
+ scanchain_207/module_data_out[2] scanchain_207/module_data_out[3] scanchain_207/module_data_out[4]
+ scanchain_207/module_data_out[5] scanchain_207/module_data_out[6] scanchain_207/module_data_out[7]
+ scanchain_207/scan_select_in scanchain_208/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_210 scanchain_210/module_data_in[0] scanchain_210/module_data_in[1]
+ scanchain_210/module_data_in[2] scanchain_210/module_data_in[3] scanchain_210/module_data_in[4]
+ scanchain_210/module_data_in[5] scanchain_210/module_data_in[6] scanchain_210/module_data_in[7]
+ scanchain_210/module_data_out[0] scanchain_210/module_data_out[1] scanchain_210/module_data_out[2]
+ scanchain_210/module_data_out[3] scanchain_210/module_data_out[4] scanchain_210/module_data_out[5]
+ scanchain_210/module_data_out[6] scanchain_210/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_218 scanchain_218/clk_in scanchain_219/clk_in scanchain_218/data_in scanchain_219/data_in
+ scanchain_218/latch_enable_in scanchain_219/latch_enable_in scanchain_218/module_data_in[0]
+ scanchain_218/module_data_in[1] scanchain_218/module_data_in[2] scanchain_218/module_data_in[3]
+ scanchain_218/module_data_in[4] scanchain_218/module_data_in[5] scanchain_218/module_data_in[6]
+ scanchain_218/module_data_in[7] scanchain_218/module_data_out[0] scanchain_218/module_data_out[1]
+ scanchain_218/module_data_out[2] scanchain_218/module_data_out[3] scanchain_218/module_data_out[4]
+ scanchain_218/module_data_out[5] scanchain_218/module_data_out[6] scanchain_218/module_data_out[7]
+ scanchain_218/scan_select_in scanchain_219/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_221 scanchain_221/module_data_in[0] scanchain_221/module_data_in[1]
+ scanchain_221/module_data_in[2] scanchain_221/module_data_in[3] scanchain_221/module_data_in[4]
+ scanchain_221/module_data_in[5] scanchain_221/module_data_in[6] scanchain_221/module_data_in[7]
+ scanchain_221/module_data_out[0] scanchain_221/module_data_out[1] scanchain_221/module_data_out[2]
+ scanchain_221/module_data_out[3] scanchain_221/module_data_out[4] scanchain_221/module_data_out[5]
+ scanchain_221/module_data_out[6] scanchain_221/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_341516949939814994_48 scanchain_48/module_data_in[0] scanchain_48/module_data_in[1]
+ scanchain_48/module_data_in[2] scanchain_48/module_data_in[3] scanchain_48/module_data_in[4]
+ scanchain_48/module_data_in[5] scanchain_48/module_data_in[6] scanchain_48/module_data_in[7]
+ scanchain_48/module_data_out[0] scanchain_48/module_data_out[1] scanchain_48/module_data_out[2]
+ scanchain_48/module_data_out[3] scanchain_48/module_data_out[4] scanchain_48/module_data_out[5]
+ scanchain_48/module_data_out[6] scanchain_48/module_data_out[7] vccd1 vssd1 user_module_341516949939814994
Xrolfmobile99_alu_fsm_top_35 scanchain_35/module_data_in[0] scanchain_35/module_data_in[1]
+ scanchain_35/module_data_in[2] scanchain_35/module_data_in[3] scanchain_35/module_data_in[4]
+ scanchain_35/module_data_in[5] scanchain_35/module_data_in[6] scanchain_35/module_data_in[7]
+ scanchain_35/module_data_out[0] scanchain_35/module_data_out[1] scanchain_35/module_data_out[2]
+ scanchain_35/module_data_out[3] scanchain_35/module_data_out[4] scanchain_35/module_data_out[5]
+ scanchain_35/module_data_out[6] scanchain_35/module_data_out[7] vccd1 vssd1 rolfmobile99_alu_fsm_top
Xscanchain_45 scanchain_45/clk_in scanchain_46/clk_in scanchain_45/data_in scanchain_46/data_in
+ scanchain_45/latch_enable_in scanchain_46/latch_enable_in scanchain_45/module_data_in[0]
+ scanchain_45/module_data_in[1] scanchain_45/module_data_in[2] scanchain_45/module_data_in[3]
+ scanchain_45/module_data_in[4] scanchain_45/module_data_in[5] scanchain_45/module_data_in[6]
+ scanchain_45/module_data_in[7] scanchain_45/module_data_out[0] scanchain_45/module_data_out[1]
+ scanchain_45/module_data_out[2] scanchain_45/module_data_out[3] scanchain_45/module_data_out[4]
+ scanchain_45/module_data_out[5] scanchain_45/module_data_out[6] scanchain_45/module_data_out[7]
+ scanchain_45/scan_select_in scanchain_46/scan_select_in vccd1 vssd1 scanchain
Xscanchain_23 scanchain_23/clk_in scanchain_24/clk_in scanchain_23/data_in scanchain_24/data_in
+ scanchain_23/latch_enable_in scanchain_24/latch_enable_in scanchain_23/module_data_in[0]
+ scanchain_23/module_data_in[1] scanchain_23/module_data_in[2] scanchain_23/module_data_in[3]
+ scanchain_23/module_data_in[4] scanchain_23/module_data_in[5] scanchain_23/module_data_in[6]
+ scanchain_23/module_data_in[7] scanchain_23/module_data_out[0] scanchain_23/module_data_out[1]
+ scanchain_23/module_data_out[2] scanchain_23/module_data_out[3] scanchain_23/module_data_out[4]
+ scanchain_23/module_data_out[5] scanchain_23/module_data_out[6] scanchain_23/module_data_out[7]
+ scanchain_23/scan_select_in scanchain_24/scan_select_in vccd1 vssd1 scanchain
Xscanchain_34 scanchain_34/clk_in scanchain_35/clk_in scanchain_34/data_in scanchain_35/data_in
+ scanchain_34/latch_enable_in scanchain_35/latch_enable_in scanchain_34/module_data_in[0]
+ scanchain_34/module_data_in[1] scanchain_34/module_data_in[2] scanchain_34/module_data_in[3]
+ scanchain_34/module_data_in[4] scanchain_34/module_data_in[5] scanchain_34/module_data_in[6]
+ scanchain_34/module_data_in[7] scanchain_34/module_data_out[0] scanchain_34/module_data_out[1]
+ scanchain_34/module_data_out[2] scanchain_34/module_data_out[3] scanchain_34/module_data_out[4]
+ scanchain_34/module_data_out[5] scanchain_34/module_data_out[6] scanchain_34/module_data_out[7]
+ scanchain_34/scan_select_in scanchain_35/scan_select_in vccd1 vssd1 scanchain
Xscanchain_12 scanchain_12/clk_in scanchain_13/clk_in scanchain_12/data_in scanchain_13/data_in
+ scanchain_12/latch_enable_in scanchain_13/latch_enable_in scanchain_12/module_data_in[0]
+ scanchain_12/module_data_in[1] scanchain_12/module_data_in[2] scanchain_12/module_data_in[3]
+ scanchain_12/module_data_in[4] scanchain_12/module_data_in[5] scanchain_12/module_data_in[6]
+ scanchain_12/module_data_in[7] scanchain_12/module_data_out[0] scanchain_12/module_data_out[1]
+ scanchain_12/module_data_out[2] scanchain_12/module_data_out[3] scanchain_12/module_data_out[4]
+ scanchain_12/module_data_out[5] scanchain_12/module_data_out[6] scanchain_12/module_data_out[7]
+ scanchain_12/scan_select_in scanchain_13/scan_select_in vccd1 vssd1 scanchain
Xscanchain_67 scanchain_67/clk_in scanchain_68/clk_in scanchain_67/data_in scanchain_68/data_in
+ scanchain_67/latch_enable_in scanchain_68/latch_enable_in scanchain_67/module_data_in[0]
+ scanchain_67/module_data_in[1] scanchain_67/module_data_in[2] scanchain_67/module_data_in[3]
+ scanchain_67/module_data_in[4] scanchain_67/module_data_in[5] scanchain_67/module_data_in[6]
+ scanchain_67/module_data_in[7] scanchain_67/module_data_out[0] scanchain_67/module_data_out[1]
+ scanchain_67/module_data_out[2] scanchain_67/module_data_out[3] scanchain_67/module_data_out[4]
+ scanchain_67/module_data_out[5] scanchain_67/module_data_out[6] scanchain_67/module_data_out[7]
+ scanchain_67/scan_select_in scanchain_68/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_63 scanchain_63/module_data_in[0] scanchain_63/module_data_in[1]
+ scanchain_63/module_data_in[2] scanchain_63/module_data_in[3] scanchain_63/module_data_in[4]
+ scanchain_63/module_data_in[5] scanchain_63/module_data_in[6] scanchain_63/module_data_in[7]
+ scanchain_63/module_data_out[0] scanchain_63/module_data_out[1] scanchain_63/module_data_out[2]
+ scanchain_63/module_data_out[3] scanchain_63/module_data_out[4] scanchain_63/module_data_out[5]
+ scanchain_63/module_data_out[6] scanchain_63/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_56 scanchain_56/clk_in scanchain_57/clk_in scanchain_56/data_in scanchain_57/data_in
+ scanchain_56/latch_enable_in scanchain_57/latch_enable_in scanchain_56/module_data_in[0]
+ scanchain_56/module_data_in[1] scanchain_56/module_data_in[2] scanchain_56/module_data_in[3]
+ scanchain_56/module_data_in[4] scanchain_56/module_data_in[5] scanchain_56/module_data_in[6]
+ scanchain_56/module_data_in[7] scanchain_56/module_data_out[0] scanchain_56/module_data_out[1]
+ scanchain_56/module_data_out[2] scanchain_56/module_data_out[3] scanchain_56/module_data_out[4]
+ scanchain_56/module_data_out[5] scanchain_56/module_data_out[6] scanchain_56/module_data_out[7]
+ scanchain_56/scan_select_in scanchain_57/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_74 scanchain_74/module_data_in[0] scanchain_74/module_data_in[1]
+ scanchain_74/module_data_in[2] scanchain_74/module_data_in[3] scanchain_74/module_data_in[4]
+ scanchain_74/module_data_in[5] scanchain_74/module_data_in[6] scanchain_74/module_data_in[7]
+ scanchain_74/module_data_out[0] scanchain_74/module_data_out[1] scanchain_74/module_data_out[2]
+ scanchain_74/module_data_out[3] scanchain_74/module_data_out[4] scanchain_74/module_data_out[5]
+ scanchain_74/module_data_out[6] scanchain_74/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_78 scanchain_78/clk_in scanchain_79/clk_in scanchain_78/data_in scanchain_79/data_in
+ scanchain_78/latch_enable_in scanchain_79/latch_enable_in scanchain_78/module_data_in[0]
+ scanchain_78/module_data_in[1] scanchain_78/module_data_in[2] scanchain_78/module_data_in[3]
+ scanchain_78/module_data_in[4] scanchain_78/module_data_in[5] scanchain_78/module_data_in[6]
+ scanchain_78/module_data_in[7] scanchain_78/module_data_out[0] scanchain_78/module_data_out[1]
+ scanchain_78/module_data_out[2] scanchain_78/module_data_out[3] scanchain_78/module_data_out[4]
+ scanchain_78/module_data_out[5] scanchain_78/module_data_out[6] scanchain_78/module_data_out[7]
+ scanchain_78/scan_select_in scanchain_79/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_85 scanchain_85/module_data_in[0] scanchain_85/module_data_in[1]
+ scanchain_85/module_data_in[2] scanchain_85/module_data_in[3] scanchain_85/module_data_in[4]
+ scanchain_85/module_data_in[5] scanchain_85/module_data_in[6] scanchain_85/module_data_in[7]
+ scanchain_85/module_data_out[0] scanchain_85/module_data_out[1] scanchain_85/module_data_out[2]
+ scanchain_85/module_data_out[3] scanchain_85/module_data_out[4] scanchain_85/module_data_out[5]
+ scanchain_85/module_data_out[6] scanchain_85/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_89 scanchain_89/clk_in scanchain_90/clk_in scanchain_89/data_in scanchain_90/data_in
+ scanchain_89/latch_enable_in scanchain_90/latch_enable_in scanchain_89/module_data_in[0]
+ scanchain_89/module_data_in[1] scanchain_89/module_data_in[2] scanchain_89/module_data_in[3]
+ scanchain_89/module_data_in[4] scanchain_89/module_data_in[5] scanchain_89/module_data_in[6]
+ scanchain_89/module_data_in[7] scanchain_89/module_data_out[0] scanchain_89/module_data_out[1]
+ scanchain_89/module_data_out[2] scanchain_89/module_data_out[3] scanchain_89/module_data_out[4]
+ scanchain_89/module_data_out[5] scanchain_89/module_data_out[6] scanchain_89/module_data_out[7]
+ scanchain_89/scan_select_in scanchain_90/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_96 scanchain_96/module_data_in[0] scanchain_96/module_data_in[1]
+ scanchain_96/module_data_in[2] scanchain_96/module_data_in[3] scanchain_96/module_data_in[4]
+ scanchain_96/module_data_in[5] scanchain_96/module_data_in[6] scanchain_96/module_data_in[7]
+ scanchain_96/module_data_out[0] scanchain_96/module_data_out[1] scanchain_96/module_data_out[2]
+ scanchain_96/module_data_out[3] scanchain_96/module_data_out[4] scanchain_96/module_data_out[5]
+ scanchain_96/module_data_out[6] scanchain_96/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_390 scanchain_390/clk_in scanchain_391/clk_in scanchain_390/data_in scanchain_391/data_in
+ scanchain_390/latch_enable_in scanchain_391/latch_enable_in scanchain_390/module_data_in[0]
+ scanchain_390/module_data_in[1] scanchain_390/module_data_in[2] scanchain_390/module_data_in[3]
+ scanchain_390/module_data_in[4] scanchain_390/module_data_in[5] scanchain_390/module_data_in[6]
+ scanchain_390/module_data_in[7] scanchain_390/module_data_out[0] scanchain_390/module_data_out[1]
+ scanchain_390/module_data_out[2] scanchain_390/module_data_out[3] scanchain_390/module_data_out[4]
+ scanchain_390/module_data_out[5] scanchain_390/module_data_out[6] scanchain_390/module_data_out[7]
+ scanchain_390/scan_select_in scanchain_391/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341614374571475540_44 scanchain_44/module_data_in[0] scanchain_44/module_data_in[1]
+ scanchain_44/module_data_in[2] scanchain_44/module_data_in[3] scanchain_44/module_data_in[4]
+ scanchain_44/module_data_in[5] scanchain_44/module_data_in[6] scanchain_44/module_data_in[7]
+ scanchain_44/module_data_out[0] scanchain_44/module_data_out[1] scanchain_44/module_data_out[2]
+ scanchain_44/module_data_out[3] scanchain_44/module_data_out[4] scanchain_44/module_data_out[5]
+ scanchain_44/module_data_out[6] scanchain_44/module_data_out[7] vccd1 vssd1 user_module_341614374571475540
Xuser_module_339501025136214612_469 scanchain_469/module_data_in[0] scanchain_469/module_data_in[1]
+ scanchain_469/module_data_in[2] scanchain_469/module_data_in[3] scanchain_469/module_data_in[4]
+ scanchain_469/module_data_in[5] scanchain_469/module_data_in[6] scanchain_469/module_data_in[7]
+ scanchain_469/module_data_out[0] scanchain_469/module_data_out[1] scanchain_469/module_data_out[2]
+ scanchain_469/module_data_out[3] scanchain_469/module_data_out[4] scanchain_469/module_data_out[5]
+ scanchain_469/module_data_out[6] scanchain_469/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_458 scanchain_458/module_data_in[0] scanchain_458/module_data_in[1]
+ scanchain_458/module_data_in[2] scanchain_458/module_data_in[3] scanchain_458/module_data_in[4]
+ scanchain_458/module_data_in[5] scanchain_458/module_data_in[6] scanchain_458/module_data_in[7]
+ scanchain_458/module_data_out[0] scanchain_458/module_data_out[1] scanchain_458/module_data_out[2]
+ scanchain_458/module_data_out[3] scanchain_458/module_data_out[4] scanchain_458/module_data_out[5]
+ scanchain_458/module_data_out[6] scanchain_458/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_436 scanchain_436/module_data_in[0] scanchain_436/module_data_in[1]
+ scanchain_436/module_data_in[2] scanchain_436/module_data_in[3] scanchain_436/module_data_in[4]
+ scanchain_436/module_data_in[5] scanchain_436/module_data_in[6] scanchain_436/module_data_in[7]
+ scanchain_436/module_data_out[0] scanchain_436/module_data_out[1] scanchain_436/module_data_out[2]
+ scanchain_436/module_data_out[3] scanchain_436/module_data_out[4] scanchain_436/module_data_out[5]
+ scanchain_436/module_data_out[6] scanchain_436/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_447 scanchain_447/module_data_in[0] scanchain_447/module_data_in[1]
+ scanchain_447/module_data_in[2] scanchain_447/module_data_in[3] scanchain_447/module_data_in[4]
+ scanchain_447/module_data_in[5] scanchain_447/module_data_in[6] scanchain_447/module_data_in[7]
+ scanchain_447/module_data_out[0] scanchain_447/module_data_out[1] scanchain_447/module_data_out[2]
+ scanchain_447/module_data_out[3] scanchain_447/module_data_out[4] scanchain_447/module_data_out[5]
+ scanchain_447/module_data_out[6] scanchain_447/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_425 scanchain_425/module_data_in[0] scanchain_425/module_data_in[1]
+ scanchain_425/module_data_in[2] scanchain_425/module_data_in[3] scanchain_425/module_data_in[4]
+ scanchain_425/module_data_in[5] scanchain_425/module_data_in[6] scanchain_425/module_data_in[7]
+ scanchain_425/module_data_out[0] scanchain_425/module_data_out[1] scanchain_425/module_data_out[2]
+ scanchain_425/module_data_out[3] scanchain_425/module_data_out[4] scanchain_425/module_data_out[5]
+ scanchain_425/module_data_out[6] scanchain_425/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_403 scanchain_403/module_data_in[0] scanchain_403/module_data_in[1]
+ scanchain_403/module_data_in[2] scanchain_403/module_data_in[3] scanchain_403/module_data_in[4]
+ scanchain_403/module_data_in[5] scanchain_403/module_data_in[6] scanchain_403/module_data_in[7]
+ scanchain_403/module_data_out[0] scanchain_403/module_data_out[1] scanchain_403/module_data_out[2]
+ scanchain_403/module_data_out[3] scanchain_403/module_data_out[4] scanchain_403/module_data_out[5]
+ scanchain_403/module_data_out[6] scanchain_403/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_414 scanchain_414/module_data_in[0] scanchain_414/module_data_in[1]
+ scanchain_414/module_data_in[2] scanchain_414/module_data_in[3] scanchain_414/module_data_in[4]
+ scanchain_414/module_data_in[5] scanchain_414/module_data_in[6] scanchain_414/module_data_in[7]
+ scanchain_414/module_data_out[0] scanchain_414/module_data_out[1] scanchain_414/module_data_out[2]
+ scanchain_414/module_data_out[3] scanchain_414/module_data_out[4] scanchain_414/module_data_out[5]
+ scanchain_414/module_data_out[6] scanchain_414/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_288 scanchain_288/module_data_in[0] scanchain_288/module_data_in[1]
+ scanchain_288/module_data_in[2] scanchain_288/module_data_in[3] scanchain_288/module_data_in[4]
+ scanchain_288/module_data_in[5] scanchain_288/module_data_in[6] scanchain_288/module_data_in[7]
+ scanchain_288/module_data_out[0] scanchain_288/module_data_out[1] scanchain_288/module_data_out[2]
+ scanchain_288/module_data_out[3] scanchain_288/module_data_out[4] scanchain_288/module_data_out[5]
+ scanchain_288/module_data_out[6] scanchain_288/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_299 scanchain_299/module_data_in[0] scanchain_299/module_data_in[1]
+ scanchain_299/module_data_in[2] scanchain_299/module_data_in[3] scanchain_299/module_data_in[4]
+ scanchain_299/module_data_in[5] scanchain_299/module_data_in[6] scanchain_299/module_data_in[7]
+ scanchain_299/module_data_out[0] scanchain_299/module_data_out[1] scanchain_299/module_data_out[2]
+ scanchain_299/module_data_out[3] scanchain_299/module_data_out[4] scanchain_299/module_data_out[5]
+ scanchain_299/module_data_out[6] scanchain_299/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_277 scanchain_277/module_data_in[0] scanchain_277/module_data_in[1]
+ scanchain_277/module_data_in[2] scanchain_277/module_data_in[3] scanchain_277/module_data_in[4]
+ scanchain_277/module_data_in[5] scanchain_277/module_data_in[6] scanchain_277/module_data_in[7]
+ scanchain_277/module_data_out[0] scanchain_277/module_data_out[1] scanchain_277/module_data_out[2]
+ scanchain_277/module_data_out[3] scanchain_277/module_data_out[4] scanchain_277/module_data_out[5]
+ scanchain_277/module_data_out[6] scanchain_277/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_266 scanchain_266/module_data_in[0] scanchain_266/module_data_in[1]
+ scanchain_266/module_data_in[2] scanchain_266/module_data_in[3] scanchain_266/module_data_in[4]
+ scanchain_266/module_data_in[5] scanchain_266/module_data_in[6] scanchain_266/module_data_in[7]
+ scanchain_266/module_data_out[0] scanchain_266/module_data_out[1] scanchain_266/module_data_out[2]
+ scanchain_266/module_data_out[3] scanchain_266/module_data_out[4] scanchain_266/module_data_out[5]
+ scanchain_266/module_data_out[6] scanchain_266/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_255 scanchain_255/module_data_in[0] scanchain_255/module_data_in[1]
+ scanchain_255/module_data_in[2] scanchain_255/module_data_in[3] scanchain_255/module_data_in[4]
+ scanchain_255/module_data_in[5] scanchain_255/module_data_in[6] scanchain_255/module_data_in[7]
+ scanchain_255/module_data_out[0] scanchain_255/module_data_out[1] scanchain_255/module_data_out[2]
+ scanchain_255/module_data_out[3] scanchain_255/module_data_out[4] scanchain_255/module_data_out[5]
+ scanchain_255/module_data_out[6] scanchain_255/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_244 scanchain_244/module_data_in[0] scanchain_244/module_data_in[1]
+ scanchain_244/module_data_in[2] scanchain_244/module_data_in[3] scanchain_244/module_data_in[4]
+ scanchain_244/module_data_in[5] scanchain_244/module_data_in[6] scanchain_244/module_data_in[7]
+ scanchain_244/module_data_out[0] scanchain_244/module_data_out[1] scanchain_244/module_data_out[2]
+ scanchain_244/module_data_out[3] scanchain_244/module_data_out[4] scanchain_244/module_data_out[5]
+ scanchain_244/module_data_out[6] scanchain_244/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_233 scanchain_233/module_data_in[0] scanchain_233/module_data_in[1]
+ scanchain_233/module_data_in[2] scanchain_233/module_data_in[3] scanchain_233/module_data_in[4]
+ scanchain_233/module_data_in[5] scanchain_233/module_data_in[6] scanchain_233/module_data_in[7]
+ scanchain_233/module_data_out[0] scanchain_233/module_data_out[1] scanchain_233/module_data_out[2]
+ scanchain_233/module_data_out[3] scanchain_233/module_data_out[4] scanchain_233/module_data_out[5]
+ scanchain_233/module_data_out[6] scanchain_233/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_208 scanchain_208/clk_in scanchain_209/clk_in scanchain_208/data_in scanchain_209/data_in
+ scanchain_208/latch_enable_in scanchain_209/latch_enable_in scanchain_208/module_data_in[0]
+ scanchain_208/module_data_in[1] scanchain_208/module_data_in[2] scanchain_208/module_data_in[3]
+ scanchain_208/module_data_in[4] scanchain_208/module_data_in[5] scanchain_208/module_data_in[6]
+ scanchain_208/module_data_in[7] scanchain_208/module_data_out[0] scanchain_208/module_data_out[1]
+ scanchain_208/module_data_out[2] scanchain_208/module_data_out[3] scanchain_208/module_data_out[4]
+ scanchain_208/module_data_out[5] scanchain_208/module_data_out[6] scanchain_208/module_data_out[7]
+ scanchain_208/scan_select_in scanchain_209/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_211 scanchain_211/module_data_in[0] scanchain_211/module_data_in[1]
+ scanchain_211/module_data_in[2] scanchain_211/module_data_in[3] scanchain_211/module_data_in[4]
+ scanchain_211/module_data_in[5] scanchain_211/module_data_in[6] scanchain_211/module_data_in[7]
+ scanchain_211/module_data_out[0] scanchain_211/module_data_out[1] scanchain_211/module_data_out[2]
+ scanchain_211/module_data_out[3] scanchain_211/module_data_out[4] scanchain_211/module_data_out[5]
+ scanchain_211/module_data_out[6] scanchain_211/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_219 scanchain_219/clk_in scanchain_220/clk_in scanchain_219/data_in scanchain_220/data_in
+ scanchain_219/latch_enable_in scanchain_220/latch_enable_in scanchain_219/module_data_in[0]
+ scanchain_219/module_data_in[1] scanchain_219/module_data_in[2] scanchain_219/module_data_in[3]
+ scanchain_219/module_data_in[4] scanchain_219/module_data_in[5] scanchain_219/module_data_in[6]
+ scanchain_219/module_data_in[7] scanchain_219/module_data_out[0] scanchain_219/module_data_out[1]
+ scanchain_219/module_data_out[2] scanchain_219/module_data_out[3] scanchain_219/module_data_out[4]
+ scanchain_219/module_data_out[5] scanchain_219/module_data_out[6] scanchain_219/module_data_out[7]
+ scanchain_219/scan_select_in scanchain_220/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_222 scanchain_222/module_data_in[0] scanchain_222/module_data_in[1]
+ scanchain_222/module_data_in[2] scanchain_222/module_data_in[3] scanchain_222/module_data_in[4]
+ scanchain_222/module_data_in[5] scanchain_222/module_data_in[6] scanchain_222/module_data_in[7]
+ scanchain_222/module_data_out[0] scanchain_222/module_data_out[1] scanchain_222/module_data_out[2]
+ scanchain_222/module_data_out[3] scanchain_222/module_data_out[4] scanchain_222/module_data_out[5]
+ scanchain_222/module_data_out[6] scanchain_222/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_200 scanchain_200/module_data_in[0] scanchain_200/module_data_in[1]
+ scanchain_200/module_data_in[2] scanchain_200/module_data_in[3] scanchain_200/module_data_in[4]
+ scanchain_200/module_data_in[5] scanchain_200/module_data_in[6] scanchain_200/module_data_in[7]
+ scanchain_200/module_data_out[0] scanchain_200/module_data_out[1] scanchain_200/module_data_out[2]
+ scanchain_200/module_data_out[3] scanchain_200/module_data_out[4] scanchain_200/module_data_out[5]
+ scanchain_200/module_data_out[6] scanchain_200/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_46 scanchain_46/clk_in scanchain_47/clk_in scanchain_46/data_in scanchain_47/data_in
+ scanchain_46/latch_enable_in scanchain_47/latch_enable_in scanchain_46/module_data_in[0]
+ scanchain_46/module_data_in[1] scanchain_46/module_data_in[2] scanchain_46/module_data_in[3]
+ scanchain_46/module_data_in[4] scanchain_46/module_data_in[5] scanchain_46/module_data_in[6]
+ scanchain_46/module_data_in[7] scanchain_46/module_data_out[0] scanchain_46/module_data_out[1]
+ scanchain_46/module_data_out[2] scanchain_46/module_data_out[3] scanchain_46/module_data_out[4]
+ scanchain_46/module_data_out[5] scanchain_46/module_data_out[6] scanchain_46/module_data_out[7]
+ scanchain_46/scan_select_in scanchain_47/scan_select_in vccd1 vssd1 scanchain
Xscanchain_24 scanchain_24/clk_in scanchain_25/clk_in scanchain_24/data_in scanchain_25/data_in
+ scanchain_24/latch_enable_in scanchain_25/latch_enable_in scanchain_24/module_data_in[0]
+ scanchain_24/module_data_in[1] scanchain_24/module_data_in[2] scanchain_24/module_data_in[3]
+ scanchain_24/module_data_in[4] scanchain_24/module_data_in[5] scanchain_24/module_data_in[6]
+ scanchain_24/module_data_in[7] scanchain_24/module_data_out[0] scanchain_24/module_data_out[1]
+ scanchain_24/module_data_out[2] scanchain_24/module_data_out[3] scanchain_24/module_data_out[4]
+ scanchain_24/module_data_out[5] scanchain_24/module_data_out[6] scanchain_24/module_data_out[7]
+ scanchain_24/scan_select_in scanchain_25/scan_select_in vccd1 vssd1 scanchain
Xscanchain_35 scanchain_35/clk_in scanchain_36/clk_in scanchain_35/data_in scanchain_36/data_in
+ scanchain_35/latch_enable_in scanchain_36/latch_enable_in scanchain_35/module_data_in[0]
+ scanchain_35/module_data_in[1] scanchain_35/module_data_in[2] scanchain_35/module_data_in[3]
+ scanchain_35/module_data_in[4] scanchain_35/module_data_in[5] scanchain_35/module_data_in[6]
+ scanchain_35/module_data_in[7] scanchain_35/module_data_out[0] scanchain_35/module_data_out[1]
+ scanchain_35/module_data_out[2] scanchain_35/module_data_out[3] scanchain_35/module_data_out[4]
+ scanchain_35/module_data_out[5] scanchain_35/module_data_out[6] scanchain_35/module_data_out[7]
+ scanchain_35/scan_select_in scanchain_36/scan_select_in vccd1 vssd1 scanchain
Xscanchain_13 scanchain_13/clk_in scanchain_14/clk_in scanchain_13/data_in scanchain_14/data_in
+ scanchain_13/latch_enable_in scanchain_14/latch_enable_in scanchain_13/module_data_in[0]
+ scanchain_13/module_data_in[1] scanchain_13/module_data_in[2] scanchain_13/module_data_in[3]
+ scanchain_13/module_data_in[4] scanchain_13/module_data_in[5] scanchain_13/module_data_in[6]
+ scanchain_13/module_data_in[7] scanchain_13/module_data_out[0] scanchain_13/module_data_out[1]
+ scanchain_13/module_data_out[2] scanchain_13/module_data_out[3] scanchain_13/module_data_out[4]
+ scanchain_13/module_data_out[5] scanchain_13/module_data_out[6] scanchain_13/module_data_out[7]
+ scanchain_13/scan_select_in scanchain_14/scan_select_in vccd1 vssd1 scanchain
Xscanchain_68 scanchain_68/clk_in scanchain_69/clk_in scanchain_68/data_in scanchain_69/data_in
+ scanchain_68/latch_enable_in scanchain_69/latch_enable_in scanchain_68/module_data_in[0]
+ scanchain_68/module_data_in[1] scanchain_68/module_data_in[2] scanchain_68/module_data_in[3]
+ scanchain_68/module_data_in[4] scanchain_68/module_data_in[5] scanchain_68/module_data_in[6]
+ scanchain_68/module_data_in[7] scanchain_68/module_data_out[0] scanchain_68/module_data_out[1]
+ scanchain_68/module_data_out[2] scanchain_68/module_data_out[3] scanchain_68/module_data_out[4]
+ scanchain_68/module_data_out[5] scanchain_68/module_data_out[6] scanchain_68/module_data_out[7]
+ scanchain_68/scan_select_in scanchain_69/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_64 scanchain_64/module_data_in[0] scanchain_64/module_data_in[1]
+ scanchain_64/module_data_in[2] scanchain_64/module_data_in[3] scanchain_64/module_data_in[4]
+ scanchain_64/module_data_in[5] scanchain_64/module_data_in[6] scanchain_64/module_data_in[7]
+ scanchain_64/module_data_out[0] scanchain_64/module_data_out[1] scanchain_64/module_data_out[2]
+ scanchain_64/module_data_out[3] scanchain_64/module_data_out[4] scanchain_64/module_data_out[5]
+ scanchain_64/module_data_out[6] scanchain_64/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_57 scanchain_57/clk_in scanchain_58/clk_in scanchain_57/data_in scanchain_58/data_in
+ scanchain_57/latch_enable_in scanchain_58/latch_enable_in scanchain_57/module_data_in[0]
+ scanchain_57/module_data_in[1] scanchain_57/module_data_in[2] scanchain_57/module_data_in[3]
+ scanchain_57/module_data_in[4] scanchain_57/module_data_in[5] scanchain_57/module_data_in[6]
+ scanchain_57/module_data_in[7] scanchain_57/module_data_out[0] scanchain_57/module_data_out[1]
+ scanchain_57/module_data_out[2] scanchain_57/module_data_out[3] scanchain_57/module_data_out[4]
+ scanchain_57/module_data_out[5] scanchain_57/module_data_out[6] scanchain_57/module_data_out[7]
+ scanchain_57/scan_select_in scanchain_58/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_75 scanchain_75/module_data_in[0] scanchain_75/module_data_in[1]
+ scanchain_75/module_data_in[2] scanchain_75/module_data_in[3] scanchain_75/module_data_in[4]
+ scanchain_75/module_data_in[5] scanchain_75/module_data_in[6] scanchain_75/module_data_in[7]
+ scanchain_75/module_data_out[0] scanchain_75/module_data_out[1] scanchain_75/module_data_out[2]
+ scanchain_75/module_data_out[3] scanchain_75/module_data_out[4] scanchain_75/module_data_out[5]
+ scanchain_75/module_data_out[6] scanchain_75/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_86 scanchain_86/module_data_in[0] scanchain_86/module_data_in[1]
+ scanchain_86/module_data_in[2] scanchain_86/module_data_in[3] scanchain_86/module_data_in[4]
+ scanchain_86/module_data_in[5] scanchain_86/module_data_in[6] scanchain_86/module_data_in[7]
+ scanchain_86/module_data_out[0] scanchain_86/module_data_out[1] scanchain_86/module_data_out[2]
+ scanchain_86/module_data_out[3] scanchain_86/module_data_out[4] scanchain_86/module_data_out[5]
+ scanchain_86/module_data_out[6] scanchain_86/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_97 scanchain_97/module_data_in[0] scanchain_97/module_data_in[1]
+ scanchain_97/module_data_in[2] scanchain_97/module_data_in[3] scanchain_97/module_data_in[4]
+ scanchain_97/module_data_in[5] scanchain_97/module_data_in[6] scanchain_97/module_data_in[7]
+ scanchain_97/module_data_out[0] scanchain_97/module_data_out[1] scanchain_97/module_data_out[2]
+ scanchain_97/module_data_out[3] scanchain_97/module_data_out[4] scanchain_97/module_data_out[5]
+ scanchain_97/module_data_out[6] scanchain_97/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_391 scanchain_391/clk_in scanchain_392/clk_in scanchain_391/data_in scanchain_392/data_in
+ scanchain_391/latch_enable_in scanchain_392/latch_enable_in scanchain_391/module_data_in[0]
+ scanchain_391/module_data_in[1] scanchain_391/module_data_in[2] scanchain_391/module_data_in[3]
+ scanchain_391/module_data_in[4] scanchain_391/module_data_in[5] scanchain_391/module_data_in[6]
+ scanchain_391/module_data_in[7] scanchain_391/module_data_out[0] scanchain_391/module_data_out[1]
+ scanchain_391/module_data_out[2] scanchain_391/module_data_out[3] scanchain_391/module_data_out[4]
+ scanchain_391/module_data_out[5] scanchain_391/module_data_out[6] scanchain_391/module_data_out[7]
+ scanchain_391/scan_select_in scanchain_392/scan_select_in vccd1 vssd1 scanchain
Xscanchain_380 scanchain_380/clk_in scanchain_381/clk_in scanchain_380/data_in scanchain_381/data_in
+ scanchain_380/latch_enable_in scanchain_381/latch_enable_in scanchain_380/module_data_in[0]
+ scanchain_380/module_data_in[1] scanchain_380/module_data_in[2] scanchain_380/module_data_in[3]
+ scanchain_380/module_data_in[4] scanchain_380/module_data_in[5] scanchain_380/module_data_in[6]
+ scanchain_380/module_data_in[7] scanchain_380/module_data_out[0] scanchain_380/module_data_out[1]
+ scanchain_380/module_data_out[2] scanchain_380/module_data_out[3] scanchain_380/module_data_out[4]
+ scanchain_380/module_data_out[5] scanchain_380/module_data_out[6] scanchain_380/module_data_out[7]
+ scanchain_380/scan_select_in scanchain_381/scan_select_in vccd1 vssd1 scanchain
Xscanchain_79 scanchain_79/clk_in scanchain_80/clk_in scanchain_79/data_in scanchain_80/data_in
+ scanchain_79/latch_enable_in scanchain_80/latch_enable_in scanchain_79/module_data_in[0]
+ scanchain_79/module_data_in[1] scanchain_79/module_data_in[2] scanchain_79/module_data_in[3]
+ scanchain_79/module_data_in[4] scanchain_79/module_data_in[5] scanchain_79/module_data_in[6]
+ scanchain_79/module_data_in[7] scanchain_79/module_data_out[0] scanchain_79/module_data_out[1]
+ scanchain_79/module_data_out[2] scanchain_79/module_data_out[3] scanchain_79/module_data_out[4]
+ scanchain_79/module_data_out[5] scanchain_79/module_data_out[6] scanchain_79/module_data_out[7]
+ scanchain_79/scan_select_in scanchain_80/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_459 scanchain_459/module_data_in[0] scanchain_459/module_data_in[1]
+ scanchain_459/module_data_in[2] scanchain_459/module_data_in[3] scanchain_459/module_data_in[4]
+ scanchain_459/module_data_in[5] scanchain_459/module_data_in[6] scanchain_459/module_data_in[7]
+ scanchain_459/module_data_out[0] scanchain_459/module_data_out[1] scanchain_459/module_data_out[2]
+ scanchain_459/module_data_out[3] scanchain_459/module_data_out[4] scanchain_459/module_data_out[5]
+ scanchain_459/module_data_out[6] scanchain_459/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_437 scanchain_437/module_data_in[0] scanchain_437/module_data_in[1]
+ scanchain_437/module_data_in[2] scanchain_437/module_data_in[3] scanchain_437/module_data_in[4]
+ scanchain_437/module_data_in[5] scanchain_437/module_data_in[6] scanchain_437/module_data_in[7]
+ scanchain_437/module_data_out[0] scanchain_437/module_data_out[1] scanchain_437/module_data_out[2]
+ scanchain_437/module_data_out[3] scanchain_437/module_data_out[4] scanchain_437/module_data_out[5]
+ scanchain_437/module_data_out[6] scanchain_437/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_448 scanchain_448/module_data_in[0] scanchain_448/module_data_in[1]
+ scanchain_448/module_data_in[2] scanchain_448/module_data_in[3] scanchain_448/module_data_in[4]
+ scanchain_448/module_data_in[5] scanchain_448/module_data_in[6] scanchain_448/module_data_in[7]
+ scanchain_448/module_data_out[0] scanchain_448/module_data_out[1] scanchain_448/module_data_out[2]
+ scanchain_448/module_data_out[3] scanchain_448/module_data_out[4] scanchain_448/module_data_out[5]
+ scanchain_448/module_data_out[6] scanchain_448/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_426 scanchain_426/module_data_in[0] scanchain_426/module_data_in[1]
+ scanchain_426/module_data_in[2] scanchain_426/module_data_in[3] scanchain_426/module_data_in[4]
+ scanchain_426/module_data_in[5] scanchain_426/module_data_in[6] scanchain_426/module_data_in[7]
+ scanchain_426/module_data_out[0] scanchain_426/module_data_out[1] scanchain_426/module_data_out[2]
+ scanchain_426/module_data_out[3] scanchain_426/module_data_out[4] scanchain_426/module_data_out[5]
+ scanchain_426/module_data_out[6] scanchain_426/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_404 scanchain_404/module_data_in[0] scanchain_404/module_data_in[1]
+ scanchain_404/module_data_in[2] scanchain_404/module_data_in[3] scanchain_404/module_data_in[4]
+ scanchain_404/module_data_in[5] scanchain_404/module_data_in[6] scanchain_404/module_data_in[7]
+ scanchain_404/module_data_out[0] scanchain_404/module_data_out[1] scanchain_404/module_data_out[2]
+ scanchain_404/module_data_out[3] scanchain_404/module_data_out[4] scanchain_404/module_data_out[5]
+ scanchain_404/module_data_out[6] scanchain_404/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_415 scanchain_415/module_data_in[0] scanchain_415/module_data_in[1]
+ scanchain_415/module_data_in[2] scanchain_415/module_data_in[3] scanchain_415/module_data_in[4]
+ scanchain_415/module_data_in[5] scanchain_415/module_data_in[6] scanchain_415/module_data_in[7]
+ scanchain_415/module_data_out[0] scanchain_415/module_data_out[1] scanchain_415/module_data_out[2]
+ scanchain_415/module_data_out[3] scanchain_415/module_data_out[4] scanchain_415/module_data_out[5]
+ scanchain_415/module_data_out[6] scanchain_415/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_289 scanchain_289/module_data_in[0] scanchain_289/module_data_in[1]
+ scanchain_289/module_data_in[2] scanchain_289/module_data_in[3] scanchain_289/module_data_in[4]
+ scanchain_289/module_data_in[5] scanchain_289/module_data_in[6] scanchain_289/module_data_in[7]
+ scanchain_289/module_data_out[0] scanchain_289/module_data_out[1] scanchain_289/module_data_out[2]
+ scanchain_289/module_data_out[3] scanchain_289/module_data_out[4] scanchain_289/module_data_out[5]
+ scanchain_289/module_data_out[6] scanchain_289/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_278 scanchain_278/module_data_in[0] scanchain_278/module_data_in[1]
+ scanchain_278/module_data_in[2] scanchain_278/module_data_in[3] scanchain_278/module_data_in[4]
+ scanchain_278/module_data_in[5] scanchain_278/module_data_in[6] scanchain_278/module_data_in[7]
+ scanchain_278/module_data_out[0] scanchain_278/module_data_out[1] scanchain_278/module_data_out[2]
+ scanchain_278/module_data_out[3] scanchain_278/module_data_out[4] scanchain_278/module_data_out[5]
+ scanchain_278/module_data_out[6] scanchain_278/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_267 scanchain_267/module_data_in[0] scanchain_267/module_data_in[1]
+ scanchain_267/module_data_in[2] scanchain_267/module_data_in[3] scanchain_267/module_data_in[4]
+ scanchain_267/module_data_in[5] scanchain_267/module_data_in[6] scanchain_267/module_data_in[7]
+ scanchain_267/module_data_out[0] scanchain_267/module_data_out[1] scanchain_267/module_data_out[2]
+ scanchain_267/module_data_out[3] scanchain_267/module_data_out[4] scanchain_267/module_data_out[5]
+ scanchain_267/module_data_out[6] scanchain_267/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_245 scanchain_245/module_data_in[0] scanchain_245/module_data_in[1]
+ scanchain_245/module_data_in[2] scanchain_245/module_data_in[3] scanchain_245/module_data_in[4]
+ scanchain_245/module_data_in[5] scanchain_245/module_data_in[6] scanchain_245/module_data_in[7]
+ scanchain_245/module_data_out[0] scanchain_245/module_data_out[1] scanchain_245/module_data_out[2]
+ scanchain_245/module_data_out[3] scanchain_245/module_data_out[4] scanchain_245/module_data_out[5]
+ scanchain_245/module_data_out[6] scanchain_245/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_256 scanchain_256/module_data_in[0] scanchain_256/module_data_in[1]
+ scanchain_256/module_data_in[2] scanchain_256/module_data_in[3] scanchain_256/module_data_in[4]
+ scanchain_256/module_data_in[5] scanchain_256/module_data_in[6] scanchain_256/module_data_in[7]
+ scanchain_256/module_data_out[0] scanchain_256/module_data_out[1] scanchain_256/module_data_out[2]
+ scanchain_256/module_data_out[3] scanchain_256/module_data_out[4] scanchain_256/module_data_out[5]
+ scanchain_256/module_data_out[6] scanchain_256/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_234 scanchain_234/module_data_in[0] scanchain_234/module_data_in[1]
+ scanchain_234/module_data_in[2] scanchain_234/module_data_in[3] scanchain_234/module_data_in[4]
+ scanchain_234/module_data_in[5] scanchain_234/module_data_in[6] scanchain_234/module_data_in[7]
+ scanchain_234/module_data_out[0] scanchain_234/module_data_out[1] scanchain_234/module_data_out[2]
+ scanchain_234/module_data_out[3] scanchain_234/module_data_out[4] scanchain_234/module_data_out[5]
+ scanchain_234/module_data_out[6] scanchain_234/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_212 scanchain_212/module_data_in[0] scanchain_212/module_data_in[1]
+ scanchain_212/module_data_in[2] scanchain_212/module_data_in[3] scanchain_212/module_data_in[4]
+ scanchain_212/module_data_in[5] scanchain_212/module_data_in[6] scanchain_212/module_data_in[7]
+ scanchain_212/module_data_out[0] scanchain_212/module_data_out[1] scanchain_212/module_data_out[2]
+ scanchain_212/module_data_out[3] scanchain_212/module_data_out[4] scanchain_212/module_data_out[5]
+ scanchain_212/module_data_out[6] scanchain_212/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_223 scanchain_223/module_data_in[0] scanchain_223/module_data_in[1]
+ scanchain_223/module_data_in[2] scanchain_223/module_data_in[3] scanchain_223/module_data_in[4]
+ scanchain_223/module_data_in[5] scanchain_223/module_data_in[6] scanchain_223/module_data_in[7]
+ scanchain_223/module_data_out[0] scanchain_223/module_data_out[1] scanchain_223/module_data_out[2]
+ scanchain_223/module_data_out[3] scanchain_223/module_data_out[4] scanchain_223/module_data_out[5]
+ scanchain_223/module_data_out[6] scanchain_223/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_201 scanchain_201/module_data_in[0] scanchain_201/module_data_in[1]
+ scanchain_201/module_data_in[2] scanchain_201/module_data_in[3] scanchain_201/module_data_in[4]
+ scanchain_201/module_data_in[5] scanchain_201/module_data_in[6] scanchain_201/module_data_in[7]
+ scanchain_201/module_data_out[0] scanchain_201/module_data_out[1] scanchain_201/module_data_out[2]
+ scanchain_201/module_data_out[3] scanchain_201/module_data_out[4] scanchain_201/module_data_out[5]
+ scanchain_201/module_data_out[6] scanchain_201/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_209 scanchain_209/clk_in scanchain_210/clk_in scanchain_209/data_in scanchain_210/data_in
+ scanchain_209/latch_enable_in scanchain_210/latch_enable_in scanchain_209/module_data_in[0]
+ scanchain_209/module_data_in[1] scanchain_209/module_data_in[2] scanchain_209/module_data_in[3]
+ scanchain_209/module_data_in[4] scanchain_209/module_data_in[5] scanchain_209/module_data_in[6]
+ scanchain_209/module_data_in[7] scanchain_209/module_data_out[0] scanchain_209/module_data_out[1]
+ scanchain_209/module_data_out[2] scanchain_209/module_data_out[3] scanchain_209/module_data_out[4]
+ scanchain_209/module_data_out[5] scanchain_209/module_data_out[6] scanchain_209/module_data_out[7]
+ scanchain_209/scan_select_in scanchain_210/scan_select_in vccd1 vssd1 scanchain
Xuser_module_347787021138264660_10 scanchain_10/module_data_in[0] scanchain_10/module_data_in[1]
+ scanchain_10/module_data_in[2] scanchain_10/module_data_in[3] scanchain_10/module_data_in[4]
+ scanchain_10/module_data_in[5] scanchain_10/module_data_in[6] scanchain_10/module_data_in[7]
+ scanchain_10/module_data_out[0] scanchain_10/module_data_out[1] scanchain_10/module_data_out[2]
+ scanchain_10/module_data_out[3] scanchain_10/module_data_out[4] scanchain_10/module_data_out[5]
+ scanchain_10/module_data_out[6] scanchain_10/module_data_out[7] vccd1 vssd1 user_module_347787021138264660
Xuser_module_339501025136214612_65 scanchain_65/module_data_in[0] scanchain_65/module_data_in[1]
+ scanchain_65/module_data_in[2] scanchain_65/module_data_in[3] scanchain_65/module_data_in[4]
+ scanchain_65/module_data_in[5] scanchain_65/module_data_in[6] scanchain_65/module_data_in[7]
+ scanchain_65/module_data_out[0] scanchain_65/module_data_out[1] scanchain_65/module_data_out[2]
+ scanchain_65/module_data_out[3] scanchain_65/module_data_out[4] scanchain_65/module_data_out[5]
+ scanchain_65/module_data_out[6] scanchain_65/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_76 scanchain_76/module_data_in[0] scanchain_76/module_data_in[1]
+ scanchain_76/module_data_in[2] scanchain_76/module_data_in[3] scanchain_76/module_data_in[4]
+ scanchain_76/module_data_in[5] scanchain_76/module_data_in[6] scanchain_76/module_data_in[7]
+ scanchain_76/module_data_out[0] scanchain_76/module_data_out[1] scanchain_76/module_data_out[2]
+ scanchain_76/module_data_out[3] scanchain_76/module_data_out[4] scanchain_76/module_data_out[5]
+ scanchain_76/module_data_out[6] scanchain_76/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_87 scanchain_87/module_data_in[0] scanchain_87/module_data_in[1]
+ scanchain_87/module_data_in[2] scanchain_87/module_data_in[3] scanchain_87/module_data_in[4]
+ scanchain_87/module_data_in[5] scanchain_87/module_data_in[6] scanchain_87/module_data_in[7]
+ scanchain_87/module_data_out[0] scanchain_87/module_data_out[1] scanchain_87/module_data_out[2]
+ scanchain_87/module_data_out[3] scanchain_87/module_data_out[4] scanchain_87/module_data_out[5]
+ scanchain_87/module_data_out[6] scanchain_87/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_98 scanchain_98/module_data_in[0] scanchain_98/module_data_in[1]
+ scanchain_98/module_data_in[2] scanchain_98/module_data_in[3] scanchain_98/module_data_in[4]
+ scanchain_98/module_data_in[5] scanchain_98/module_data_in[6] scanchain_98/module_data_in[7]
+ scanchain_98/module_data_out[0] scanchain_98/module_data_out[1] scanchain_98/module_data_out[2]
+ scanchain_98/module_data_out[3] scanchain_98/module_data_out[4] scanchain_98/module_data_out[5]
+ scanchain_98/module_data_out[6] scanchain_98/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_392 scanchain_392/clk_in scanchain_393/clk_in scanchain_392/data_in scanchain_393/data_in
+ scanchain_392/latch_enable_in scanchain_393/latch_enable_in scanchain_392/module_data_in[0]
+ scanchain_392/module_data_in[1] scanchain_392/module_data_in[2] scanchain_392/module_data_in[3]
+ scanchain_392/module_data_in[4] scanchain_392/module_data_in[5] scanchain_392/module_data_in[6]
+ scanchain_392/module_data_in[7] scanchain_392/module_data_out[0] scanchain_392/module_data_out[1]
+ scanchain_392/module_data_out[2] scanchain_392/module_data_out[3] scanchain_392/module_data_out[4]
+ scanchain_392/module_data_out[5] scanchain_392/module_data_out[6] scanchain_392/module_data_out[7]
+ scanchain_392/scan_select_in scanchain_393/scan_select_in vccd1 vssd1 scanchain
Xscanchain_381 scanchain_381/clk_in scanchain_382/clk_in scanchain_381/data_in scanchain_382/data_in
+ scanchain_381/latch_enable_in scanchain_382/latch_enable_in scanchain_381/module_data_in[0]
+ scanchain_381/module_data_in[1] scanchain_381/module_data_in[2] scanchain_381/module_data_in[3]
+ scanchain_381/module_data_in[4] scanchain_381/module_data_in[5] scanchain_381/module_data_in[6]
+ scanchain_381/module_data_in[7] scanchain_381/module_data_out[0] scanchain_381/module_data_out[1]
+ scanchain_381/module_data_out[2] scanchain_381/module_data_out[3] scanchain_381/module_data_out[4]
+ scanchain_381/module_data_out[5] scanchain_381/module_data_out[6] scanchain_381/module_data_out[7]
+ scanchain_381/scan_select_in scanchain_382/scan_select_in vccd1 vssd1 scanchain
Xscanchain_370 scanchain_370/clk_in scanchain_371/clk_in scanchain_370/data_in scanchain_371/data_in
+ scanchain_370/latch_enable_in scanchain_371/latch_enable_in scanchain_370/module_data_in[0]
+ scanchain_370/module_data_in[1] scanchain_370/module_data_in[2] scanchain_370/module_data_in[3]
+ scanchain_370/module_data_in[4] scanchain_370/module_data_in[5] scanchain_370/module_data_in[6]
+ scanchain_370/module_data_in[7] scanchain_370/module_data_out[0] scanchain_370/module_data_out[1]
+ scanchain_370/module_data_out[2] scanchain_370/module_data_out[3] scanchain_370/module_data_out[4]
+ scanchain_370/module_data_out[5] scanchain_370/module_data_out[6] scanchain_370/module_data_out[7]
+ scanchain_370/scan_select_in scanchain_371/scan_select_in vccd1 vssd1 scanchain
Xscanchain_47 scanchain_47/clk_in scanchain_48/clk_in scanchain_47/data_in scanchain_48/data_in
+ scanchain_47/latch_enable_in scanchain_48/latch_enable_in scanchain_47/module_data_in[0]
+ scanchain_47/module_data_in[1] scanchain_47/module_data_in[2] scanchain_47/module_data_in[3]
+ scanchain_47/module_data_in[4] scanchain_47/module_data_in[5] scanchain_47/module_data_in[6]
+ scanchain_47/module_data_in[7] scanchain_47/module_data_out[0] scanchain_47/module_data_out[1]
+ scanchain_47/module_data_out[2] scanchain_47/module_data_out[3] scanchain_47/module_data_out[4]
+ scanchain_47/module_data_out[5] scanchain_47/module_data_out[6] scanchain_47/module_data_out[7]
+ scanchain_47/scan_select_in scanchain_48/scan_select_in vccd1 vssd1 scanchain
Xscanchain_36 scanchain_36/clk_in scanchain_37/clk_in scanchain_36/data_in scanchain_37/data_in
+ scanchain_36/latch_enable_in scanchain_37/latch_enable_in jar_illegal_logic_36/io_in[0]
+ jar_illegal_logic_36/io_in[1] jar_illegal_logic_36/io_in[2] jar_illegal_logic_36/io_in[3]
+ jar_illegal_logic_36/io_in[4] jar_illegal_logic_36/io_in[5] jar_illegal_logic_36/io_in[6]
+ jar_illegal_logic_36/io_in[7] jar_illegal_logic_36/io_out[0] jar_illegal_logic_36/io_out[1]
+ jar_illegal_logic_36/io_out[2] jar_illegal_logic_36/io_out[3] jar_illegal_logic_36/io_out[4]
+ jar_illegal_logic_36/io_out[5] jar_illegal_logic_36/io_out[6] jar_illegal_logic_36/io_out[7]
+ scanchain_36/scan_select_in scanchain_37/scan_select_in vccd1 vssd1 scanchain
Xscanchain_25 scanchain_25/clk_in scanchain_26/clk_in scanchain_25/data_in scanchain_26/data_in
+ scanchain_25/latch_enable_in scanchain_26/latch_enable_in scanchain_25/module_data_in[0]
+ scanchain_25/module_data_in[1] scanchain_25/module_data_in[2] scanchain_25/module_data_in[3]
+ scanchain_25/module_data_in[4] scanchain_25/module_data_in[5] scanchain_25/module_data_in[6]
+ scanchain_25/module_data_in[7] scanchain_25/module_data_out[0] scanchain_25/module_data_out[1]
+ scanchain_25/module_data_out[2] scanchain_25/module_data_out[3] scanchain_25/module_data_out[4]
+ scanchain_25/module_data_out[5] scanchain_25/module_data_out[6] scanchain_25/module_data_out[7]
+ scanchain_25/scan_select_in scanchain_26/scan_select_in vccd1 vssd1 scanchain
Xscanchain_14 scanchain_14/clk_in scanchain_15/clk_in scanchain_14/data_in scanchain_15/data_in
+ scanchain_14/latch_enable_in scanchain_15/latch_enable_in scanchain_14/module_data_in[0]
+ scanchain_14/module_data_in[1] scanchain_14/module_data_in[2] scanchain_14/module_data_in[3]
+ scanchain_14/module_data_in[4] scanchain_14/module_data_in[5] scanchain_14/module_data_in[6]
+ scanchain_14/module_data_in[7] scanchain_14/module_data_out[0] scanchain_14/module_data_out[1]
+ scanchain_14/module_data_out[2] scanchain_14/module_data_out[3] scanchain_14/module_data_out[4]
+ scanchain_14/module_data_out[5] scanchain_14/module_data_out[6] scanchain_14/module_data_out[7]
+ scanchain_14/scan_select_in scanchain_15/scan_select_in vccd1 vssd1 scanchain
Xscanchain_69 scanchain_69/clk_in scanchain_70/clk_in scanchain_69/data_in scanchain_70/data_in
+ scanchain_69/latch_enable_in scanchain_70/latch_enable_in scanchain_69/module_data_in[0]
+ scanchain_69/module_data_in[1] scanchain_69/module_data_in[2] scanchain_69/module_data_in[3]
+ scanchain_69/module_data_in[4] scanchain_69/module_data_in[5] scanchain_69/module_data_in[6]
+ scanchain_69/module_data_in[7] scanchain_69/module_data_out[0] scanchain_69/module_data_out[1]
+ scanchain_69/module_data_out[2] scanchain_69/module_data_out[3] scanchain_69/module_data_out[4]
+ scanchain_69/module_data_out[5] scanchain_69/module_data_out[6] scanchain_69/module_data_out[7]
+ scanchain_69/scan_select_in scanchain_70/scan_select_in vccd1 vssd1 scanchain
Xscanchain_58 scanchain_58/clk_in scanchain_59/clk_in scanchain_58/data_in scanchain_59/data_in
+ scanchain_58/latch_enable_in scanchain_59/latch_enable_in scanchain_58/module_data_in[0]
+ scanchain_58/module_data_in[1] scanchain_58/module_data_in[2] scanchain_58/module_data_in[3]
+ scanchain_58/module_data_in[4] scanchain_58/module_data_in[5] scanchain_58/module_data_in[6]
+ scanchain_58/module_data_in[7] scanchain_58/module_data_out[0] scanchain_58/module_data_out[1]
+ scanchain_58/module_data_out[2] scanchain_58/module_data_out[3] scanchain_58/module_data_out[4]
+ scanchain_58/module_data_out[5] scanchain_58/module_data_out[6] scanchain_58/module_data_out[7]
+ scanchain_58/scan_select_in scanchain_59/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_438 scanchain_438/module_data_in[0] scanchain_438/module_data_in[1]
+ scanchain_438/module_data_in[2] scanchain_438/module_data_in[3] scanchain_438/module_data_in[4]
+ scanchain_438/module_data_in[5] scanchain_438/module_data_in[6] scanchain_438/module_data_in[7]
+ scanchain_438/module_data_out[0] scanchain_438/module_data_out[1] scanchain_438/module_data_out[2]
+ scanchain_438/module_data_out[3] scanchain_438/module_data_out[4] scanchain_438/module_data_out[5]
+ scanchain_438/module_data_out[6] scanchain_438/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_449 scanchain_449/module_data_in[0] scanchain_449/module_data_in[1]
+ scanchain_449/module_data_in[2] scanchain_449/module_data_in[3] scanchain_449/module_data_in[4]
+ scanchain_449/module_data_in[5] scanchain_449/module_data_in[6] scanchain_449/module_data_in[7]
+ scanchain_449/module_data_out[0] scanchain_449/module_data_out[1] scanchain_449/module_data_out[2]
+ scanchain_449/module_data_out[3] scanchain_449/module_data_out[4] scanchain_449/module_data_out[5]
+ scanchain_449/module_data_out[6] scanchain_449/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_427 scanchain_427/module_data_in[0] scanchain_427/module_data_in[1]
+ scanchain_427/module_data_in[2] scanchain_427/module_data_in[3] scanchain_427/module_data_in[4]
+ scanchain_427/module_data_in[5] scanchain_427/module_data_in[6] scanchain_427/module_data_in[7]
+ scanchain_427/module_data_out[0] scanchain_427/module_data_out[1] scanchain_427/module_data_out[2]
+ scanchain_427/module_data_out[3] scanchain_427/module_data_out[4] scanchain_427/module_data_out[5]
+ scanchain_427/module_data_out[6] scanchain_427/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_416 scanchain_416/module_data_in[0] scanchain_416/module_data_in[1]
+ scanchain_416/module_data_in[2] scanchain_416/module_data_in[3] scanchain_416/module_data_in[4]
+ scanchain_416/module_data_in[5] scanchain_416/module_data_in[6] scanchain_416/module_data_in[7]
+ scanchain_416/module_data_out[0] scanchain_416/module_data_out[1] scanchain_416/module_data_out[2]
+ scanchain_416/module_data_out[3] scanchain_416/module_data_out[4] scanchain_416/module_data_out[5]
+ scanchain_416/module_data_out[6] scanchain_416/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_405 scanchain_405/module_data_in[0] scanchain_405/module_data_in[1]
+ scanchain_405/module_data_in[2] scanchain_405/module_data_in[3] scanchain_405/module_data_in[4]
+ scanchain_405/module_data_in[5] scanchain_405/module_data_in[6] scanchain_405/module_data_in[7]
+ scanchain_405/module_data_out[0] scanchain_405/module_data_out[1] scanchain_405/module_data_out[2]
+ scanchain_405/module_data_out[3] scanchain_405/module_data_out[4] scanchain_405/module_data_out[5]
+ scanchain_405/module_data_out[6] scanchain_405/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_279 scanchain_279/module_data_in[0] scanchain_279/module_data_in[1]
+ scanchain_279/module_data_in[2] scanchain_279/module_data_in[3] scanchain_279/module_data_in[4]
+ scanchain_279/module_data_in[5] scanchain_279/module_data_in[6] scanchain_279/module_data_in[7]
+ scanchain_279/module_data_out[0] scanchain_279/module_data_out[1] scanchain_279/module_data_out[2]
+ scanchain_279/module_data_out[3] scanchain_279/module_data_out[4] scanchain_279/module_data_out[5]
+ scanchain_279/module_data_out[6] scanchain_279/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_268 scanchain_268/module_data_in[0] scanchain_268/module_data_in[1]
+ scanchain_268/module_data_in[2] scanchain_268/module_data_in[3] scanchain_268/module_data_in[4]
+ scanchain_268/module_data_in[5] scanchain_268/module_data_in[6] scanchain_268/module_data_in[7]
+ scanchain_268/module_data_out[0] scanchain_268/module_data_out[1] scanchain_268/module_data_out[2]
+ scanchain_268/module_data_out[3] scanchain_268/module_data_out[4] scanchain_268/module_data_out[5]
+ scanchain_268/module_data_out[6] scanchain_268/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_246 scanchain_246/module_data_in[0] scanchain_246/module_data_in[1]
+ scanchain_246/module_data_in[2] scanchain_246/module_data_in[3] scanchain_246/module_data_in[4]
+ scanchain_246/module_data_in[5] scanchain_246/module_data_in[6] scanchain_246/module_data_in[7]
+ scanchain_246/module_data_out[0] scanchain_246/module_data_out[1] scanchain_246/module_data_out[2]
+ scanchain_246/module_data_out[3] scanchain_246/module_data_out[4] scanchain_246/module_data_out[5]
+ scanchain_246/module_data_out[6] scanchain_246/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_257 scanchain_257/module_data_in[0] scanchain_257/module_data_in[1]
+ scanchain_257/module_data_in[2] scanchain_257/module_data_in[3] scanchain_257/module_data_in[4]
+ scanchain_257/module_data_in[5] scanchain_257/module_data_in[6] scanchain_257/module_data_in[7]
+ scanchain_257/module_data_out[0] scanchain_257/module_data_out[1] scanchain_257/module_data_out[2]
+ scanchain_257/module_data_out[3] scanchain_257/module_data_out[4] scanchain_257/module_data_out[5]
+ scanchain_257/module_data_out[6] scanchain_257/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_235 scanchain_235/module_data_in[0] scanchain_235/module_data_in[1]
+ scanchain_235/module_data_in[2] scanchain_235/module_data_in[3] scanchain_235/module_data_in[4]
+ scanchain_235/module_data_in[5] scanchain_235/module_data_in[6] scanchain_235/module_data_in[7]
+ scanchain_235/module_data_out[0] scanchain_235/module_data_out[1] scanchain_235/module_data_out[2]
+ scanchain_235/module_data_out[3] scanchain_235/module_data_out[4] scanchain_235/module_data_out[5]
+ scanchain_235/module_data_out[6] scanchain_235/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_213 scanchain_213/module_data_in[0] scanchain_213/module_data_in[1]
+ scanchain_213/module_data_in[2] scanchain_213/module_data_in[3] scanchain_213/module_data_in[4]
+ scanchain_213/module_data_in[5] scanchain_213/module_data_in[6] scanchain_213/module_data_in[7]
+ scanchain_213/module_data_out[0] scanchain_213/module_data_out[1] scanchain_213/module_data_out[2]
+ scanchain_213/module_data_out[3] scanchain_213/module_data_out[4] scanchain_213/module_data_out[5]
+ scanchain_213/module_data_out[6] scanchain_213/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_224 scanchain_224/module_data_in[0] scanchain_224/module_data_in[1]
+ scanchain_224/module_data_in[2] scanchain_224/module_data_in[3] scanchain_224/module_data_in[4]
+ scanchain_224/module_data_in[5] scanchain_224/module_data_in[6] scanchain_224/module_data_in[7]
+ scanchain_224/module_data_out[0] scanchain_224/module_data_out[1] scanchain_224/module_data_out[2]
+ scanchain_224/module_data_out[3] scanchain_224/module_data_out[4] scanchain_224/module_data_out[5]
+ scanchain_224/module_data_out[6] scanchain_224/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_202 scanchain_202/module_data_in[0] scanchain_202/module_data_in[1]
+ scanchain_202/module_data_in[2] scanchain_202/module_data_in[3] scanchain_202/module_data_in[4]
+ scanchain_202/module_data_in[5] scanchain_202/module_data_in[6] scanchain_202/module_data_in[7]
+ scanchain_202/module_data_out[0] scanchain_202/module_data_out[1] scanchain_202/module_data_out[2]
+ scanchain_202/module_data_out[3] scanchain_202/module_data_out[4] scanchain_202/module_data_out[5]
+ scanchain_202/module_data_out[6] scanchain_202/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscan_controller io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18]
+ io_in[19] io_in[20] wb_clk_i io_in[8] io_in[9] io_in[21] io_in[22] io_in[23] io_in[24]
+ io_in[25] io_in[26] io_in[27] io_in[28] la_data_in[0] la_data_in[1] la_data_out[0]
+ la_data_in[3] la_data_in[2] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[29] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35]
+ io_out[36] io_out[37] wb_rst_i scanchain_472/clk_out scanchain_0/clk_in scanchain_472/data_out
+ scanchain_0/data_in scanchain_0/latch_enable_in scanchain_0/scan_select_in io_in[11]
+ io_out[10] vccd1 vssd1 scan_controller
Xuser_module_339501025136214612_66 scanchain_66/module_data_in[0] scanchain_66/module_data_in[1]
+ scanchain_66/module_data_in[2] scanchain_66/module_data_in[3] scanchain_66/module_data_in[4]
+ scanchain_66/module_data_in[5] scanchain_66/module_data_in[6] scanchain_66/module_data_in[7]
+ scanchain_66/module_data_out[0] scanchain_66/module_data_out[1] scanchain_66/module_data_out[2]
+ scanchain_66/module_data_out[3] scanchain_66/module_data_out[4] scanchain_66/module_data_out[5]
+ scanchain_66/module_data_out[6] scanchain_66/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_77 scanchain_77/module_data_in[0] scanchain_77/module_data_in[1]
+ scanchain_77/module_data_in[2] scanchain_77/module_data_in[3] scanchain_77/module_data_in[4]
+ scanchain_77/module_data_in[5] scanchain_77/module_data_in[6] scanchain_77/module_data_in[7]
+ scanchain_77/module_data_out[0] scanchain_77/module_data_out[1] scanchain_77/module_data_out[2]
+ scanchain_77/module_data_out[3] scanchain_77/module_data_out[4] scanchain_77/module_data_out[5]
+ scanchain_77/module_data_out[6] scanchain_77/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_88 scanchain_88/module_data_in[0] scanchain_88/module_data_in[1]
+ scanchain_88/module_data_in[2] scanchain_88/module_data_in[3] scanchain_88/module_data_in[4]
+ scanchain_88/module_data_in[5] scanchain_88/module_data_in[6] scanchain_88/module_data_in[7]
+ scanchain_88/module_data_out[0] scanchain_88/module_data_out[1] scanchain_88/module_data_out[2]
+ scanchain_88/module_data_out[3] scanchain_88/module_data_out[4] scanchain_88/module_data_out[5]
+ scanchain_88/module_data_out[6] scanchain_88/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_99 scanchain_99/module_data_in[0] scanchain_99/module_data_in[1]
+ scanchain_99/module_data_in[2] scanchain_99/module_data_in[3] scanchain_99/module_data_in[4]
+ scanchain_99/module_data_in[5] scanchain_99/module_data_in[6] scanchain_99/module_data_in[7]
+ scanchain_99/module_data_out[0] scanchain_99/module_data_out[1] scanchain_99/module_data_out[2]
+ scanchain_99/module_data_out[3] scanchain_99/module_data_out[4] scanchain_99/module_data_out[5]
+ scanchain_99/module_data_out[6] scanchain_99/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_393 scanchain_393/clk_in scanchain_394/clk_in scanchain_393/data_in scanchain_394/data_in
+ scanchain_393/latch_enable_in scanchain_394/latch_enable_in scanchain_393/module_data_in[0]
+ scanchain_393/module_data_in[1] scanchain_393/module_data_in[2] scanchain_393/module_data_in[3]
+ scanchain_393/module_data_in[4] scanchain_393/module_data_in[5] scanchain_393/module_data_in[6]
+ scanchain_393/module_data_in[7] scanchain_393/module_data_out[0] scanchain_393/module_data_out[1]
+ scanchain_393/module_data_out[2] scanchain_393/module_data_out[3] scanchain_393/module_data_out[4]
+ scanchain_393/module_data_out[5] scanchain_393/module_data_out[6] scanchain_393/module_data_out[7]
+ scanchain_393/scan_select_in scanchain_394/scan_select_in vccd1 vssd1 scanchain
Xscanchain_382 scanchain_382/clk_in scanchain_383/clk_in scanchain_382/data_in scanchain_383/data_in
+ scanchain_382/latch_enable_in scanchain_383/latch_enable_in scanchain_382/module_data_in[0]
+ scanchain_382/module_data_in[1] scanchain_382/module_data_in[2] scanchain_382/module_data_in[3]
+ scanchain_382/module_data_in[4] scanchain_382/module_data_in[5] scanchain_382/module_data_in[6]
+ scanchain_382/module_data_in[7] scanchain_382/module_data_out[0] scanchain_382/module_data_out[1]
+ scanchain_382/module_data_out[2] scanchain_382/module_data_out[3] scanchain_382/module_data_out[4]
+ scanchain_382/module_data_out[5] scanchain_382/module_data_out[6] scanchain_382/module_data_out[7]
+ scanchain_382/scan_select_in scanchain_383/scan_select_in vccd1 vssd1 scanchain
Xscanchain_360 scanchain_360/clk_in scanchain_361/clk_in scanchain_360/data_in scanchain_361/data_in
+ scanchain_360/latch_enable_in scanchain_361/latch_enable_in scanchain_360/module_data_in[0]
+ scanchain_360/module_data_in[1] scanchain_360/module_data_in[2] scanchain_360/module_data_in[3]
+ scanchain_360/module_data_in[4] scanchain_360/module_data_in[5] scanchain_360/module_data_in[6]
+ scanchain_360/module_data_in[7] scanchain_360/module_data_out[0] scanchain_360/module_data_out[1]
+ scanchain_360/module_data_out[2] scanchain_360/module_data_out[3] scanchain_360/module_data_out[4]
+ scanchain_360/module_data_out[5] scanchain_360/module_data_out[6] scanchain_360/module_data_out[7]
+ scanchain_360/scan_select_in scanchain_361/scan_select_in vccd1 vssd1 scanchain
Xscanchain_371 scanchain_371/clk_in scanchain_372/clk_in scanchain_371/data_in scanchain_372/data_in
+ scanchain_371/latch_enable_in scanchain_372/latch_enable_in scanchain_371/module_data_in[0]
+ scanchain_371/module_data_in[1] scanchain_371/module_data_in[2] scanchain_371/module_data_in[3]
+ scanchain_371/module_data_in[4] scanchain_371/module_data_in[5] scanchain_371/module_data_in[6]
+ scanchain_371/module_data_in[7] scanchain_371/module_data_out[0] scanchain_371/module_data_out[1]
+ scanchain_371/module_data_out[2] scanchain_371/module_data_out[3] scanchain_371/module_data_out[4]
+ scanchain_371/module_data_out[5] scanchain_371/module_data_out[6] scanchain_371/module_data_out[7]
+ scanchain_371/scan_select_in scanchain_372/scan_select_in vccd1 vssd1 scanchain
Xscanchain_37 scanchain_37/clk_in scanchain_38/clk_in scanchain_37/data_in scanchain_38/data_in
+ scanchain_37/latch_enable_in scanchain_38/latch_enable_in scanchain_37/module_data_in[0]
+ scanchain_37/module_data_in[1] scanchain_37/module_data_in[2] scanchain_37/module_data_in[3]
+ scanchain_37/module_data_in[4] scanchain_37/module_data_in[5] scanchain_37/module_data_in[6]
+ scanchain_37/module_data_in[7] scanchain_37/module_data_out[0] scanchain_37/module_data_out[1]
+ scanchain_37/module_data_out[2] scanchain_37/module_data_out[3] scanchain_37/module_data_out[4]
+ scanchain_37/module_data_out[5] scanchain_37/module_data_out[6] scanchain_37/module_data_out[7]
+ scanchain_37/scan_select_in scanchain_38/scan_select_in vccd1 vssd1 scanchain
Xscanchain_26 scanchain_26/clk_in scanchain_27/clk_in scanchain_26/data_in scanchain_27/data_in
+ scanchain_26/latch_enable_in scanchain_27/latch_enable_in mm21_LEDMatrixTop_26/io_in[0]
+ mm21_LEDMatrixTop_26/io_in[1] mm21_LEDMatrixTop_26/io_in[2] mm21_LEDMatrixTop_26/io_in[3]
+ mm21_LEDMatrixTop_26/io_in[4] mm21_LEDMatrixTop_26/io_in[5] mm21_LEDMatrixTop_26/io_in[6]
+ mm21_LEDMatrixTop_26/io_in[7] mm21_LEDMatrixTop_26/io_out[0] mm21_LEDMatrixTop_26/io_out[1]
+ mm21_LEDMatrixTop_26/io_out[2] mm21_LEDMatrixTop_26/io_out[3] mm21_LEDMatrixTop_26/io_out[4]
+ mm21_LEDMatrixTop_26/io_out[5] mm21_LEDMatrixTop_26/io_out[6] mm21_LEDMatrixTop_26/io_out[7]
+ scanchain_26/scan_select_in scanchain_27/scan_select_in vccd1 vssd1 scanchain
Xscanchain_15 scanchain_15/clk_in scanchain_16/clk_in scanchain_15/data_in scanchain_16/data_in
+ scanchain_15/latch_enable_in scanchain_16/latch_enable_in tiny_fft_15/io_in[0] tiny_fft_15/io_in[1]
+ tiny_fft_15/io_in[2] tiny_fft_15/io_in[3] tiny_fft_15/io_in[4] tiny_fft_15/io_in[5]
+ tiny_fft_15/io_in[6] tiny_fft_15/io_in[7] tiny_fft_15/io_out[0] tiny_fft_15/io_out[1]
+ tiny_fft_15/io_out[2] tiny_fft_15/io_out[3] tiny_fft_15/io_out[4] tiny_fft_15/io_out[5]
+ tiny_fft_15/io_out[6] tiny_fft_15/io_out[7] scanchain_15/scan_select_in scanchain_16/scan_select_in
+ vccd1 vssd1 scanchain
Xscanchain_48 scanchain_48/clk_in scanchain_49/clk_in scanchain_48/data_in scanchain_49/data_in
+ scanchain_48/latch_enable_in scanchain_49/latch_enable_in scanchain_48/module_data_in[0]
+ scanchain_48/module_data_in[1] scanchain_48/module_data_in[2] scanchain_48/module_data_in[3]
+ scanchain_48/module_data_in[4] scanchain_48/module_data_in[5] scanchain_48/module_data_in[6]
+ scanchain_48/module_data_in[7] scanchain_48/module_data_out[0] scanchain_48/module_data_out[1]
+ scanchain_48/module_data_out[2] scanchain_48/module_data_out[3] scanchain_48/module_data_out[4]
+ scanchain_48/module_data_out[5] scanchain_48/module_data_out[6] scanchain_48/module_data_out[7]
+ scanchain_48/scan_select_in scanchain_49/scan_select_in vccd1 vssd1 scanchain
Xscanchain_59 scanchain_59/clk_in scanchain_60/clk_in scanchain_59/data_in scanchain_60/data_in
+ scanchain_59/latch_enable_in scanchain_60/latch_enable_in scanchain_59/module_data_in[0]
+ scanchain_59/module_data_in[1] scanchain_59/module_data_in[2] scanchain_59/module_data_in[3]
+ scanchain_59/module_data_in[4] scanchain_59/module_data_in[5] scanchain_59/module_data_in[6]
+ scanchain_59/module_data_in[7] scanchain_59/module_data_out[0] scanchain_59/module_data_out[1]
+ scanchain_59/module_data_out[2] scanchain_59/module_data_out[3] scanchain_59/module_data_out[4]
+ scanchain_59/module_data_out[5] scanchain_59/module_data_out[6] scanchain_59/module_data_out[7]
+ scanchain_59/scan_select_in scanchain_60/scan_select_in vccd1 vssd1 scanchain
Xscanchain_190 scanchain_190/clk_in scanchain_191/clk_in scanchain_190/data_in scanchain_191/data_in
+ scanchain_190/latch_enable_in scanchain_191/latch_enable_in scanchain_190/module_data_in[0]
+ scanchain_190/module_data_in[1] scanchain_190/module_data_in[2] scanchain_190/module_data_in[3]
+ scanchain_190/module_data_in[4] scanchain_190/module_data_in[5] scanchain_190/module_data_in[6]
+ scanchain_190/module_data_in[7] scanchain_190/module_data_out[0] scanchain_190/module_data_out[1]
+ scanchain_190/module_data_out[2] scanchain_190/module_data_out[3] scanchain_190/module_data_out[4]
+ scanchain_190/module_data_out[5] scanchain_190/module_data_out[6] scanchain_190/module_data_out[7]
+ scanchain_190/scan_select_in scanchain_191/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_439 scanchain_439/module_data_in[0] scanchain_439/module_data_in[1]
+ scanchain_439/module_data_in[2] scanchain_439/module_data_in[3] scanchain_439/module_data_in[4]
+ scanchain_439/module_data_in[5] scanchain_439/module_data_in[6] scanchain_439/module_data_in[7]
+ scanchain_439/module_data_out[0] scanchain_439/module_data_out[1] scanchain_439/module_data_out[2]
+ scanchain_439/module_data_out[3] scanchain_439/module_data_out[4] scanchain_439/module_data_out[5]
+ scanchain_439/module_data_out[6] scanchain_439/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_428 scanchain_428/module_data_in[0] scanchain_428/module_data_in[1]
+ scanchain_428/module_data_in[2] scanchain_428/module_data_in[3] scanchain_428/module_data_in[4]
+ scanchain_428/module_data_in[5] scanchain_428/module_data_in[6] scanchain_428/module_data_in[7]
+ scanchain_428/module_data_out[0] scanchain_428/module_data_out[1] scanchain_428/module_data_out[2]
+ scanchain_428/module_data_out[3] scanchain_428/module_data_out[4] scanchain_428/module_data_out[5]
+ scanchain_428/module_data_out[6] scanchain_428/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_417 scanchain_417/module_data_in[0] scanchain_417/module_data_in[1]
+ scanchain_417/module_data_in[2] scanchain_417/module_data_in[3] scanchain_417/module_data_in[4]
+ scanchain_417/module_data_in[5] scanchain_417/module_data_in[6] scanchain_417/module_data_in[7]
+ scanchain_417/module_data_out[0] scanchain_417/module_data_out[1] scanchain_417/module_data_out[2]
+ scanchain_417/module_data_out[3] scanchain_417/module_data_out[4] scanchain_417/module_data_out[5]
+ scanchain_417/module_data_out[6] scanchain_417/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_406 scanchain_406/module_data_in[0] scanchain_406/module_data_in[1]
+ scanchain_406/module_data_in[2] scanchain_406/module_data_in[3] scanchain_406/module_data_in[4]
+ scanchain_406/module_data_in[5] scanchain_406/module_data_in[6] scanchain_406/module_data_in[7]
+ scanchain_406/module_data_out[0] scanchain_406/module_data_out[1] scanchain_406/module_data_out[2]
+ scanchain_406/module_data_out[3] scanchain_406/module_data_out[4] scanchain_406/module_data_out[5]
+ scanchain_406/module_data_out[6] scanchain_406/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_214 scanchain_214/module_data_in[0] scanchain_214/module_data_in[1]
+ scanchain_214/module_data_in[2] scanchain_214/module_data_in[3] scanchain_214/module_data_in[4]
+ scanchain_214/module_data_in[5] scanchain_214/module_data_in[6] scanchain_214/module_data_in[7]
+ scanchain_214/module_data_out[0] scanchain_214/module_data_out[1] scanchain_214/module_data_out[2]
+ scanchain_214/module_data_out[3] scanchain_214/module_data_out[4] scanchain_214/module_data_out[5]
+ scanchain_214/module_data_out[6] scanchain_214/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_225 scanchain_225/module_data_in[0] scanchain_225/module_data_in[1]
+ scanchain_225/module_data_in[2] scanchain_225/module_data_in[3] scanchain_225/module_data_in[4]
+ scanchain_225/module_data_in[5] scanchain_225/module_data_in[6] scanchain_225/module_data_in[7]
+ scanchain_225/module_data_out[0] scanchain_225/module_data_out[1] scanchain_225/module_data_out[2]
+ scanchain_225/module_data_out[3] scanchain_225/module_data_out[4] scanchain_225/module_data_out[5]
+ scanchain_225/module_data_out[6] scanchain_225/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_203 scanchain_203/module_data_in[0] scanchain_203/module_data_in[1]
+ scanchain_203/module_data_in[2] scanchain_203/module_data_in[3] scanchain_203/module_data_in[4]
+ scanchain_203/module_data_in[5] scanchain_203/module_data_in[6] scanchain_203/module_data_in[7]
+ scanchain_203/module_data_out[0] scanchain_203/module_data_out[1] scanchain_203/module_data_out[2]
+ scanchain_203/module_data_out[3] scanchain_203/module_data_out[4] scanchain_203/module_data_out[5]
+ scanchain_203/module_data_out[6] scanchain_203/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xyupferris_bitslam_40 yupferris_bitslam_40/io_in[0] yupferris_bitslam_40/io_in[1]
+ yupferris_bitslam_40/io_in[2] yupferris_bitslam_40/io_in[3] yupferris_bitslam_40/io_in[4]
+ yupferris_bitslam_40/io_in[5] yupferris_bitslam_40/io_in[6] yupferris_bitslam_40/io_in[7]
+ yupferris_bitslam_40/io_out[0] yupferris_bitslam_40/io_out[1] yupferris_bitslam_40/io_out[2]
+ yupferris_bitslam_40/io_out[3] yupferris_bitslam_40/io_out[4] yupferris_bitslam_40/io_out[5]
+ yupferris_bitslam_40/io_out[6] yupferris_bitslam_40/io_out[7] vccd1 vssd1 yupferris_bitslam
Xxyz_peppergray_Potato1_top_30 scanchain_30/module_data_in[0] scanchain_30/module_data_in[1]
+ scanchain_30/module_data_in[2] scanchain_30/module_data_in[3] scanchain_30/module_data_in[4]
+ scanchain_30/module_data_in[5] scanchain_30/module_data_in[6] scanchain_30/module_data_in[7]
+ scanchain_30/module_data_out[0] scanchain_30/module_data_out[1] scanchain_30/module_data_out[2]
+ scanchain_30/module_data_out[3] scanchain_30/module_data_out[4] scanchain_30/module_data_out[5]
+ scanchain_30/module_data_out[6] scanchain_30/module_data_out[7] vccd1 vssd1 xyz_peppergray_Potato1_top
Xuser_module_339501025136214612_269 scanchain_269/module_data_in[0] scanchain_269/module_data_in[1]
+ scanchain_269/module_data_in[2] scanchain_269/module_data_in[3] scanchain_269/module_data_in[4]
+ scanchain_269/module_data_in[5] scanchain_269/module_data_in[6] scanchain_269/module_data_in[7]
+ scanchain_269/module_data_out[0] scanchain_269/module_data_out[1] scanchain_269/module_data_out[2]
+ scanchain_269/module_data_out[3] scanchain_269/module_data_out[4] scanchain_269/module_data_out[5]
+ scanchain_269/module_data_out[6] scanchain_269/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_247 scanchain_247/module_data_in[0] scanchain_247/module_data_in[1]
+ scanchain_247/module_data_in[2] scanchain_247/module_data_in[3] scanchain_247/module_data_in[4]
+ scanchain_247/module_data_in[5] scanchain_247/module_data_in[6] scanchain_247/module_data_in[7]
+ scanchain_247/module_data_out[0] scanchain_247/module_data_out[1] scanchain_247/module_data_out[2]
+ scanchain_247/module_data_out[3] scanchain_247/module_data_out[4] scanchain_247/module_data_out[5]
+ scanchain_247/module_data_out[6] scanchain_247/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_258 scanchain_258/module_data_in[0] scanchain_258/module_data_in[1]
+ scanchain_258/module_data_in[2] scanchain_258/module_data_in[3] scanchain_258/module_data_in[4]
+ scanchain_258/module_data_in[5] scanchain_258/module_data_in[6] scanchain_258/module_data_in[7]
+ scanchain_258/module_data_out[0] scanchain_258/module_data_out[1] scanchain_258/module_data_out[2]
+ scanchain_258/module_data_out[3] scanchain_258/module_data_out[4] scanchain_258/module_data_out[5]
+ scanchain_258/module_data_out[6] scanchain_258/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_236 scanchain_236/module_data_in[0] scanchain_236/module_data_in[1]
+ scanchain_236/module_data_in[2] scanchain_236/module_data_in[3] scanchain_236/module_data_in[4]
+ scanchain_236/module_data_in[5] scanchain_236/module_data_in[6] scanchain_236/module_data_in[7]
+ scanchain_236/module_data_out[0] scanchain_236/module_data_out[1] scanchain_236/module_data_out[2]
+ scanchain_236/module_data_out[3] scanchain_236/module_data_out[4] scanchain_236/module_data_out[5]
+ scanchain_236/module_data_out[6] scanchain_236/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xchase_the_beat_20 chase_the_beat_20/io_in[0] chase_the_beat_20/io_in[1] chase_the_beat_20/io_in[2]
+ chase_the_beat_20/io_in[3] chase_the_beat_20/io_in[4] chase_the_beat_20/io_in[5]
+ chase_the_beat_20/io_in[6] chase_the_beat_20/io_in[7] chase_the_beat_20/io_out[0]
+ chase_the_beat_20/io_out[1] chase_the_beat_20/io_out[2] chase_the_beat_20/io_out[3]
+ chase_the_beat_20/io_out[4] chase_the_beat_20/io_out[5] chase_the_beat_20/io_out[6]
+ chase_the_beat_20/io_out[7] vccd1 vssd1 chase_the_beat
Xuser_module_339501025136214612_67 scanchain_67/module_data_in[0] scanchain_67/module_data_in[1]
+ scanchain_67/module_data_in[2] scanchain_67/module_data_in[3] scanchain_67/module_data_in[4]
+ scanchain_67/module_data_in[5] scanchain_67/module_data_in[6] scanchain_67/module_data_in[7]
+ scanchain_67/module_data_out[0] scanchain_67/module_data_out[1] scanchain_67/module_data_out[2]
+ scanchain_67/module_data_out[3] scanchain_67/module_data_out[4] scanchain_67/module_data_out[5]
+ scanchain_67/module_data_out[6] scanchain_67/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_78 scanchain_78/module_data_in[0] scanchain_78/module_data_in[1]
+ scanchain_78/module_data_in[2] scanchain_78/module_data_in[3] scanchain_78/module_data_in[4]
+ scanchain_78/module_data_in[5] scanchain_78/module_data_in[6] scanchain_78/module_data_in[7]
+ scanchain_78/module_data_out[0] scanchain_78/module_data_out[1] scanchain_78/module_data_out[2]
+ scanchain_78/module_data_out[3] scanchain_78/module_data_out[4] scanchain_78/module_data_out[5]
+ scanchain_78/module_data_out[6] scanchain_78/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_89 scanchain_89/module_data_in[0] scanchain_89/module_data_in[1]
+ scanchain_89/module_data_in[2] scanchain_89/module_data_in[3] scanchain_89/module_data_in[4]
+ scanchain_89/module_data_in[5] scanchain_89/module_data_in[6] scanchain_89/module_data_in[7]
+ scanchain_89/module_data_out[0] scanchain_89/module_data_out[1] scanchain_89/module_data_out[2]
+ scanchain_89/module_data_out[3] scanchain_89/module_data_out[4] scanchain_89/module_data_out[5]
+ scanchain_89/module_data_out[6] scanchain_89/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_394 scanchain_394/clk_in scanchain_395/clk_in scanchain_394/data_in scanchain_395/data_in
+ scanchain_394/latch_enable_in scanchain_395/latch_enable_in scanchain_394/module_data_in[0]
+ scanchain_394/module_data_in[1] scanchain_394/module_data_in[2] scanchain_394/module_data_in[3]
+ scanchain_394/module_data_in[4] scanchain_394/module_data_in[5] scanchain_394/module_data_in[6]
+ scanchain_394/module_data_in[7] scanchain_394/module_data_out[0] scanchain_394/module_data_out[1]
+ scanchain_394/module_data_out[2] scanchain_394/module_data_out[3] scanchain_394/module_data_out[4]
+ scanchain_394/module_data_out[5] scanchain_394/module_data_out[6] scanchain_394/module_data_out[7]
+ scanchain_394/scan_select_in scanchain_395/scan_select_in vccd1 vssd1 scanchain
Xscanchain_383 scanchain_383/clk_in scanchain_384/clk_in scanchain_383/data_in scanchain_384/data_in
+ scanchain_383/latch_enable_in scanchain_384/latch_enable_in scanchain_383/module_data_in[0]
+ scanchain_383/module_data_in[1] scanchain_383/module_data_in[2] scanchain_383/module_data_in[3]
+ scanchain_383/module_data_in[4] scanchain_383/module_data_in[5] scanchain_383/module_data_in[6]
+ scanchain_383/module_data_in[7] scanchain_383/module_data_out[0] scanchain_383/module_data_out[1]
+ scanchain_383/module_data_out[2] scanchain_383/module_data_out[3] scanchain_383/module_data_out[4]
+ scanchain_383/module_data_out[5] scanchain_383/module_data_out[6] scanchain_383/module_data_out[7]
+ scanchain_383/scan_select_in scanchain_384/scan_select_in vccd1 vssd1 scanchain
Xscanchain_361 scanchain_361/clk_in scanchain_362/clk_in scanchain_361/data_in scanchain_362/data_in
+ scanchain_361/latch_enable_in scanchain_362/latch_enable_in scanchain_361/module_data_in[0]
+ scanchain_361/module_data_in[1] scanchain_361/module_data_in[2] scanchain_361/module_data_in[3]
+ scanchain_361/module_data_in[4] scanchain_361/module_data_in[5] scanchain_361/module_data_in[6]
+ scanchain_361/module_data_in[7] scanchain_361/module_data_out[0] scanchain_361/module_data_out[1]
+ scanchain_361/module_data_out[2] scanchain_361/module_data_out[3] scanchain_361/module_data_out[4]
+ scanchain_361/module_data_out[5] scanchain_361/module_data_out[6] scanchain_361/module_data_out[7]
+ scanchain_361/scan_select_in scanchain_362/scan_select_in vccd1 vssd1 scanchain
Xscanchain_372 scanchain_372/clk_in scanchain_373/clk_in scanchain_372/data_in scanchain_373/data_in
+ scanchain_372/latch_enable_in scanchain_373/latch_enable_in scanchain_372/module_data_in[0]
+ scanchain_372/module_data_in[1] scanchain_372/module_data_in[2] scanchain_372/module_data_in[3]
+ scanchain_372/module_data_in[4] scanchain_372/module_data_in[5] scanchain_372/module_data_in[6]
+ scanchain_372/module_data_in[7] scanchain_372/module_data_out[0] scanchain_372/module_data_out[1]
+ scanchain_372/module_data_out[2] scanchain_372/module_data_out[3] scanchain_372/module_data_out[4]
+ scanchain_372/module_data_out[5] scanchain_372/module_data_out[6] scanchain_372/module_data_out[7]
+ scanchain_372/scan_select_in scanchain_373/scan_select_in vccd1 vssd1 scanchain
Xscanchain_350 scanchain_350/clk_in scanchain_351/clk_in scanchain_350/data_in scanchain_351/data_in
+ scanchain_350/latch_enable_in scanchain_351/latch_enable_in scanchain_350/module_data_in[0]
+ scanchain_350/module_data_in[1] scanchain_350/module_data_in[2] scanchain_350/module_data_in[3]
+ scanchain_350/module_data_in[4] scanchain_350/module_data_in[5] scanchain_350/module_data_in[6]
+ scanchain_350/module_data_in[7] scanchain_350/module_data_out[0] scanchain_350/module_data_out[1]
+ scanchain_350/module_data_out[2] scanchain_350/module_data_out[3] scanchain_350/module_data_out[4]
+ scanchain_350/module_data_out[5] scanchain_350/module_data_out[6] scanchain_350/module_data_out[7]
+ scanchain_350/scan_select_in scanchain_351/scan_select_in vccd1 vssd1 scanchain
Xscanchain_38 scanchain_38/clk_in scanchain_39/clk_in scanchain_38/data_in scanchain_39/data_in
+ scanchain_38/latch_enable_in scanchain_39/latch_enable_in thezoq2_yafpga_38/io_in[0]
+ thezoq2_yafpga_38/io_in[1] thezoq2_yafpga_38/io_in[2] thezoq2_yafpga_38/io_in[3]
+ thezoq2_yafpga_38/io_in[4] thezoq2_yafpga_38/io_in[5] thezoq2_yafpga_38/io_in[6]
+ thezoq2_yafpga_38/io_in[7] thezoq2_yafpga_38/io_out[0] thezoq2_yafpga_38/io_out[1]
+ thezoq2_yafpga_38/io_out[2] thezoq2_yafpga_38/io_out[3] thezoq2_yafpga_38/io_out[4]
+ thezoq2_yafpga_38/io_out[5] thezoq2_yafpga_38/io_out[6] thezoq2_yafpga_38/io_out[7]
+ scanchain_38/scan_select_in scanchain_39/scan_select_in vccd1 vssd1 scanchain
Xscanchain_27 scanchain_27/clk_in scanchain_28/clk_in scanchain_27/data_in scanchain_28/data_in
+ scanchain_27/latch_enable_in scanchain_28/latch_enable_in scanchain_27/module_data_in[0]
+ scanchain_27/module_data_in[1] scanchain_27/module_data_in[2] scanchain_27/module_data_in[3]
+ scanchain_27/module_data_in[4] scanchain_27/module_data_in[5] scanchain_27/module_data_in[6]
+ scanchain_27/module_data_in[7] scanchain_27/module_data_out[0] scanchain_27/module_data_out[1]
+ scanchain_27/module_data_out[2] scanchain_27/module_data_out[3] scanchain_27/module_data_out[4]
+ scanchain_27/module_data_out[5] scanchain_27/module_data_out[6] scanchain_27/module_data_out[7]
+ scanchain_27/scan_select_in scanchain_28/scan_select_in vccd1 vssd1 scanchain
Xscanchain_16 scanchain_16/clk_in scanchain_17/clk_in scanchain_16/data_in scanchain_17/data_in
+ scanchain_16/latch_enable_in scanchain_17/latch_enable_in scanchain_16/module_data_in[0]
+ scanchain_16/module_data_in[1] scanchain_16/module_data_in[2] scanchain_16/module_data_in[3]
+ scanchain_16/module_data_in[4] scanchain_16/module_data_in[5] scanchain_16/module_data_in[6]
+ scanchain_16/module_data_in[7] scanchain_16/module_data_out[0] scanchain_16/module_data_out[1]
+ scanchain_16/module_data_out[2] scanchain_16/module_data_out[3] scanchain_16/module_data_out[4]
+ scanchain_16/module_data_out[5] scanchain_16/module_data_out[6] scanchain_16/module_data_out[7]
+ scanchain_16/scan_select_in scanchain_17/scan_select_in vccd1 vssd1 scanchain
Xscanchain_49 scanchain_49/clk_in scanchain_50/clk_in scanchain_49/data_in scanchain_50/data_in
+ scanchain_49/latch_enable_in scanchain_50/latch_enable_in scanchain_49/module_data_in[0]
+ scanchain_49/module_data_in[1] scanchain_49/module_data_in[2] scanchain_49/module_data_in[3]
+ scanchain_49/module_data_in[4] scanchain_49/module_data_in[5] scanchain_49/module_data_in[6]
+ scanchain_49/module_data_in[7] scanchain_49/module_data_out[0] scanchain_49/module_data_out[1]
+ scanchain_49/module_data_out[2] scanchain_49/module_data_out[3] scanchain_49/module_data_out[4]
+ scanchain_49/module_data_out[5] scanchain_49/module_data_out[6] scanchain_49/module_data_out[7]
+ scanchain_49/scan_select_in scanchain_50/scan_select_in vccd1 vssd1 scanchain
Xscanchain_180 scanchain_180/clk_in scanchain_181/clk_in scanchain_180/data_in scanchain_181/data_in
+ scanchain_180/latch_enable_in scanchain_181/latch_enable_in scanchain_180/module_data_in[0]
+ scanchain_180/module_data_in[1] scanchain_180/module_data_in[2] scanchain_180/module_data_in[3]
+ scanchain_180/module_data_in[4] scanchain_180/module_data_in[5] scanchain_180/module_data_in[6]
+ scanchain_180/module_data_in[7] scanchain_180/module_data_out[0] scanchain_180/module_data_out[1]
+ scanchain_180/module_data_out[2] scanchain_180/module_data_out[3] scanchain_180/module_data_out[4]
+ scanchain_180/module_data_out[5] scanchain_180/module_data_out[6] scanchain_180/module_data_out[7]
+ scanchain_180/scan_select_in scanchain_181/scan_select_in vccd1 vssd1 scanchain
Xscanchain_191 scanchain_191/clk_in scanchain_192/clk_in scanchain_191/data_in scanchain_192/data_in
+ scanchain_191/latch_enable_in scanchain_192/latch_enable_in scanchain_191/module_data_in[0]
+ scanchain_191/module_data_in[1] scanchain_191/module_data_in[2] scanchain_191/module_data_in[3]
+ scanchain_191/module_data_in[4] scanchain_191/module_data_in[5] scanchain_191/module_data_in[6]
+ scanchain_191/module_data_in[7] scanchain_191/module_data_out[0] scanchain_191/module_data_out[1]
+ scanchain_191/module_data_out[2] scanchain_191/module_data_out[3] scanchain_191/module_data_out[4]
+ scanchain_191/module_data_out[5] scanchain_191/module_data_out[6] scanchain_191/module_data_out[7]
+ scanchain_191/scan_select_in scanchain_192/scan_select_in vccd1 vssd1 scanchain
Xuser_module_342981109408072274_22 scanchain_22/module_data_in[0] scanchain_22/module_data_in[1]
+ scanchain_22/module_data_in[2] scanchain_22/module_data_in[3] scanchain_22/module_data_in[4]
+ scanchain_22/module_data_in[5] scanchain_22/module_data_in[6] scanchain_22/module_data_in[7]
+ scanchain_22/module_data_out[0] scanchain_22/module_data_out[1] scanchain_22/module_data_out[2]
+ scanchain_22/module_data_out[3] scanchain_22/module_data_out[4] scanchain_22/module_data_out[5]
+ scanchain_22/module_data_out[6] scanchain_22/module_data_out[7] vccd1 vssd1 user_module_342981109408072274
Xuser_module_339501025136214612_429 scanchain_429/module_data_in[0] scanchain_429/module_data_in[1]
+ scanchain_429/module_data_in[2] scanchain_429/module_data_in[3] scanchain_429/module_data_in[4]
+ scanchain_429/module_data_in[5] scanchain_429/module_data_in[6] scanchain_429/module_data_in[7]
+ scanchain_429/module_data_out[0] scanchain_429/module_data_out[1] scanchain_429/module_data_out[2]
+ scanchain_429/module_data_out[3] scanchain_429/module_data_out[4] scanchain_429/module_data_out[5]
+ scanchain_429/module_data_out[6] scanchain_429/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_418 scanchain_418/module_data_in[0] scanchain_418/module_data_in[1]
+ scanchain_418/module_data_in[2] scanchain_418/module_data_in[3] scanchain_418/module_data_in[4]
+ scanchain_418/module_data_in[5] scanchain_418/module_data_in[6] scanchain_418/module_data_in[7]
+ scanchain_418/module_data_out[0] scanchain_418/module_data_out[1] scanchain_418/module_data_out[2]
+ scanchain_418/module_data_out[3] scanchain_418/module_data_out[4] scanchain_418/module_data_out[5]
+ scanchain_418/module_data_out[6] scanchain_418/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_407 scanchain_407/module_data_in[0] scanchain_407/module_data_in[1]
+ scanchain_407/module_data_in[2] scanchain_407/module_data_in[3] scanchain_407/module_data_in[4]
+ scanchain_407/module_data_in[5] scanchain_407/module_data_in[6] scanchain_407/module_data_in[7]
+ scanchain_407/module_data_out[0] scanchain_407/module_data_out[1] scanchain_407/module_data_out[2]
+ scanchain_407/module_data_out[3] scanchain_407/module_data_out[4] scanchain_407/module_data_out[5]
+ scanchain_407/module_data_out[6] scanchain_407/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_348255968419643987_32 scanchain_32/module_data_in[0] scanchain_32/module_data_in[1]
+ scanchain_32/module_data_in[2] scanchain_32/module_data_in[3] scanchain_32/module_data_in[4]
+ scanchain_32/module_data_in[5] scanchain_32/module_data_in[6] scanchain_32/module_data_in[7]
+ scanchain_32/module_data_out[0] scanchain_32/module_data_out[1] scanchain_32/module_data_out[2]
+ scanchain_32/module_data_out[3] scanchain_32/module_data_out[4] scanchain_32/module_data_out[5]
+ scanchain_32/module_data_out[6] scanchain_32/module_data_out[7] vccd1 vssd1 user_module_348255968419643987
Xuser_module_339501025136214612_248 scanchain_248/module_data_in[0] scanchain_248/module_data_in[1]
+ scanchain_248/module_data_in[2] scanchain_248/module_data_in[3] scanchain_248/module_data_in[4]
+ scanchain_248/module_data_in[5] scanchain_248/module_data_in[6] scanchain_248/module_data_in[7]
+ scanchain_248/module_data_out[0] scanchain_248/module_data_out[1] scanchain_248/module_data_out[2]
+ scanchain_248/module_data_out[3] scanchain_248/module_data_out[4] scanchain_248/module_data_out[5]
+ scanchain_248/module_data_out[6] scanchain_248/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_259 scanchain_259/module_data_in[0] scanchain_259/module_data_in[1]
+ scanchain_259/module_data_in[2] scanchain_259/module_data_in[3] scanchain_259/module_data_in[4]
+ scanchain_259/module_data_in[5] scanchain_259/module_data_in[6] scanchain_259/module_data_in[7]
+ scanchain_259/module_data_out[0] scanchain_259/module_data_out[1] scanchain_259/module_data_out[2]
+ scanchain_259/module_data_out[3] scanchain_259/module_data_out[4] scanchain_259/module_data_out[5]
+ scanchain_259/module_data_out[6] scanchain_259/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_237 scanchain_237/module_data_in[0] scanchain_237/module_data_in[1]
+ scanchain_237/module_data_in[2] scanchain_237/module_data_in[3] scanchain_237/module_data_in[4]
+ scanchain_237/module_data_in[5] scanchain_237/module_data_in[6] scanchain_237/module_data_in[7]
+ scanchain_237/module_data_out[0] scanchain_237/module_data_out[1] scanchain_237/module_data_out[2]
+ scanchain_237/module_data_out[3] scanchain_237/module_data_out[4] scanchain_237/module_data_out[5]
+ scanchain_237/module_data_out[6] scanchain_237/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_226 scanchain_226/module_data_in[0] scanchain_226/module_data_in[1]
+ scanchain_226/module_data_in[2] scanchain_226/module_data_in[3] scanchain_226/module_data_in[4]
+ scanchain_226/module_data_in[5] scanchain_226/module_data_in[6] scanchain_226/module_data_in[7]
+ scanchain_226/module_data_out[0] scanchain_226/module_data_out[1] scanchain_226/module_data_out[2]
+ scanchain_226/module_data_out[3] scanchain_226/module_data_out[4] scanchain_226/module_data_out[5]
+ scanchain_226/module_data_out[6] scanchain_226/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_215 scanchain_215/module_data_in[0] scanchain_215/module_data_in[1]
+ scanchain_215/module_data_in[2] scanchain_215/module_data_in[3] scanchain_215/module_data_in[4]
+ scanchain_215/module_data_in[5] scanchain_215/module_data_in[6] scanchain_215/module_data_in[7]
+ scanchain_215/module_data_out[0] scanchain_215/module_data_out[1] scanchain_215/module_data_out[2]
+ scanchain_215/module_data_out[3] scanchain_215/module_data_out[4] scanchain_215/module_data_out[5]
+ scanchain_215/module_data_out[6] scanchain_215/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_204 scanchain_204/module_data_in[0] scanchain_204/module_data_in[1]
+ scanchain_204/module_data_in[2] scanchain_204/module_data_in[3] scanchain_204/module_data_in[4]
+ scanchain_204/module_data_in[5] scanchain_204/module_data_in[6] scanchain_204/module_data_in[7]
+ scanchain_204/module_data_out[0] scanchain_204/module_data_out[1] scanchain_204/module_data_out[2]
+ scanchain_204/module_data_out[3] scanchain_204/module_data_out[4] scanchain_204/module_data_out[5]
+ scanchain_204/module_data_out[6] scanchain_204/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_395 scanchain_395/clk_in scanchain_396/clk_in scanchain_395/data_in scanchain_396/data_in
+ scanchain_395/latch_enable_in scanchain_396/latch_enable_in scanchain_395/module_data_in[0]
+ scanchain_395/module_data_in[1] scanchain_395/module_data_in[2] scanchain_395/module_data_in[3]
+ scanchain_395/module_data_in[4] scanchain_395/module_data_in[5] scanchain_395/module_data_in[6]
+ scanchain_395/module_data_in[7] scanchain_395/module_data_out[0] scanchain_395/module_data_out[1]
+ scanchain_395/module_data_out[2] scanchain_395/module_data_out[3] scanchain_395/module_data_out[4]
+ scanchain_395/module_data_out[5] scanchain_395/module_data_out[6] scanchain_395/module_data_out[7]
+ scanchain_395/scan_select_in scanchain_396/scan_select_in vccd1 vssd1 scanchain
Xscanchain_384 scanchain_384/clk_in scanchain_385/clk_in scanchain_384/data_in scanchain_385/data_in
+ scanchain_384/latch_enable_in scanchain_385/latch_enable_in scanchain_384/module_data_in[0]
+ scanchain_384/module_data_in[1] scanchain_384/module_data_in[2] scanchain_384/module_data_in[3]
+ scanchain_384/module_data_in[4] scanchain_384/module_data_in[5] scanchain_384/module_data_in[6]
+ scanchain_384/module_data_in[7] scanchain_384/module_data_out[0] scanchain_384/module_data_out[1]
+ scanchain_384/module_data_out[2] scanchain_384/module_data_out[3] scanchain_384/module_data_out[4]
+ scanchain_384/module_data_out[5] scanchain_384/module_data_out[6] scanchain_384/module_data_out[7]
+ scanchain_384/scan_select_in scanchain_385/scan_select_in vccd1 vssd1 scanchain
Xscanchain_362 scanchain_362/clk_in scanchain_363/clk_in scanchain_362/data_in scanchain_363/data_in
+ scanchain_362/latch_enable_in scanchain_363/latch_enable_in scanchain_362/module_data_in[0]
+ scanchain_362/module_data_in[1] scanchain_362/module_data_in[2] scanchain_362/module_data_in[3]
+ scanchain_362/module_data_in[4] scanchain_362/module_data_in[5] scanchain_362/module_data_in[6]
+ scanchain_362/module_data_in[7] scanchain_362/module_data_out[0] scanchain_362/module_data_out[1]
+ scanchain_362/module_data_out[2] scanchain_362/module_data_out[3] scanchain_362/module_data_out[4]
+ scanchain_362/module_data_out[5] scanchain_362/module_data_out[6] scanchain_362/module_data_out[7]
+ scanchain_362/scan_select_in scanchain_363/scan_select_in vccd1 vssd1 scanchain
Xscanchain_373 scanchain_373/clk_in scanchain_374/clk_in scanchain_373/data_in scanchain_374/data_in
+ scanchain_373/latch_enable_in scanchain_374/latch_enable_in scanchain_373/module_data_in[0]
+ scanchain_373/module_data_in[1] scanchain_373/module_data_in[2] scanchain_373/module_data_in[3]
+ scanchain_373/module_data_in[4] scanchain_373/module_data_in[5] scanchain_373/module_data_in[6]
+ scanchain_373/module_data_in[7] scanchain_373/module_data_out[0] scanchain_373/module_data_out[1]
+ scanchain_373/module_data_out[2] scanchain_373/module_data_out[3] scanchain_373/module_data_out[4]
+ scanchain_373/module_data_out[5] scanchain_373/module_data_out[6] scanchain_373/module_data_out[7]
+ scanchain_373/scan_select_in scanchain_374/scan_select_in vccd1 vssd1 scanchain
Xscanchain_351 scanchain_351/clk_in scanchain_352/clk_in scanchain_351/data_in scanchain_352/data_in
+ scanchain_351/latch_enable_in scanchain_352/latch_enable_in scanchain_351/module_data_in[0]
+ scanchain_351/module_data_in[1] scanchain_351/module_data_in[2] scanchain_351/module_data_in[3]
+ scanchain_351/module_data_in[4] scanchain_351/module_data_in[5] scanchain_351/module_data_in[6]
+ scanchain_351/module_data_in[7] scanchain_351/module_data_out[0] scanchain_351/module_data_out[1]
+ scanchain_351/module_data_out[2] scanchain_351/module_data_out[3] scanchain_351/module_data_out[4]
+ scanchain_351/module_data_out[5] scanchain_351/module_data_out[6] scanchain_351/module_data_out[7]
+ scanchain_351/scan_select_in scanchain_352/scan_select_in vccd1 vssd1 scanchain
Xscanchain_340 scanchain_340/clk_in scanchain_341/clk_in scanchain_340/data_in scanchain_341/data_in
+ scanchain_340/latch_enable_in scanchain_341/latch_enable_in scanchain_340/module_data_in[0]
+ scanchain_340/module_data_in[1] scanchain_340/module_data_in[2] scanchain_340/module_data_in[3]
+ scanchain_340/module_data_in[4] scanchain_340/module_data_in[5] scanchain_340/module_data_in[6]
+ scanchain_340/module_data_in[7] scanchain_340/module_data_out[0] scanchain_340/module_data_out[1]
+ scanchain_340/module_data_out[2] scanchain_340/module_data_out[3] scanchain_340/module_data_out[4]
+ scanchain_340/module_data_out[5] scanchain_340/module_data_out[6] scanchain_340/module_data_out[7]
+ scanchain_340/scan_select_in scanchain_341/scan_select_in vccd1 vssd1 scanchain
Xscanchain_39 scanchain_39/clk_in scanchain_40/clk_in scanchain_39/data_in scanchain_40/data_in
+ scanchain_39/latch_enable_in scanchain_40/latch_enable_in moyes0_top_module_39/io_in[0]
+ moyes0_top_module_39/io_in[1] moyes0_top_module_39/io_in[2] moyes0_top_module_39/io_in[3]
+ moyes0_top_module_39/io_in[4] moyes0_top_module_39/io_in[5] moyes0_top_module_39/io_in[6]
+ moyes0_top_module_39/io_in[7] moyes0_top_module_39/io_out[0] moyes0_top_module_39/io_out[1]
+ moyes0_top_module_39/io_out[2] moyes0_top_module_39/io_out[3] moyes0_top_module_39/io_out[4]
+ moyes0_top_module_39/io_out[5] moyes0_top_module_39/io_out[6] moyes0_top_module_39/io_out[7]
+ scanchain_39/scan_select_in scanchain_40/scan_select_in vccd1 vssd1 scanchain
Xscanchain_17 scanchain_17/clk_in scanchain_18/clk_in scanchain_17/data_in scanchain_18/data_in
+ scanchain_17/latch_enable_in scanchain_18/latch_enable_in scanchain_17/module_data_in[0]
+ scanchain_17/module_data_in[1] scanchain_17/module_data_in[2] scanchain_17/module_data_in[3]
+ scanchain_17/module_data_in[4] scanchain_17/module_data_in[5] scanchain_17/module_data_in[6]
+ scanchain_17/module_data_in[7] scanchain_17/module_data_out[0] scanchain_17/module_data_out[1]
+ scanchain_17/module_data_out[2] scanchain_17/module_data_out[3] scanchain_17/module_data_out[4]
+ scanchain_17/module_data_out[5] scanchain_17/module_data_out[6] scanchain_17/module_data_out[7]
+ scanchain_17/scan_select_in scanchain_18/scan_select_in vccd1 vssd1 scanchain
Xscanchain_28 scanchain_28/clk_in scanchain_29/clk_in scanchain_28/data_in scanchain_29/data_in
+ scanchain_28/latch_enable_in scanchain_29/latch_enable_in scanchain_28/module_data_in[0]
+ scanchain_28/module_data_in[1] scanchain_28/module_data_in[2] scanchain_28/module_data_in[3]
+ scanchain_28/module_data_in[4] scanchain_28/module_data_in[5] scanchain_28/module_data_in[6]
+ scanchain_28/module_data_in[7] scanchain_28/module_data_out[0] scanchain_28/module_data_out[1]
+ scanchain_28/module_data_out[2] scanchain_28/module_data_out[3] scanchain_28/module_data_out[4]
+ scanchain_28/module_data_out[5] scanchain_28/module_data_out[6] scanchain_28/module_data_out[7]
+ scanchain_28/scan_select_in scanchain_29/scan_select_in vccd1 vssd1 scanchain
Xuser_module_347592305412145748_13 scanchain_13/module_data_in[0] scanchain_13/module_data_in[1]
+ scanchain_13/module_data_in[2] scanchain_13/module_data_in[3] scanchain_13/module_data_in[4]
+ scanchain_13/module_data_in[5] scanchain_13/module_data_in[6] scanchain_13/module_data_in[7]
+ scanchain_13/module_data_out[0] scanchain_13/module_data_out[1] scanchain_13/module_data_out[2]
+ scanchain_13/module_data_out[3] scanchain_13/module_data_out[4] scanchain_13/module_data_out[5]
+ scanchain_13/module_data_out[6] scanchain_13/module_data_out[7] vccd1 vssd1 user_module_347592305412145748
Xuser_module_339501025136214612_68 scanchain_68/module_data_in[0] scanchain_68/module_data_in[1]
+ scanchain_68/module_data_in[2] scanchain_68/module_data_in[3] scanchain_68/module_data_in[4]
+ scanchain_68/module_data_in[5] scanchain_68/module_data_in[6] scanchain_68/module_data_in[7]
+ scanchain_68/module_data_out[0] scanchain_68/module_data_out[1] scanchain_68/module_data_out[2]
+ scanchain_68/module_data_out[3] scanchain_68/module_data_out[4] scanchain_68/module_data_out[5]
+ scanchain_68/module_data_out[6] scanchain_68/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_57 scanchain_57/module_data_in[0] scanchain_57/module_data_in[1]
+ scanchain_57/module_data_in[2] scanchain_57/module_data_in[3] scanchain_57/module_data_in[4]
+ scanchain_57/module_data_in[5] scanchain_57/module_data_in[6] scanchain_57/module_data_in[7]
+ scanchain_57/module_data_out[0] scanchain_57/module_data_out[1] scanchain_57/module_data_out[2]
+ scanchain_57/module_data_out[3] scanchain_57/module_data_out[4] scanchain_57/module_data_out[5]
+ scanchain_57/module_data_out[6] scanchain_57/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_79 scanchain_79/module_data_in[0] scanchain_79/module_data_in[1]
+ scanchain_79/module_data_in[2] scanchain_79/module_data_in[3] scanchain_79/module_data_in[4]
+ scanchain_79/module_data_in[5] scanchain_79/module_data_in[6] scanchain_79/module_data_in[7]
+ scanchain_79/module_data_out[0] scanchain_79/module_data_out[1] scanchain_79/module_data_out[2]
+ scanchain_79/module_data_out[3] scanchain_79/module_data_out[4] scanchain_79/module_data_out[5]
+ scanchain_79/module_data_out[6] scanchain_79/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_192 scanchain_192/clk_in scanchain_193/clk_in scanchain_192/data_in scanchain_193/data_in
+ scanchain_192/latch_enable_in scanchain_193/latch_enable_in scanchain_192/module_data_in[0]
+ scanchain_192/module_data_in[1] scanchain_192/module_data_in[2] scanchain_192/module_data_in[3]
+ scanchain_192/module_data_in[4] scanchain_192/module_data_in[5] scanchain_192/module_data_in[6]
+ scanchain_192/module_data_in[7] scanchain_192/module_data_out[0] scanchain_192/module_data_out[1]
+ scanchain_192/module_data_out[2] scanchain_192/module_data_out[3] scanchain_192/module_data_out[4]
+ scanchain_192/module_data_out[5] scanchain_192/module_data_out[6] scanchain_192/module_data_out[7]
+ scanchain_192/scan_select_in scanchain_193/scan_select_in vccd1 vssd1 scanchain
Xscanchain_181 scanchain_181/clk_in scanchain_182/clk_in scanchain_181/data_in scanchain_182/data_in
+ scanchain_181/latch_enable_in scanchain_182/latch_enable_in scanchain_181/module_data_in[0]
+ scanchain_181/module_data_in[1] scanchain_181/module_data_in[2] scanchain_181/module_data_in[3]
+ scanchain_181/module_data_in[4] scanchain_181/module_data_in[5] scanchain_181/module_data_in[6]
+ scanchain_181/module_data_in[7] scanchain_181/module_data_out[0] scanchain_181/module_data_out[1]
+ scanchain_181/module_data_out[2] scanchain_181/module_data_out[3] scanchain_181/module_data_out[4]
+ scanchain_181/module_data_out[5] scanchain_181/module_data_out[6] scanchain_181/module_data_out[7]
+ scanchain_181/scan_select_in scanchain_182/scan_select_in vccd1 vssd1 scanchain
Xscanchain_170 scanchain_170/clk_in scanchain_171/clk_in scanchain_170/data_in scanchain_171/data_in
+ scanchain_170/latch_enable_in scanchain_171/latch_enable_in scanchain_170/module_data_in[0]
+ scanchain_170/module_data_in[1] scanchain_170/module_data_in[2] scanchain_170/module_data_in[3]
+ scanchain_170/module_data_in[4] scanchain_170/module_data_in[5] scanchain_170/module_data_in[6]
+ scanchain_170/module_data_in[7] scanchain_170/module_data_out[0] scanchain_170/module_data_out[1]
+ scanchain_170/module_data_out[2] scanchain_170/module_data_out[3] scanchain_170/module_data_out[4]
+ scanchain_170/module_data_out[5] scanchain_170/module_data_out[6] scanchain_170/module_data_out[7]
+ scanchain_170/scan_select_in scanchain_171/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_419 scanchain_419/module_data_in[0] scanchain_419/module_data_in[1]
+ scanchain_419/module_data_in[2] scanchain_419/module_data_in[3] scanchain_419/module_data_in[4]
+ scanchain_419/module_data_in[5] scanchain_419/module_data_in[6] scanchain_419/module_data_in[7]
+ scanchain_419/module_data_out[0] scanchain_419/module_data_out[1] scanchain_419/module_data_out[2]
+ scanchain_419/module_data_out[3] scanchain_419/module_data_out[4] scanchain_419/module_data_out[5]
+ scanchain_419/module_data_out[6] scanchain_419/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_408 scanchain_408/module_data_in[0] scanchain_408/module_data_in[1]
+ scanchain_408/module_data_in[2] scanchain_408/module_data_in[3] scanchain_408/module_data_in[4]
+ scanchain_408/module_data_in[5] scanchain_408/module_data_in[6] scanchain_408/module_data_in[7]
+ scanchain_408/module_data_out[0] scanchain_408/module_data_out[1] scanchain_408/module_data_out[2]
+ scanchain_408/module_data_out[3] scanchain_408/module_data_out[4] scanchain_408/module_data_out[5]
+ scanchain_408/module_data_out[6] scanchain_408/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_249 scanchain_249/module_data_in[0] scanchain_249/module_data_in[1]
+ scanchain_249/module_data_in[2] scanchain_249/module_data_in[3] scanchain_249/module_data_in[4]
+ scanchain_249/module_data_in[5] scanchain_249/module_data_in[6] scanchain_249/module_data_in[7]
+ scanchain_249/module_data_out[0] scanchain_249/module_data_out[1] scanchain_249/module_data_out[2]
+ scanchain_249/module_data_out[3] scanchain_249/module_data_out[4] scanchain_249/module_data_out[5]
+ scanchain_249/module_data_out[6] scanchain_249/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_238 scanchain_238/module_data_in[0] scanchain_238/module_data_in[1]
+ scanchain_238/module_data_in[2] scanchain_238/module_data_in[3] scanchain_238/module_data_in[4]
+ scanchain_238/module_data_in[5] scanchain_238/module_data_in[6] scanchain_238/module_data_in[7]
+ scanchain_238/module_data_out[0] scanchain_238/module_data_out[1] scanchain_238/module_data_out[2]
+ scanchain_238/module_data_out[3] scanchain_238/module_data_out[4] scanchain_238/module_data_out[5]
+ scanchain_238/module_data_out[6] scanchain_238/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_227 scanchain_227/module_data_in[0] scanchain_227/module_data_in[1]
+ scanchain_227/module_data_in[2] scanchain_227/module_data_in[3] scanchain_227/module_data_in[4]
+ scanchain_227/module_data_in[5] scanchain_227/module_data_in[6] scanchain_227/module_data_in[7]
+ scanchain_227/module_data_out[0] scanchain_227/module_data_out[1] scanchain_227/module_data_out[2]
+ scanchain_227/module_data_out[3] scanchain_227/module_data_out[4] scanchain_227/module_data_out[5]
+ scanchain_227/module_data_out[6] scanchain_227/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_216 scanchain_216/module_data_in[0] scanchain_216/module_data_in[1]
+ scanchain_216/module_data_in[2] scanchain_216/module_data_in[3] scanchain_216/module_data_in[4]
+ scanchain_216/module_data_in[5] scanchain_216/module_data_in[6] scanchain_216/module_data_in[7]
+ scanchain_216/module_data_out[0] scanchain_216/module_data_out[1] scanchain_216/module_data_out[2]
+ scanchain_216/module_data_out[3] scanchain_216/module_data_out[4] scanchain_216/module_data_out[5]
+ scanchain_216/module_data_out[6] scanchain_216/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_205 scanchain_205/module_data_in[0] scanchain_205/module_data_in[1]
+ scanchain_205/module_data_in[2] scanchain_205/module_data_in[3] scanchain_205/module_data_in[4]
+ scanchain_205/module_data_in[5] scanchain_205/module_data_in[6] scanchain_205/module_data_in[7]
+ scanchain_205/module_data_out[0] scanchain_205/module_data_out[1] scanchain_205/module_data_out[2]
+ scanchain_205/module_data_out[3] scanchain_205/module_data_out[4] scanchain_205/module_data_out[5]
+ scanchain_205/module_data_out[6] scanchain_205/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_18 scanchain_18/clk_in scanchain_19/clk_in scanchain_18/data_in scanchain_19/data_in
+ scanchain_18/latch_enable_in scanchain_19/latch_enable_in scanchain_18/module_data_in[0]
+ scanchain_18/module_data_in[1] scanchain_18/module_data_in[2] scanchain_18/module_data_in[3]
+ scanchain_18/module_data_in[4] scanchain_18/module_data_in[5] scanchain_18/module_data_in[6]
+ scanchain_18/module_data_in[7] scanchain_18/module_data_out[0] scanchain_18/module_data_out[1]
+ scanchain_18/module_data_out[2] scanchain_18/module_data_out[3] scanchain_18/module_data_out[4]
+ scanchain_18/module_data_out[5] scanchain_18/module_data_out[6] scanchain_18/module_data_out[7]
+ scanchain_18/scan_select_in scanchain_19/scan_select_in vccd1 vssd1 scanchain
Xscanchain_29 scanchain_29/clk_in scanchain_30/clk_in scanchain_29/data_in scanchain_30/data_in
+ scanchain_29/latch_enable_in scanchain_30/latch_enable_in yubex_egg_timer_29/io_in[0]
+ yubex_egg_timer_29/io_in[1] yubex_egg_timer_29/io_in[2] yubex_egg_timer_29/io_in[3]
+ yubex_egg_timer_29/io_in[4] yubex_egg_timer_29/io_in[5] yubex_egg_timer_29/io_in[6]
+ yubex_egg_timer_29/io_in[7] yubex_egg_timer_29/io_out[0] yubex_egg_timer_29/io_out[1]
+ yubex_egg_timer_29/io_out[2] yubex_egg_timer_29/io_out[3] yubex_egg_timer_29/io_out[4]
+ yubex_egg_timer_29/io_out[5] yubex_egg_timer_29/io_out[6] yubex_egg_timer_29/io_out[7]
+ scanchain_29/scan_select_in scanchain_30/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_69 scanchain_69/module_data_in[0] scanchain_69/module_data_in[1]
+ scanchain_69/module_data_in[2] scanchain_69/module_data_in[3] scanchain_69/module_data_in[4]
+ scanchain_69/module_data_in[5] scanchain_69/module_data_in[6] scanchain_69/module_data_in[7]
+ scanchain_69/module_data_out[0] scanchain_69/module_data_out[1] scanchain_69/module_data_out[2]
+ scanchain_69/module_data_out[3] scanchain_69/module_data_out[4] scanchain_69/module_data_out[5]
+ scanchain_69/module_data_out[6] scanchain_69/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_58 scanchain_58/module_data_in[0] scanchain_58/module_data_in[1]
+ scanchain_58/module_data_in[2] scanchain_58/module_data_in[3] scanchain_58/module_data_in[4]
+ scanchain_58/module_data_in[5] scanchain_58/module_data_in[6] scanchain_58/module_data_in[7]
+ scanchain_58/module_data_out[0] scanchain_58/module_data_out[1] scanchain_58/module_data_out[2]
+ scanchain_58/module_data_out[3] scanchain_58/module_data_out[4] scanchain_58/module_data_out[5]
+ scanchain_58/module_data_out[6] scanchain_58/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xscanchain_396 scanchain_396/clk_in scanchain_397/clk_in scanchain_396/data_in scanchain_397/data_in
+ scanchain_396/latch_enable_in scanchain_397/latch_enable_in scanchain_396/module_data_in[0]
+ scanchain_396/module_data_in[1] scanchain_396/module_data_in[2] scanchain_396/module_data_in[3]
+ scanchain_396/module_data_in[4] scanchain_396/module_data_in[5] scanchain_396/module_data_in[6]
+ scanchain_396/module_data_in[7] scanchain_396/module_data_out[0] scanchain_396/module_data_out[1]
+ scanchain_396/module_data_out[2] scanchain_396/module_data_out[3] scanchain_396/module_data_out[4]
+ scanchain_396/module_data_out[5] scanchain_396/module_data_out[6] scanchain_396/module_data_out[7]
+ scanchain_396/scan_select_in scanchain_397/scan_select_in vccd1 vssd1 scanchain
Xscanchain_385 scanchain_385/clk_in scanchain_386/clk_in scanchain_385/data_in scanchain_386/data_in
+ scanchain_385/latch_enable_in scanchain_386/latch_enable_in scanchain_385/module_data_in[0]
+ scanchain_385/module_data_in[1] scanchain_385/module_data_in[2] scanchain_385/module_data_in[3]
+ scanchain_385/module_data_in[4] scanchain_385/module_data_in[5] scanchain_385/module_data_in[6]
+ scanchain_385/module_data_in[7] scanchain_385/module_data_out[0] scanchain_385/module_data_out[1]
+ scanchain_385/module_data_out[2] scanchain_385/module_data_out[3] scanchain_385/module_data_out[4]
+ scanchain_385/module_data_out[5] scanchain_385/module_data_out[6] scanchain_385/module_data_out[7]
+ scanchain_385/scan_select_in scanchain_386/scan_select_in vccd1 vssd1 scanchain
Xscanchain_363 scanchain_363/clk_in scanchain_364/clk_in scanchain_363/data_in scanchain_364/data_in
+ scanchain_363/latch_enable_in scanchain_364/latch_enable_in scanchain_363/module_data_in[0]
+ scanchain_363/module_data_in[1] scanchain_363/module_data_in[2] scanchain_363/module_data_in[3]
+ scanchain_363/module_data_in[4] scanchain_363/module_data_in[5] scanchain_363/module_data_in[6]
+ scanchain_363/module_data_in[7] scanchain_363/module_data_out[0] scanchain_363/module_data_out[1]
+ scanchain_363/module_data_out[2] scanchain_363/module_data_out[3] scanchain_363/module_data_out[4]
+ scanchain_363/module_data_out[5] scanchain_363/module_data_out[6] scanchain_363/module_data_out[7]
+ scanchain_363/scan_select_in scanchain_364/scan_select_in vccd1 vssd1 scanchain
Xscanchain_374 scanchain_374/clk_in scanchain_375/clk_in scanchain_374/data_in scanchain_375/data_in
+ scanchain_374/latch_enable_in scanchain_375/latch_enable_in scanchain_374/module_data_in[0]
+ scanchain_374/module_data_in[1] scanchain_374/module_data_in[2] scanchain_374/module_data_in[3]
+ scanchain_374/module_data_in[4] scanchain_374/module_data_in[5] scanchain_374/module_data_in[6]
+ scanchain_374/module_data_in[7] scanchain_374/module_data_out[0] scanchain_374/module_data_out[1]
+ scanchain_374/module_data_out[2] scanchain_374/module_data_out[3] scanchain_374/module_data_out[4]
+ scanchain_374/module_data_out[5] scanchain_374/module_data_out[6] scanchain_374/module_data_out[7]
+ scanchain_374/scan_select_in scanchain_375/scan_select_in vccd1 vssd1 scanchain
Xscanchain_352 scanchain_352/clk_in scanchain_353/clk_in scanchain_352/data_in scanchain_353/data_in
+ scanchain_352/latch_enable_in scanchain_353/latch_enable_in scanchain_352/module_data_in[0]
+ scanchain_352/module_data_in[1] scanchain_352/module_data_in[2] scanchain_352/module_data_in[3]
+ scanchain_352/module_data_in[4] scanchain_352/module_data_in[5] scanchain_352/module_data_in[6]
+ scanchain_352/module_data_in[7] scanchain_352/module_data_out[0] scanchain_352/module_data_out[1]
+ scanchain_352/module_data_out[2] scanchain_352/module_data_out[3] scanchain_352/module_data_out[4]
+ scanchain_352/module_data_out[5] scanchain_352/module_data_out[6] scanchain_352/module_data_out[7]
+ scanchain_352/scan_select_in scanchain_353/scan_select_in vccd1 vssd1 scanchain
Xscanchain_341 scanchain_341/clk_in scanchain_342/clk_in scanchain_341/data_in scanchain_342/data_in
+ scanchain_341/latch_enable_in scanchain_342/latch_enable_in scanchain_341/module_data_in[0]
+ scanchain_341/module_data_in[1] scanchain_341/module_data_in[2] scanchain_341/module_data_in[3]
+ scanchain_341/module_data_in[4] scanchain_341/module_data_in[5] scanchain_341/module_data_in[6]
+ scanchain_341/module_data_in[7] scanchain_341/module_data_out[0] scanchain_341/module_data_out[1]
+ scanchain_341/module_data_out[2] scanchain_341/module_data_out[3] scanchain_341/module_data_out[4]
+ scanchain_341/module_data_out[5] scanchain_341/module_data_out[6] scanchain_341/module_data_out[7]
+ scanchain_341/scan_select_in scanchain_342/scan_select_in vccd1 vssd1 scanchain
Xscanchain_330 scanchain_330/clk_in scanchain_331/clk_in scanchain_330/data_in scanchain_331/data_in
+ scanchain_330/latch_enable_in scanchain_331/latch_enable_in scanchain_330/module_data_in[0]
+ scanchain_330/module_data_in[1] scanchain_330/module_data_in[2] scanchain_330/module_data_in[3]
+ scanchain_330/module_data_in[4] scanchain_330/module_data_in[5] scanchain_330/module_data_in[6]
+ scanchain_330/module_data_in[7] scanchain_330/module_data_out[0] scanchain_330/module_data_out[1]
+ scanchain_330/module_data_out[2] scanchain_330/module_data_out[3] scanchain_330/module_data_out[4]
+ scanchain_330/module_data_out[5] scanchain_330/module_data_out[6] scanchain_330/module_data_out[7]
+ scanchain_330/scan_select_in scanchain_331/scan_select_in vccd1 vssd1 scanchain
Xscanchain_193 scanchain_193/clk_in scanchain_194/clk_in scanchain_193/data_in scanchain_194/data_in
+ scanchain_193/latch_enable_in scanchain_194/latch_enable_in scanchain_193/module_data_in[0]
+ scanchain_193/module_data_in[1] scanchain_193/module_data_in[2] scanchain_193/module_data_in[3]
+ scanchain_193/module_data_in[4] scanchain_193/module_data_in[5] scanchain_193/module_data_in[6]
+ scanchain_193/module_data_in[7] scanchain_193/module_data_out[0] scanchain_193/module_data_out[1]
+ scanchain_193/module_data_out[2] scanchain_193/module_data_out[3] scanchain_193/module_data_out[4]
+ scanchain_193/module_data_out[5] scanchain_193/module_data_out[6] scanchain_193/module_data_out[7]
+ scanchain_193/scan_select_in scanchain_194/scan_select_in vccd1 vssd1 scanchain
Xscanchain_160 scanchain_160/clk_in scanchain_161/clk_in scanchain_160/data_in scanchain_161/data_in
+ scanchain_160/latch_enable_in scanchain_161/latch_enable_in scanchain_160/module_data_in[0]
+ scanchain_160/module_data_in[1] scanchain_160/module_data_in[2] scanchain_160/module_data_in[3]
+ scanchain_160/module_data_in[4] scanchain_160/module_data_in[5] scanchain_160/module_data_in[6]
+ scanchain_160/module_data_in[7] scanchain_160/module_data_out[0] scanchain_160/module_data_out[1]
+ scanchain_160/module_data_out[2] scanchain_160/module_data_out[3] scanchain_160/module_data_out[4]
+ scanchain_160/module_data_out[5] scanchain_160/module_data_out[6] scanchain_160/module_data_out[7]
+ scanchain_160/scan_select_in scanchain_161/scan_select_in vccd1 vssd1 scanchain
Xscanchain_182 scanchain_182/clk_in scanchain_183/clk_in scanchain_182/data_in scanchain_183/data_in
+ scanchain_182/latch_enable_in scanchain_183/latch_enable_in scanchain_182/module_data_in[0]
+ scanchain_182/module_data_in[1] scanchain_182/module_data_in[2] scanchain_182/module_data_in[3]
+ scanchain_182/module_data_in[4] scanchain_182/module_data_in[5] scanchain_182/module_data_in[6]
+ scanchain_182/module_data_in[7] scanchain_182/module_data_out[0] scanchain_182/module_data_out[1]
+ scanchain_182/module_data_out[2] scanchain_182/module_data_out[3] scanchain_182/module_data_out[4]
+ scanchain_182/module_data_out[5] scanchain_182/module_data_out[6] scanchain_182/module_data_out[7]
+ scanchain_182/scan_select_in scanchain_183/scan_select_in vccd1 vssd1 scanchain
Xscanchain_171 scanchain_171/clk_in scanchain_172/clk_in scanchain_171/data_in scanchain_172/data_in
+ scanchain_171/latch_enable_in scanchain_172/latch_enable_in scanchain_171/module_data_in[0]
+ scanchain_171/module_data_in[1] scanchain_171/module_data_in[2] scanchain_171/module_data_in[3]
+ scanchain_171/module_data_in[4] scanchain_171/module_data_in[5] scanchain_171/module_data_in[6]
+ scanchain_171/module_data_in[7] scanchain_171/module_data_out[0] scanchain_171/module_data_out[1]
+ scanchain_171/module_data_out[2] scanchain_171/module_data_out[3] scanchain_171/module_data_out[4]
+ scanchain_171/module_data_out[5] scanchain_171/module_data_out[6] scanchain_171/module_data_out[7]
+ scanchain_171/scan_select_in scanchain_172/scan_select_in vccd1 vssd1 scanchain
Xuser_module_339501025136214612_409 scanchain_409/module_data_in[0] scanchain_409/module_data_in[1]
+ scanchain_409/module_data_in[2] scanchain_409/module_data_in[3] scanchain_409/module_data_in[4]
+ scanchain_409/module_data_in[5] scanchain_409/module_data_in[6] scanchain_409/module_data_in[7]
+ scanchain_409/module_data_out[0] scanchain_409/module_data_out[1] scanchain_409/module_data_out[2]
+ scanchain_409/module_data_out[3] scanchain_409/module_data_out[4] scanchain_409/module_data_out[5]
+ scanchain_409/module_data_out[6] scanchain_409/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_239 scanchain_239/module_data_in[0] scanchain_239/module_data_in[1]
+ scanchain_239/module_data_in[2] scanchain_239/module_data_in[3] scanchain_239/module_data_in[4]
+ scanchain_239/module_data_in[5] scanchain_239/module_data_in[6] scanchain_239/module_data_in[7]
+ scanchain_239/module_data_out[0] scanchain_239/module_data_out[1] scanchain_239/module_data_out[2]
+ scanchain_239/module_data_out[3] scanchain_239/module_data_out[4] scanchain_239/module_data_out[5]
+ scanchain_239/module_data_out[6] scanchain_239/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_228 scanchain_228/module_data_in[0] scanchain_228/module_data_in[1]
+ scanchain_228/module_data_in[2] scanchain_228/module_data_in[3] scanchain_228/module_data_in[4]
+ scanchain_228/module_data_in[5] scanchain_228/module_data_in[6] scanchain_228/module_data_in[7]
+ scanchain_228/module_data_out[0] scanchain_228/module_data_out[1] scanchain_228/module_data_out[2]
+ scanchain_228/module_data_out[3] scanchain_228/module_data_out[4] scanchain_228/module_data_out[5]
+ scanchain_228/module_data_out[6] scanchain_228/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_217 scanchain_217/module_data_in[0] scanchain_217/module_data_in[1]
+ scanchain_217/module_data_in[2] scanchain_217/module_data_in[3] scanchain_217/module_data_in[4]
+ scanchain_217/module_data_in[5] scanchain_217/module_data_in[6] scanchain_217/module_data_in[7]
+ scanchain_217/module_data_out[0] scanchain_217/module_data_out[1] scanchain_217/module_data_out[2]
+ scanchain_217/module_data_out[3] scanchain_217/module_data_out[4] scanchain_217/module_data_out[5]
+ scanchain_217/module_data_out[6] scanchain_217/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xuser_module_339501025136214612_206 scanchain_206/module_data_in[0] scanchain_206/module_data_in[1]
+ scanchain_206/module_data_in[2] scanchain_206/module_data_in[3] scanchain_206/module_data_in[4]
+ scanchain_206/module_data_in[5] scanchain_206/module_data_in[6] scanchain_206/module_data_in[7]
+ scanchain_206/module_data_out[0] scanchain_206/module_data_out[1] scanchain_206/module_data_out[2]
+ scanchain_206/module_data_out[3] scanchain_206/module_data_out[4] scanchain_206/module_data_out[5]
+ scanchain_206/module_data_out[6] scanchain_206/module_data_out[7] vccd1 vssd1 user_module_339501025136214612
Xfraserbc_simon_1 fraserbc_simon_1/io_in[0] fraserbc_simon_1/io_in[1] fraserbc_simon_1/io_in[2]
+ fraserbc_simon_1/io_in[3] fraserbc_simon_1/io_in[4] fraserbc_simon_1/io_in[5] fraserbc_simon_1/io_in[6]
+ fraserbc_simon_1/io_in[7] fraserbc_simon_1/io_out[0] fraserbc_simon_1/io_out[1]
+ fraserbc_simon_1/io_out[2] fraserbc_simon_1/io_out[3] fraserbc_simon_1/io_out[4]
+ fraserbc_simon_1/io_out[5] fraserbc_simon_1/io_out[6] fraserbc_simon_1/io_out[7]
+ vccd1 vssd1 fraserbc_simon
.ends

