VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu_top
  CLASS BLOCK ;
  FOREIGN alu_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 120.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 118.000 3.590 120.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 118.000 9.110 120.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 118.000 14.630 120.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 118.000 20.150 120.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 118.000 25.670 120.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 118.000 31.190 120.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 118.000 36.710 120.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 118.000 42.230 120.000 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 118.000 47.750 120.000 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 118.000 53.270 120.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 118.000 58.790 120.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 118.000 64.310 120.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 118.000 69.830 120.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 118.000 75.350 120.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 118.000 80.870 120.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 118.000 86.390 120.000 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.590 5.200 16.190 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.330 5.200 35.930 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.070 5.200 55.670 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.810 5.200 75.410 114.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.460 5.200 26.060 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.200 5.200 45.800 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.940 5.200 65.540 114.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 84.180 114.325 ;
      LAYER met1 ;
        RECT 0.070 5.200 86.410 114.480 ;
      LAYER met2 ;
        RECT 0.100 117.720 3.030 118.730 ;
        RECT 3.870 117.720 8.550 118.730 ;
        RECT 9.390 117.720 14.070 118.730 ;
        RECT 14.910 117.720 19.590 118.730 ;
        RECT 20.430 117.720 25.110 118.730 ;
        RECT 25.950 117.720 30.630 118.730 ;
        RECT 31.470 117.720 36.150 118.730 ;
        RECT 36.990 117.720 41.670 118.730 ;
        RECT 42.510 117.720 47.190 118.730 ;
        RECT 48.030 117.720 52.710 118.730 ;
        RECT 53.550 117.720 58.230 118.730 ;
        RECT 59.070 117.720 63.750 118.730 ;
        RECT 64.590 117.720 69.270 118.730 ;
        RECT 70.110 117.720 74.790 118.730 ;
        RECT 75.630 117.720 80.310 118.730 ;
        RECT 81.150 117.720 85.830 118.730 ;
        RECT 0.100 5.255 86.380 117.720 ;
      LAYER met3 ;
        RECT 7.425 5.275 78.595 114.405 ;
      LAYER met4 ;
        RECT 12.255 66.815 14.190 112.705 ;
        RECT 16.590 66.815 24.060 112.705 ;
        RECT 26.460 66.815 33.930 112.705 ;
        RECT 36.330 66.815 43.800 112.705 ;
        RECT 46.200 66.815 53.670 112.705 ;
        RECT 56.070 66.815 63.540 112.705 ;
        RECT 65.940 66.815 73.305 112.705 ;
  END
END alu_top
END LIBRARY

