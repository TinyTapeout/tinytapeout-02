VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tiny_kinda_pic
  CLASS BLOCK ;
  FOREIGN tiny_kinda_pic ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 170.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.000 8.800 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.000 19.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.000 29.200 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.000 39.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.000 49.600 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.000 59.800 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.000 70.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.000 80.200 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.000 90.400 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.000 100.600 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.000 110.800 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 2.000 121.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.000 131.200 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 2.000 141.400 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 2.000 151.600 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 2.000 161.800 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.090 5.200 23.690 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.830 5.200 58.430 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.570 5.200 93.170 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.310 5.200 127.910 163.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.460 5.200 41.060 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.200 5.200 75.800 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.940 5.200 110.540 163.440 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 144.440 163.285 ;
      LAYER met1 ;
        RECT 5.520 1.740 144.440 166.220 ;
      LAYER met2 ;
        RECT 6.530 1.710 143.880 166.250 ;
      LAYER met3 ;
        RECT 2.000 162.200 143.455 163.365 ;
        RECT 2.400 160.800 143.455 162.200 ;
        RECT 2.000 152.000 143.455 160.800 ;
        RECT 2.400 150.600 143.455 152.000 ;
        RECT 2.000 141.800 143.455 150.600 ;
        RECT 2.400 140.400 143.455 141.800 ;
        RECT 2.000 131.600 143.455 140.400 ;
        RECT 2.400 130.200 143.455 131.600 ;
        RECT 2.000 121.400 143.455 130.200 ;
        RECT 2.400 120.000 143.455 121.400 ;
        RECT 2.000 111.200 143.455 120.000 ;
        RECT 2.400 109.800 143.455 111.200 ;
        RECT 2.000 101.000 143.455 109.800 ;
        RECT 2.400 99.600 143.455 101.000 ;
        RECT 2.000 90.800 143.455 99.600 ;
        RECT 2.400 89.400 143.455 90.800 ;
        RECT 2.000 80.600 143.455 89.400 ;
        RECT 2.400 79.200 143.455 80.600 ;
        RECT 2.000 70.400 143.455 79.200 ;
        RECT 2.400 69.000 143.455 70.400 ;
        RECT 2.000 60.200 143.455 69.000 ;
        RECT 2.400 58.800 143.455 60.200 ;
        RECT 2.000 50.000 143.455 58.800 ;
        RECT 2.400 48.600 143.455 50.000 ;
        RECT 2.000 39.800 143.455 48.600 ;
        RECT 2.400 38.400 143.455 39.800 ;
        RECT 2.000 29.600 143.455 38.400 ;
        RECT 2.400 28.200 143.455 29.600 ;
        RECT 2.000 19.400 143.455 28.200 ;
        RECT 2.400 18.000 143.455 19.400 ;
        RECT 2.000 9.200 143.455 18.000 ;
        RECT 2.400 7.800 143.455 9.200 ;
        RECT 2.000 5.275 143.455 7.800 ;
      LAYER met4 ;
        RECT 19.615 15.815 21.690 156.225 ;
        RECT 24.090 15.815 39.060 156.225 ;
        RECT 41.460 15.815 56.430 156.225 ;
        RECT 58.830 15.815 73.800 156.225 ;
        RECT 76.200 15.815 91.170 156.225 ;
        RECT 93.570 15.815 108.540 156.225 ;
        RECT 110.940 15.815 125.910 156.225 ;
        RECT 128.310 15.815 137.705 156.225 ;
  END
END tiny_kinda_pic
END LIBRARY

