/* Automatically generated from https://wokwi.com/projects/349405063877231188 */

`default_nettype none

module user_module_349405063877231188(
  input [7:0] io_in,
  output [7:0] io_out
);
  wire net1 = io_in[3];
  wire net2 = io_in[4];
  wire net3 = io_in[5];
  wire net4 = io_in[6];
  wire net5 = io_in[7];
  wire net6 = 1'b1;
  wire net7 = 1'b1;
  wire net8 = 1'b1;
  wire net9;
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16;
  wire net17;
  wire net18;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81 = 1'b1;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152 = 1'b1;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234 = 1'b0;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;

  and_cell gate1 (

  );
  or_cell gate2 (

  );
  xor_cell gate3 (

  );
  nand_cell gate4 (

  );
  not_cell gate5 (

  );
  buffer_cell gate6 (

  );
  mux_cell mux1 (

  );
  dff_cell flipflop1 (

  );
  dff_cell flipflop2 (
    .d (net9),
    .clk (net10),
    .q (net11),
    .notq (net12)
  );
  and_cell gate7 (
    .a (net12),
    .b (net8),
    .out (net13)
  );
  and_cell gate8 (
    .a (net14),
    .b (net11),
    .out (net15)
  );
  or_cell gate9 (
    .a (net13),
    .b (net15),
    .out (net9)
  );
  not_cell gate10 (
    .in (net8),
    .out (net14)
  );
  dff_cell flipflop3 (
    .d (net16),
    .clk (net10),
    .q (net17),
    .notq (net18)
  );
  and_cell gate11 (
    .a (net18),
    .b (net19),
    .out (net20)
  );
  and_cell gate12 (
    .a (net21),
    .b (net17),
    .out (net22)
  );
  or_cell gate13 (
    .a (net20),
    .b (net22),
    .out (net16)
  );
  not_cell gate14 (
    .in (net19),
    .out (net21)
  );
  and_cell gate15 (
    .a (net23),
    .b (net11),
    .out (net24)
  );
  and_cell gate16 (
    .a (net5),
    .b (net12),
    .out (net25)
  );
  or_cell gate17 (
    .a (net24),
    .b (net25),
    .out (net19)
  );
  not_cell gate18 (
    .in (net5),
    .out (net23)
  );
  dff_cell flipflop4 (
    .d (net26),
    .clk (net10),
    .q (net27),
    .notq (net28)
  );
  and_cell gate19 (
    .a (net28),
    .b (net29),
    .out (net30)
  );
  and_cell gate20 (
    .a (net31),
    .b (net27),
    .out (net32)
  );
  or_cell gate21 (
    .a (net30),
    .b (net32),
    .out (net26)
  );
  not_cell gate22 (
    .in (net29),
    .out (net31)
  );
  and_cell gate23 (
    .a (net24),
    .b (net17),
    .out (net33)
  );
  and_cell gate24 (
    .a (net18),
    .b (net25),
    .out (net34)
  );
  or_cell gate25 (
    .a (net33),
    .b (net34),
    .out (net29)
  );
  dff_cell flipflop5 (
    .d (net35),
    .clk (net10),
    .q (net36),
    .notq (net37)
  );
  and_cell gate26 (
    .a (net37),
    .b (net38),
    .out (net39)
  );
  and_cell gate27 (
    .a (net40),
    .b (net36),
    .out (net41)
  );
  or_cell gate28 (
    .a (net39),
    .b (net41),
    .out (net35)
  );
  not_cell gate29 (
    .in (net38),
    .out (net40)
  );
  and_cell gate30 (
    .a (net33),
    .b (net27),
    .out (net42)
  );
  and_cell gate31 (
    .a (net28),
    .b (net34),
    .out (net43)
  );
  or_cell gate32 (
    .a (net42),
    .b (net43),
    .out (net38)
  );
  dff_cell flipflop6 (
    .d (net44),
    .clk (net10),
    .q (net45),
    .notq (net46)
  );
  and_cell gate33 (
    .a (net46),
    .b (net47),
    .out (net48)
  );
  and_cell gate34 (
    .a (net49),
    .b (net45),
    .out (net50)
  );
  or_cell gate35 (
    .a (net48),
    .b (net50),
    .out (net44)
  );
  not_cell gate36 (
    .in (net47),
    .out (net49)
  );
  and_cell gate37 (
    .a (net42),
    .b (net36),
    .out (net51)
  );
  and_cell gate38 (
    .a (net37),
    .b (net43),
    .out (net52)
  );
  or_cell gate39 (
    .a (net51),
    .b (net52),
    .out (net47)
  );
  dff_cell flipflop7 (
    .d (net53),
    .clk (net10),
    .q (net54),
    .notq (net55)
  );
  and_cell gate40 (
    .a (net55),
    .b (net56),
    .out (net57)
  );
  and_cell gate41 (
    .a (net58),
    .b (net54),
    .out (net59)
  );
  or_cell gate42 (
    .a (net57),
    .b (net59),
    .out (net53)
  );
  not_cell gate43 (
    .in (net56),
    .out (net58)
  );
  and_cell gate44 (
    .a (net51),
    .b (net45),
    .out (net60)
  );
  and_cell gate45 (
    .a (net46),
    .b (net52),
    .out (net61)
  );
  or_cell gate46 (
    .a (net60),
    .b (net61),
    .out (net56)
  );
  dff_cell flipflop8 (
    .d (net62),
    .clk (net10),
    .q (net63),
    .notq (net64)
  );
  and_cell gate47 (
    .a (net64),
    .b (net65),
    .out (net66)
  );
  and_cell gate48 (
    .a (net67),
    .b (net63),
    .out (net68)
  );
  or_cell gate49 (
    .a (net66),
    .b (net68),
    .out (net62)
  );
  not_cell gate50 (
    .in (net65),
    .out (net67)
  );
  and_cell gate51 (
    .a (net60),
    .b (net54),
    .out (net69)
  );
  and_cell gate52 (
    .a (net55),
    .b (net61),
    .out (net70)
  );
  or_cell gate53 (
    .a (net69),
    .b (net70),
    .out (net65)
  );
  dff_cell flipflop9 (
    .d (net71),
    .clk (net10),
    .q (net72),
    .notq (net73)
  );
  and_cell gate54 (
    .a (net73),
    .b (net74),
    .out (net75)
  );
  and_cell gate55 (
    .a (net76),
    .b (net72),
    .out (net77)
  );
  or_cell gate56 (
    .a (net75),
    .b (net77),
    .out (net71)
  );
  not_cell gate57 (
    .in (net74),
    .out (net76)
  );
  and_cell gate58 (
    .a (net69),
    .b (net63),
    .out (net78)
  );
  and_cell gate59 (
    .a (net64),
    .b (net70),
    .out (net79)
  );
  or_cell gate60 (
    .a (net78),
    .b (net79),
    .out (net74)
  );
  not_cell gate114 (
    .in (net5),
    .out (net80)
  );
  dff_cell flipflop10 (
    .d (net82),
    .clk (net83),
    .q (net84),
    .notq (net85)
  );
  and_cell gate61 (
    .a (net85),
    .b (net81),
    .out (net86)
  );
  and_cell gate62 (
    .a (net87),
    .b (net84),
    .out (net88)
  );
  or_cell gate63 (
    .a (net86),
    .b (net88),
    .out (net82)
  );
  not_cell gate64 (
    .in (net81),
    .out (net87)
  );
  dff_cell flipflop11 (
    .d (net89),
    .clk (net83),
    .q (net90),
    .notq (net91)
  );
  and_cell gate65 (
    .a (net91),
    .b (net92),
    .out (net93)
  );
  and_cell gate66 (
    .a (net94),
    .b (net90),
    .out (net95)
  );
  or_cell gate67 (
    .a (net93),
    .b (net95),
    .out (net89)
  );
  not_cell gate68 (
    .in (net92),
    .out (net94)
  );
  and_cell gate69 (
    .a (net80),
    .b (net84),
    .out (net96)
  );
  and_cell gate70 (
    .a (net5),
    .b (net85),
    .out (net97)
  );
  or_cell gate71 (
    .a (net96),
    .b (net97),
    .out (net92)
  );
  dff_cell flipflop12 (
    .d (net98),
    .clk (net83),
    .q (net99),
    .notq (net100)
  );
  and_cell gate72 (
    .a (net100),
    .b (net101),
    .out (net102)
  );
  and_cell gate73 (
    .a (net103),
    .b (net99),
    .out (net104)
  );
  or_cell gate74 (
    .a (net102),
    .b (net104),
    .out (net98)
  );
  not_cell gate75 (
    .in (net101),
    .out (net103)
  );
  and_cell gate76 (
    .a (net96),
    .b (net90),
    .out (net105)
  );
  and_cell gate77 (
    .a (net91),
    .b (net97),
    .out (net106)
  );
  or_cell gate78 (
    .a (net105),
    .b (net106),
    .out (net101)
  );
  dff_cell flipflop13 (
    .d (net107),
    .clk (net83),
    .q (net108),
    .notq (net109)
  );
  and_cell gate79 (
    .a (net109),
    .b (net110),
    .out (net111)
  );
  and_cell gate80 (
    .a (net112),
    .b (net108),
    .out (net113)
  );
  or_cell gate81 (
    .a (net111),
    .b (net113),
    .out (net107)
  );
  not_cell gate82 (
    .in (net110),
    .out (net112)
  );
  and_cell gate83 (
    .a (net105),
    .b (net99),
    .out (net114)
  );
  and_cell gate84 (
    .a (net100),
    .b (net106),
    .out (net115)
  );
  or_cell gate85 (
    .a (net114),
    .b (net115),
    .out (net110)
  );
  dff_cell flipflop14 (
    .d (net116),
    .clk (net83),
    .q (net117),
    .notq (net118)
  );
  and_cell gate86 (
    .a (net118),
    .b (net119),
    .out (net120)
  );
  and_cell gate87 (
    .a (net121),
    .b (net117),
    .out (net122)
  );
  or_cell gate88 (
    .a (net120),
    .b (net122),
    .out (net116)
  );
  not_cell gate89 (
    .in (net119),
    .out (net121)
  );
  and_cell gate90 (
    .a (net114),
    .b (net108),
    .out (net123)
  );
  and_cell gate91 (
    .a (net109),
    .b (net115),
    .out (net124)
  );
  or_cell gate92 (
    .a (net123),
    .b (net124),
    .out (net119)
  );
  dff_cell flipflop15 (
    .d (net125),
    .clk (net83),
    .q (net126),
    .notq (net127)
  );
  and_cell gate93 (
    .a (net127),
    .b (net128),
    .out (net129)
  );
  and_cell gate94 (
    .a (net130),
    .b (net126),
    .out (net131)
  );
  or_cell gate95 (
    .a (net129),
    .b (net131),
    .out (net125)
  );
  not_cell gate96 (
    .in (net128),
    .out (net130)
  );
  and_cell gate97 (
    .a (net123),
    .b (net117),
    .out (net132)
  );
  and_cell gate98 (
    .a (net118),
    .b (net124),
    .out (net133)
  );
  or_cell gate99 (
    .a (net132),
    .b (net133),
    .out (net128)
  );
  dff_cell flipflop16 (
    .d (net134),
    .clk (net83),
    .q (net135),
    .notq (net136)
  );
  and_cell gate100 (
    .a (net136),
    .b (net137),
    .out (net138)
  );
  and_cell gate101 (
    .a (net139),
    .b (net135),
    .out (net140)
  );
  or_cell gate102 (
    .a (net138),
    .b (net140),
    .out (net134)
  );
  not_cell gate103 (
    .in (net137),
    .out (net139)
  );
  and_cell gate104 (
    .a (net132),
    .b (net126),
    .out (net141)
  );
  and_cell gate105 (
    .a (net127),
    .b (net133),
    .out (net142)
  );
  or_cell gate106 (
    .a (net141),
    .b (net142),
    .out (net137)
  );
  dff_cell flipflop17 (
    .d (net143),
    .clk (net83),
    .q (net144),
    .notq (net145)
  );
  and_cell gate107 (
    .a (net145),
    .b (net146),
    .out (net147)
  );
  and_cell gate108 (
    .a (net148),
    .b (net144),
    .out (net149)
  );
  or_cell gate109 (
    .a (net147),
    .b (net149),
    .out (net143)
  );
  not_cell gate110 (
    .in (net146),
    .out (net148)
  );
  and_cell gate111 (
    .a (net141),
    .b (net135),
    .out (net150)
  );
  and_cell gate112 (
    .a (net136),
    .b (net142),
    .out (net151)
  );
  or_cell gate113 (
    .a (net150),
    .b (net151),
    .out (net146)
  );
  and_cell gate115 (
    .a (net1),
    .b (net4),
    .out (net10)
  );
  and_cell gate116 (
    .a (net153),
    .b (net1),
    .out (net83)
  );
  not_cell gate117 (
    .in (net4),
    .out (net153)
  );
  not_cell gate118 (

  );
  not_cell gate130 (

  );
  not_cell gate131 (

  );
  buffer_cell gate132 (
    .in (net154),
    .out (net155)
  );
  buffer_cell gate133 (
    .in (net156),
    .out (net157)
  );
  buffer_cell gate134 (
    .in (net158),
    .out (net159)
  );
  buffer_cell gate135 (
    .in (net160),
    .out (net161)
  );
  not_cell gate136 (
    .in (net159),
    .out (net162)
  );
  not_cell gate137 (
    .in (net161),
    .out (net163)
  );
  not_cell gate138 (
    .in (net157),
    .out (net164)
  );
  not_cell gate139 (
    .in (net155),
    .out (net165)
  );
  and_cell gate140 (
    .a (net159),
    .b (net166),
    .out (net167)
  );
  and_cell gate141 (
    .a (net165),
    .b (net157),
    .out (net166)
  );
  or_cell gate142 (
    .a (net168),
    .b (net169),
    .out (net170)
  );
  and_cell gate143 (
    .a (net155),
    .b (net162),
    .out (net171)
  );
  and_cell gate144 (
    .a (net163),
    .b (net172),
    .out (net173)
  );
  and_cell gate145 (
    .a (net164),
    .b (net155),
    .out (net172)
  );
  and_cell gate146 (
    .a (net161),
    .b (net165),
    .out (net174)
  );
  and_cell gate147 (
    .a (net157),
    .b (net161),
    .out (net175)
  );
  or_cell gate148 (
    .a (net176),
    .b (net175),
    .out (net177)
  );
  or_cell gate149 (
    .a (net174),
    .b (net167),
    .out (net178)
  );
  or_cell gate150 (
    .a (net173),
    .b (net171),
    .out (net169)
  );
  or_cell gate151 (
    .a (net177),
    .b (net178),
    .out (net168)
  );
  and_cell gate152 (
    .a (net155),
    .b (net179),
    .out (net180)
  );
  and_cell gate153 (
    .a (net163),
    .b (net159),
    .out (net179)
  );
  and_cell gate154 (
    .a (net164),
    .b (net162),
    .out (net176)
  );
  and_cell gate155 (
    .a (net165),
    .b (net181),
    .out (net182)
  );
  and_cell gate156 (
    .a (net163),
    .b (net162),
    .out (net181)
  );
  and_cell gate157 (
    .a (net165),
    .b (net161),
    .out (net183)
  );
  and_cell gate158 (
    .a (net183),
    .b (net159),
    .out (net184)
  );
  and_cell gate159 (
    .a (net165),
    .b (net164),
    .out (net185)
  );
  or_cell gate160 (
    .a (net180),
    .b (net185),
    .out (net186)
  );
  or_cell gate161 (
    .a (net184),
    .b (net182),
    .out (net187)
  );
  or_cell gate162 (
    .a (net186),
    .b (net187),
    .out (net188)
  );
  or_cell gate163 (
    .a (net188),
    .b (net176),
    .out (net189)
  );
  and_cell gate164 (
    .a (net155),
    .b (net164),
    .out (net190)
  );
  and_cell gate165 (
    .a (net165),
    .b (net157),
    .out (net191)
  );
  and_cell gate166 (
    .a (net165),
    .b (net163),
    .out (net192)
  );
  and_cell gate167 (
    .a (net165),
    .b (net159),
    .out (net193)
  );
  and_cell gate168 (
    .a (net159),
    .b (net163),
    .out (net194)
  );
  or_cell gate169 (
    .a (net190),
    .b (net191),
    .out (net195)
  );
  or_cell gate170 (
    .a (net192),
    .b (net193),
    .out (net196)
  );
  or_cell gate171 (
    .a (net195),
    .b (net196),
    .out (net197)
  );
  or_cell gate172 (
    .a (net197),
    .b (net194),
    .out (net198)
  );
  and_cell gate173 (
    .a (net157),
    .b (net163),
    .out (net199)
  );
  and_cell gate174 (
    .a (net165),
    .b (net161),
    .out (net200)
  );
  and_cell gate175 (
    .a (net155),
    .b (net157),
    .out (net201)
  );
  and_cell gate176 (
    .a (net199),
    .b (net159),
    .out (net202)
  );
  and_cell gate177 (
    .a (net200),
    .b (net162),
    .out (net203)
  );
  and_cell gate178 (
    .a (net201),
    .b (net162),
    .out (net204)
  );
  and_cell gate179 (
    .a (net164),
    .b (net163),
    .out (net205)
  );
  and_cell gate180 (
    .a (net164),
    .b (net161),
    .out (net206)
  );
  and_cell gate181 (
    .a (net205),
    .b (net162),
    .out (net207)
  );
  and_cell gate182 (
    .a (net206),
    .b (net159),
    .out (net208)
  );
  or_cell gate183 (
    .a (net204),
    .b (net203),
    .out (net209)
  );
  or_cell gate184 (
    .a (net202),
    .b (net208),
    .out (net210)
  );
  or_cell gate185 (
    .a (net209),
    .b (net210),
    .out (net211)
  );
  or_cell gate186 (
    .a (net211),
    .b (net207),
    .out (net212)
  );
  and_cell gate187 (
    .a (net155),
    .b (net161),
    .out (net213)
  );
  and_cell gate188 (
    .a (net155),
    .b (net157),
    .out (net214)
  );
  and_cell gate189 (
    .a (net161),
    .b (net162),
    .out (net215)
  );
  or_cell gate190 (
    .a (net214),
    .b (net213),
    .out (net216)
  );
  or_cell gate191 (
    .a (net176),
    .b (net215),
    .out (net217)
  );
  or_cell gate192 (
    .a (net216),
    .b (net217),
    .out (net218)
  );
  and_cell gate193 (
    .a (net155),
    .b (net164),
    .out (net219)
  );
  and_cell gate194 (
    .a (net192),
    .b (net157),
    .out (net220)
  );
  and_cell gate195 (
    .a (net157),
    .b (net162),
    .out (net221)
  );
  or_cell gate196 (
    .a (net219),
    .b (net213),
    .out (net222)
  );
  or_cell gate197 (
    .a (net220),
    .b (net221),
    .out (net223)
  );
  or_cell gate198 (
    .a (net222),
    .b (net223),
    .out (net224)
  );
  or_cell gate199 (
    .a (net224),
    .b (net181),
    .out (net225)
  );
  and_cell gate200 (
    .a (net219),
    .b (net226),
    .out (net227)
  );
  and_cell gate201 (
    .a (net155),
    .b (net159),
    .out (net228)
  );
  or_cell gate202 (
    .a (net219),
    .b (net220),
    .out (net229)
  );
  or_cell gate203 (
    .a (net228),
    .b (net230),
    .out (net231)
  );
  and_cell gate204 (
    .a (net164),
    .b (net161),
    .out (net230)
  );
  or_cell gate205 (
    .a (net229),
    .b (net231),
    .out (net232)
  );
  or_cell gate206 (
    .a (net215),
    .b (net232),
    .out (net233)
  );
  and_cell gate207 (
    .a (net161),
    .b (net159),
    .out (net226)
  );
  mux_cell mux5 (
    .a (net11),
    .b (net84),
    .sel (net235),
    .out (net236)
  );
  or_cell gate208 (
    .a (net237),
    .b (net238),
    .out (net158)
  );
  not_cell gate209 (
    .in (net2),
    .out (net239)
  );
  and_cell gate210 (
    .a (net2),
    .b (net240),
    .out (net241)
  );
  mux_cell mux6 (
    .a (net36),
    .b (net108),
    .sel (net235),
    .out (net242)
  );
  mux_cell mux7 (
    .a (net27),
    .b (net99),
    .sel (net235),
    .out (net243)
  );
  mux_cell mux8 (
    .a (net17),
    .b (net90),
    .sel (net235),
    .out (net240)
  );
  mux_cell mux9 (
    .a (net45),
    .b (net117),
    .sel (net235),
    .out (net244)
  );
  mux_cell mux10 (
    .a (net72),
    .b (net144),
    .sel (net235),
    .out (net245)
  );
  mux_cell mux11 (
    .a (net63),
    .b (net135),
    .sel (net235),
    .out (net246)
  );
  mux_cell mux12 (
    .a (net54),
    .b (net126),
    .sel (net235),
    .out (net247)
  );
  and_cell gate211 (
    .a (net2),
    .b (net236),
    .out (net237)
  );
  and_cell gate212 (
    .a (net2),
    .b (net243),
    .out (net248)
  );
  and_cell gate213 (
    .a (net2),
    .b (net242),
    .out (net249)
  );
  and_cell gate214 (
    .a (net250),
    .b (net247),
    .out (net251)
  );
  and_cell gate215 (
    .a (net239),
    .b (net244),
    .out (net238)
  );
  and_cell gate216 (
    .a (net252),
    .b (net246),
    .out (net253)
  );
  and_cell gate217 (
    .a (net254),
    .b (net245),
    .out (net255)
  );
  not_cell gate218 (
    .in (net2),
    .out (net250)
  );
  not_cell gate219 (
    .in (net2),
    .out (net252)
  );
  not_cell gate220 (
    .in (net2),
    .out (net254)
  );
  or_cell gate221 (
    .a (net249),
    .b (net255),
    .out (net154)
  );
  or_cell gate222 (
    .a (net248),
    .b (net253),
    .out (net156)
  );
  or_cell gate223 (
    .a (net241),
    .b (net251),
    .out (net160)
  );
  not_cell not1 (
    .in (net3),
    .out (net235)
  );
endmodule
