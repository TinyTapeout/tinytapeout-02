magic
tech sky130B
magscale 1 2
timestamp 1665589554
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 26234 700816 26240 700868
rect 26292 700856 26298 700868
rect 105446 700856 105452 700868
rect 26292 700828 105452 700856
rect 26292 700816 26298 700828
rect 105446 700816 105452 700828
rect 105504 700816 105510 700868
rect 56594 700748 56600 700800
rect 56652 700788 56658 700800
rect 202782 700788 202788 700800
rect 56652 700760 202788 700788
rect 56652 700748 56658 700760
rect 202782 700748 202788 700760
rect 202840 700748 202846 700800
rect 65518 700680 65524 700732
rect 65576 700720 65582 700732
rect 267642 700720 267648 700732
rect 65576 700692 267648 700720
rect 65576 700680 65582 700692
rect 267642 700680 267648 700692
rect 267700 700680 267706 700732
rect 17954 700612 17960 700664
rect 18012 700652 18018 700664
rect 235166 700652 235172 700664
rect 18012 700624 235172 700652
rect 18012 700612 18018 700624
rect 235166 700612 235172 700624
rect 235224 700612 235230 700664
rect 59354 700544 59360 700596
rect 59412 700584 59418 700596
rect 332502 700584 332508 700596
rect 59412 700556 332508 700584
rect 59412 700544 59418 700556
rect 332502 700544 332508 700556
rect 332560 700544 332566 700596
rect 13722 700476 13728 700528
rect 13780 700516 13786 700528
rect 300118 700516 300124 700528
rect 13780 700488 300124 700516
rect 13780 700476 13786 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 64138 700408 64144 700460
rect 64196 700448 64202 700460
rect 364978 700448 364984 700460
rect 64196 700420 364984 700448
rect 64196 700408 64202 700420
rect 364978 700408 364984 700420
rect 365036 700408 365042 700460
rect 23474 700340 23480 700392
rect 23532 700380 23538 700392
rect 462314 700380 462320 700392
rect 23532 700352 462320 700380
rect 23532 700340 23538 700352
rect 462314 700340 462320 700352
rect 462372 700340 462378 700392
rect 47026 700272 47032 700324
rect 47084 700312 47090 700324
rect 494790 700312 494796 700324
rect 47084 700284 494796 700312
rect 47084 700272 47090 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 52454 696940 52460 696992
rect 52512 696980 52518 696992
rect 580166 696980 580172 696992
rect 52512 696952 580172 696980
rect 52512 696940 52518 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 657432 3424 657484
rect 3476 657472 3482 657484
rect 8938 657472 8944 657484
rect 3476 657444 8944 657472
rect 3476 657432 3482 657444
rect 8938 657432 8944 657444
rect 8996 657432 9002 657484
rect 2774 632068 2780 632120
rect 2832 632108 2838 632120
rect 4798 632108 4804 632120
rect 2832 632080 4804 632108
rect 2832 632068 2838 632080
rect 4798 632068 4804 632080
rect 4856 632068 4862 632120
rect 64230 590656 64236 590708
rect 64288 590696 64294 590708
rect 580166 590696 580172 590708
rect 64288 590668 580172 590696
rect 64288 590656 64294 590668
rect 580166 590656 580172 590668
rect 580224 590656 580230 590708
rect 2958 579640 2964 579692
rect 3016 579680 3022 579692
rect 6178 579680 6184 579692
rect 3016 579652 6184 579680
rect 3016 579640 3022 579652
rect 6178 579640 6184 579652
rect 6236 579640 6242 579692
rect 16574 563048 16580 563100
rect 16632 563088 16638 563100
rect 580166 563088 580172 563100
rect 16632 563060 580172 563088
rect 16632 563048 16638 563060
rect 580166 563048 580172 563060
rect 580224 563048 580230 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 11698 553432 11704 553444
rect 3476 553404 11704 553432
rect 3476 553392 3482 553404
rect 11698 553392 11704 553404
rect 11756 553392 11762 553444
rect 64322 536800 64328 536852
rect 64380 536840 64386 536852
rect 580166 536840 580172 536852
rect 64380 536812 580172 536840
rect 64380 536800 64386 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 7558 527184 7564 527196
rect 3476 527156 7564 527184
rect 3476 527144 3482 527156
rect 7558 527144 7564 527156
rect 7616 527144 7622 527196
rect 24854 510620 24860 510672
rect 24912 510660 24918 510672
rect 580166 510660 580172 510672
rect 24912 510632 580172 510660
rect 24912 510620 24918 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 64414 470568 64420 470620
rect 64472 470608 64478 470620
rect 579982 470608 579988 470620
rect 64472 470580 579988 470608
rect 64472 470568 64478 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 19978 448576 19984 448588
rect 3200 448548 19984 448576
rect 3200 448536 3206 448548
rect 19978 448536 19984 448548
rect 20036 448536 20042 448588
rect 13630 430584 13636 430636
rect 13688 430624 13694 430636
rect 579614 430624 579620 430636
rect 13688 430596 579620 430624
rect 13688 430584 13694 430596
rect 579614 430584 579620 430596
rect 579672 430584 579678 430636
rect 15194 404336 15200 404388
rect 15252 404376 15258 404388
rect 580166 404376 580172 404388
rect 15252 404348 580172 404376
rect 15252 404336 15258 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 64506 378156 64512 378208
rect 64564 378196 64570 378208
rect 580166 378196 580172 378208
rect 64564 378168 580172 378196
rect 64564 378156 64570 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 3326 357416 3332 357468
rect 3384 357456 3390 357468
rect 61286 357456 61292 357468
rect 3384 357428 61292 357456
rect 3384 357416 3390 357428
rect 61286 357416 61292 357428
rect 61344 357416 61350 357468
rect 2774 345176 2780 345228
rect 2832 345216 2838 345228
rect 4890 345216 4896 345228
rect 2832 345188 4896 345216
rect 2832 345176 2838 345188
rect 4890 345176 4896 345188
rect 4948 345176 4954 345228
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 9030 292584 9036 292596
rect 3384 292556 9036 292584
rect 3384 292544 3390 292556
rect 9030 292544 9036 292556
rect 9088 292544 9094 292596
rect 3142 253920 3148 253972
rect 3200 253960 3206 253972
rect 29638 253960 29644 253972
rect 3200 253932 29644 253960
rect 3200 253920 3206 253932
rect 29638 253920 29644 253932
rect 29696 253920 29702 253972
rect 34514 231820 34520 231872
rect 34572 231860 34578 231872
rect 579798 231860 579804 231872
rect 34572 231832 579804 231860
rect 34572 231820 34578 231832
rect 579798 231820 579804 231832
rect 579856 231820 579862 231872
rect 3326 201492 3332 201544
rect 3384 201532 3390 201544
rect 61194 201532 61200 201544
rect 3384 201504 61200 201532
rect 3384 201492 3390 201504
rect 61194 201492 61200 201504
rect 61252 201492 61258 201544
rect 60826 191836 60832 191888
rect 60884 191876 60890 191888
rect 580166 191876 580172 191888
rect 60884 191848 580172 191876
rect 60884 191836 60890 191848
rect 580166 191836 580172 191848
rect 580224 191836 580230 191888
rect 51074 151784 51080 151836
rect 51132 151824 51138 151836
rect 579982 151824 579988 151836
rect 51132 151796 579988 151824
rect 51132 151784 51138 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 3326 136620 3332 136672
rect 3384 136660 3390 136672
rect 11790 136660 11796 136672
rect 3384 136632 11796 136660
rect 3384 136620 3390 136632
rect 11790 136620 11796 136632
rect 11848 136620 11854 136672
rect 64598 111800 64604 111852
rect 64656 111840 64662 111852
rect 579982 111840 579988 111852
rect 64656 111812 579988 111840
rect 64656 111800 64662 111812
rect 579982 111800 579988 111812
rect 580040 111800 580046 111852
rect 3234 44208 3240 44260
rect 3292 44248 3298 44260
rect 9122 44248 9128 44260
rect 3292 44220 9128 44248
rect 3292 44208 3298 44220
rect 9122 44208 9128 44220
rect 9180 44208 9186 44260
rect 248506 44044 248512 44056
rect 220188 44016 248512 44044
rect 220188 43988 220216 44016
rect 248506 44004 248512 44016
rect 248564 44004 248570 44056
rect 249058 44004 249064 44056
rect 249116 44044 249122 44056
rect 277486 44044 277492 44056
rect 249116 44016 277492 44044
rect 249116 44004 249122 44016
rect 277486 44004 277492 44016
rect 277544 44004 277550 44056
rect 306466 44044 306472 44056
rect 278148 44016 306472 44044
rect 278148 43988 278176 44016
rect 306466 44004 306472 44016
rect 306524 44004 306530 44056
rect 307018 44004 307024 44056
rect 307076 44044 307082 44056
rect 333146 44044 333152 44056
rect 307076 44016 333152 44044
rect 307076 44004 307082 44016
rect 333146 44004 333152 44016
rect 333204 44004 333210 44056
rect 335998 44004 336004 44056
rect 336056 44044 336062 44056
rect 362126 44044 362132 44056
rect 336056 44016 362132 44044
rect 336056 44004 336062 44016
rect 362126 44004 362132 44016
rect 362184 44004 362190 44056
rect 364978 44004 364984 44056
rect 365036 44044 365042 44056
rect 391106 44044 391112 44056
rect 365036 44016 391112 44044
rect 365036 44004 365042 44016
rect 391106 44004 391112 44016
rect 391164 44004 391170 44056
rect 393958 44004 393964 44056
rect 394016 44044 394022 44056
rect 420086 44044 420092 44056
rect 394016 44016 420092 44044
rect 394016 44004 394022 44016
rect 420086 44004 420092 44016
rect 420144 44004 420150 44056
rect 423030 44004 423036 44056
rect 423088 44044 423094 44056
rect 451366 44044 451372 44056
rect 423088 44016 451372 44044
rect 423088 44004 423094 44016
rect 451366 44004 451372 44016
rect 451424 44004 451430 44056
rect 480346 44044 480352 44056
rect 451936 44016 480352 44044
rect 220170 43936 220176 43988
rect 220228 43936 220234 43988
rect 220354 43936 220360 43988
rect 220412 43976 220418 43988
rect 248414 43976 248420 43988
rect 220412 43948 248420 43976
rect 220412 43936 220418 43948
rect 248414 43936 248420 43948
rect 248472 43936 248478 43988
rect 249242 43936 249248 43988
rect 249300 43976 249306 43988
rect 277394 43976 277400 43988
rect 249300 43948 277400 43976
rect 249300 43936 249306 43948
rect 277394 43936 277400 43948
rect 277452 43936 277458 43988
rect 278130 43936 278136 43988
rect 278188 43936 278194 43988
rect 304074 43976 304080 43988
rect 278240 43948 304080 43976
rect 278038 43868 278044 43920
rect 278096 43908 278102 43920
rect 278240 43908 278268 43948
rect 304074 43936 304080 43948
rect 304132 43936 304138 43988
rect 307110 43936 307116 43988
rect 307168 43976 307174 43988
rect 335446 43976 335452 43988
rect 307168 43948 335452 43976
rect 307168 43936 307174 43948
rect 335446 43936 335452 43948
rect 335504 43936 335510 43988
rect 336090 43936 336096 43988
rect 336148 43976 336154 43988
rect 364426 43976 364432 43988
rect 336148 43948 364432 43976
rect 336148 43936 336154 43948
rect 364426 43936 364432 43948
rect 364484 43936 364490 43988
rect 365070 43936 365076 43988
rect 365128 43976 365134 43988
rect 393406 43976 393412 43988
rect 365128 43948 393412 43976
rect 365128 43936 365134 43948
rect 393406 43936 393412 43948
rect 393464 43936 393470 43988
rect 394050 43936 394056 43988
rect 394108 43976 394114 43988
rect 422386 43976 422392 43988
rect 394108 43948 422392 43976
rect 394108 43936 394114 43948
rect 422386 43936 422392 43948
rect 422444 43936 422450 43988
rect 422938 43936 422944 43988
rect 422996 43976 423002 43988
rect 449066 43976 449072 43988
rect 422996 43948 449072 43976
rect 422996 43936 423002 43948
rect 449066 43936 449072 43948
rect 449124 43936 449130 43988
rect 278096 43880 278268 43908
rect 278096 43868 278102 43880
rect 278314 43868 278320 43920
rect 278372 43908 278378 43920
rect 306558 43908 306564 43920
rect 278372 43880 306564 43908
rect 278372 43868 278378 43880
rect 306558 43868 306564 43880
rect 306616 43868 306622 43920
rect 307202 43868 307208 43920
rect 307260 43908 307266 43920
rect 335354 43908 335360 43920
rect 307260 43880 335360 43908
rect 307260 43868 307266 43880
rect 335354 43868 335360 43880
rect 335412 43868 335418 43920
rect 336182 43868 336188 43920
rect 336240 43908 336246 43920
rect 364334 43908 364340 43920
rect 336240 43880 364340 43908
rect 336240 43868 336246 43880
rect 364334 43868 364340 43880
rect 364392 43868 364398 43920
rect 365162 43868 365168 43920
rect 365220 43908 365226 43920
rect 393314 43908 393320 43920
rect 365220 43880 393320 43908
rect 365220 43868 365226 43880
rect 393314 43868 393320 43880
rect 393372 43868 393378 43920
rect 394142 43868 394148 43920
rect 394200 43908 394206 43920
rect 422294 43908 422300 43920
rect 394200 43880 422300 43908
rect 394200 43868 394206 43880
rect 422294 43868 422300 43880
rect 422352 43868 422358 43920
rect 423122 43868 423128 43920
rect 423180 43908 423186 43920
rect 451458 43908 451464 43920
rect 423180 43880 451464 43908
rect 423180 43868 423186 43880
rect 451458 43868 451464 43880
rect 451516 43868 451522 43920
rect 451936 43908 451964 44016
rect 480346 44004 480352 44016
rect 480404 44004 480410 44056
rect 509326 44044 509332 44056
rect 481100 44016 509332 44044
rect 481100 43988 481128 44016
rect 509326 44004 509332 44016
rect 509384 44004 509390 44056
rect 509970 44004 509976 44056
rect 510028 44044 510034 44056
rect 538214 44044 538220 44056
rect 510028 44016 538220 44044
rect 510028 44004 510034 44016
rect 538214 44004 538220 44016
rect 538272 44004 538278 44056
rect 538858 44004 538864 44056
rect 538916 44044 538922 44056
rect 565078 44044 565084 44056
rect 538916 44016 565084 44044
rect 538916 44004 538922 44016
rect 565078 44004 565084 44016
rect 565136 44004 565142 44056
rect 452010 43936 452016 43988
rect 452068 43976 452074 43988
rect 480254 43976 480260 43988
rect 452068 43948 480260 43976
rect 452068 43936 452074 43948
rect 480254 43936 480260 43948
rect 480312 43936 480318 43988
rect 481082 43936 481088 43988
rect 481140 43936 481146 43988
rect 509234 43976 509240 43988
rect 481192 43948 509240 43976
rect 452102 43908 452108 43920
rect 451936 43880 452108 43908
rect 452102 43868 452108 43880
rect 452160 43868 452166 43920
rect 452194 43868 452200 43920
rect 452252 43908 452258 43920
rect 480438 43908 480444 43920
rect 452252 43880 480444 43908
rect 452252 43868 452258 43880
rect 480438 43868 480444 43880
rect 480496 43868 480502 43920
rect 480990 43868 480996 43920
rect 481048 43908 481054 43920
rect 481192 43908 481220 43948
rect 509234 43936 509240 43948
rect 509292 43936 509298 43988
rect 510062 43936 510068 43988
rect 510120 43976 510126 43988
rect 538306 43976 538312 43988
rect 510120 43948 538312 43976
rect 510120 43936 510126 43948
rect 538306 43936 538312 43948
rect 538364 43936 538370 43988
rect 538950 43936 538956 43988
rect 539008 43976 539014 43988
rect 567194 43976 567200 43988
rect 539008 43948 567200 43976
rect 539008 43936 539014 43948
rect 567194 43936 567200 43948
rect 567252 43936 567258 43988
rect 481048 43880 481220 43908
rect 481048 43868 481054 43880
rect 481266 43868 481272 43920
rect 481324 43908 481330 43920
rect 509418 43908 509424 43920
rect 481324 43880 509424 43908
rect 481324 43868 481330 43880
rect 509418 43868 509424 43880
rect 509476 43868 509482 43920
rect 510154 43868 510160 43920
rect 510212 43908 510218 43920
rect 538398 43908 538404 43920
rect 510212 43880 538404 43908
rect 510212 43868 510218 43880
rect 538398 43868 538404 43880
rect 538456 43868 538462 43920
rect 539042 43868 539048 43920
rect 539100 43908 539106 43920
rect 567654 43908 567660 43920
rect 539100 43880 567660 43908
rect 539100 43868 539106 43880
rect 567654 43868 567660 43880
rect 567712 43868 567718 43920
rect 539134 43800 539140 43852
rect 539192 43840 539198 43852
rect 567562 43840 567568 43852
rect 539192 43812 567568 43840
rect 539192 43800 539198 43812
rect 567562 43800 567568 43812
rect 567620 43800 567626 43852
rect 32122 40672 32128 40724
rect 32180 40712 32186 40724
rect 219434 40712 219440 40724
rect 32180 40684 219440 40712
rect 32180 40672 32186 40684
rect 219434 40672 219440 40684
rect 219492 40672 219498 40724
rect 538122 40672 538128 40724
rect 538180 40712 538186 40724
rect 567286 40712 567292 40724
rect 538180 40684 567292 40712
rect 538180 40672 538186 40684
rect 567286 40672 567292 40684
rect 567344 40672 567350 40724
rect 536558 39516 536564 39568
rect 536616 39556 536622 39568
rect 567378 39556 567384 39568
rect 536616 39528 567384 39556
rect 536616 39516 536622 39528
rect 567378 39516 567384 39528
rect 567436 39516 567442 39568
rect 536742 39380 536748 39432
rect 536800 39420 536806 39432
rect 567746 39420 567752 39432
rect 536800 39392 567752 39420
rect 536800 39380 536806 39392
rect 567746 39380 567752 39392
rect 567804 39380 567810 39432
rect 536650 39312 536656 39364
rect 536708 39352 536714 39364
rect 567470 39352 567476 39364
rect 536708 39324 567476 39352
rect 536708 39312 536714 39324
rect 567470 39312 567476 39324
rect 567528 39312 567534 39364
rect 71406 39108 71412 39160
rect 71464 39148 71470 39160
rect 100018 39148 100024 39160
rect 71464 39120 100024 39148
rect 71464 39108 71470 39120
rect 100018 39108 100024 39120
rect 100076 39108 100082 39160
rect 100386 39108 100392 39160
rect 100444 39148 100450 39160
rect 128998 39148 129004 39160
rect 100444 39120 129004 39148
rect 100444 39108 100450 39120
rect 128998 39108 129004 39120
rect 129056 39108 129062 39160
rect 129642 39108 129648 39160
rect 129700 39148 129706 39160
rect 157978 39148 157984 39160
rect 129700 39120 157984 39148
rect 129700 39108 129706 39120
rect 157978 39108 157984 39120
rect 158036 39108 158042 39160
rect 158622 39108 158628 39160
rect 158680 39148 158686 39160
rect 186958 39148 186964 39160
rect 158680 39120 186964 39148
rect 158680 39108 158686 39120
rect 186958 39108 186964 39120
rect 187016 39108 187022 39160
rect 187602 39108 187608 39160
rect 187660 39148 187666 39160
rect 215938 39148 215944 39160
rect 187660 39120 215944 39148
rect 187660 39108 187666 39120
rect 215938 39108 215944 39120
rect 215996 39108 216002 39160
rect 216582 39108 216588 39160
rect 216640 39148 216646 39160
rect 246298 39148 246304 39160
rect 216640 39120 246304 39148
rect 216640 39108 216646 39120
rect 246298 39108 246304 39120
rect 246356 39108 246362 39160
rect 246942 39108 246948 39160
rect 247000 39148 247006 39160
rect 275278 39148 275284 39160
rect 247000 39120 275284 39148
rect 247000 39108 247006 39120
rect 275278 39108 275284 39120
rect 275336 39108 275342 39160
rect 275922 39108 275928 39160
rect 275980 39148 275986 39160
rect 304258 39148 304264 39160
rect 275980 39120 304264 39148
rect 275980 39108 275986 39120
rect 304258 39108 304264 39120
rect 304316 39108 304322 39160
rect 304902 39108 304908 39160
rect 304960 39148 304966 39160
rect 333238 39148 333244 39160
rect 304960 39120 333244 39148
rect 304960 39108 304966 39120
rect 333238 39108 333244 39120
rect 333296 39108 333302 39160
rect 333882 39108 333888 39160
rect 333940 39148 333946 39160
rect 362218 39148 362224 39160
rect 333940 39120 362224 39148
rect 333940 39108 333946 39120
rect 362218 39108 362224 39120
rect 362276 39108 362282 39160
rect 362862 39108 362868 39160
rect 362920 39148 362926 39160
rect 391198 39148 391204 39160
rect 362920 39120 391204 39148
rect 362920 39108 362926 39120
rect 391198 39108 391204 39120
rect 391256 39108 391262 39160
rect 391842 39108 391848 39160
rect 391900 39148 391906 39160
rect 420178 39148 420184 39160
rect 391900 39120 420184 39148
rect 391900 39108 391906 39120
rect 420178 39108 420184 39120
rect 420236 39108 420242 39160
rect 420822 39108 420828 39160
rect 420880 39148 420886 39160
rect 449158 39148 449164 39160
rect 420880 39120 449164 39148
rect 420880 39108 420886 39120
rect 449158 39108 449164 39120
rect 449216 39108 449222 39160
rect 449802 39108 449808 39160
rect 449860 39148 449866 39160
rect 478138 39148 478144 39160
rect 449860 39120 478144 39148
rect 449860 39108 449866 39120
rect 478138 39108 478144 39120
rect 478196 39108 478202 39160
rect 478782 39108 478788 39160
rect 478840 39148 478846 39160
rect 507118 39148 507124 39160
rect 478840 39120 507124 39148
rect 478840 39108 478846 39120
rect 507118 39108 507124 39120
rect 507176 39108 507182 39160
rect 507762 39108 507768 39160
rect 507820 39148 507826 39160
rect 536098 39148 536104 39160
rect 507820 39120 536104 39148
rect 507820 39108 507826 39120
rect 536098 39108 536104 39120
rect 536156 39108 536162 39160
rect 71498 39040 71504 39092
rect 71556 39080 71562 39092
rect 100110 39080 100116 39092
rect 71556 39052 100116 39080
rect 71556 39040 71562 39052
rect 100110 39040 100116 39052
rect 100168 39040 100174 39092
rect 100478 39040 100484 39092
rect 100536 39080 100542 39092
rect 129090 39080 129096 39092
rect 100536 39052 129096 39080
rect 100536 39040 100542 39052
rect 129090 39040 129096 39052
rect 129148 39040 129154 39092
rect 129458 39040 129464 39092
rect 129516 39080 129522 39092
rect 158070 39080 158076 39092
rect 129516 39052 158076 39080
rect 129516 39040 129522 39052
rect 158070 39040 158076 39052
rect 158128 39040 158134 39092
rect 158438 39040 158444 39092
rect 158496 39080 158502 39092
rect 187050 39080 187056 39092
rect 158496 39052 187056 39080
rect 158496 39040 158502 39052
rect 187050 39040 187056 39052
rect 187108 39040 187114 39092
rect 187418 39040 187424 39092
rect 187476 39080 187482 39092
rect 216030 39080 216036 39092
rect 187476 39052 216036 39080
rect 187476 39040 187482 39052
rect 216030 39040 216036 39052
rect 216088 39040 216094 39092
rect 216398 39040 216404 39092
rect 216456 39080 216462 39092
rect 246390 39080 246396 39092
rect 216456 39052 246396 39080
rect 216456 39040 216462 39052
rect 246390 39040 246396 39052
rect 246448 39040 246454 39092
rect 246758 39040 246764 39092
rect 246816 39080 246822 39092
rect 275370 39080 275376 39092
rect 246816 39052 275376 39080
rect 246816 39040 246822 39052
rect 275370 39040 275376 39052
rect 275428 39040 275434 39092
rect 275738 39040 275744 39092
rect 275796 39080 275802 39092
rect 304350 39080 304356 39092
rect 275796 39052 304356 39080
rect 275796 39040 275802 39052
rect 304350 39040 304356 39052
rect 304408 39040 304414 39092
rect 304718 39040 304724 39092
rect 304776 39080 304782 39092
rect 333330 39080 333336 39092
rect 304776 39052 333336 39080
rect 304776 39040 304782 39052
rect 333330 39040 333336 39052
rect 333388 39040 333394 39092
rect 333698 39040 333704 39092
rect 333756 39080 333762 39092
rect 362310 39080 362316 39092
rect 333756 39052 362316 39080
rect 333756 39040 333762 39052
rect 362310 39040 362316 39052
rect 362368 39040 362374 39092
rect 362678 39040 362684 39092
rect 362736 39080 362742 39092
rect 391290 39080 391296 39092
rect 362736 39052 391296 39080
rect 362736 39040 362742 39052
rect 391290 39040 391296 39052
rect 391348 39040 391354 39092
rect 391658 39040 391664 39092
rect 391716 39080 391722 39092
rect 420270 39080 420276 39092
rect 391716 39052 420276 39080
rect 391716 39040 391722 39052
rect 420270 39040 420276 39052
rect 420328 39040 420334 39092
rect 420638 39040 420644 39092
rect 420696 39080 420702 39092
rect 449250 39080 449256 39092
rect 420696 39052 449256 39080
rect 420696 39040 420702 39052
rect 449250 39040 449256 39052
rect 449308 39040 449314 39092
rect 449618 39040 449624 39092
rect 449676 39080 449682 39092
rect 478230 39080 478236 39092
rect 449676 39052 478236 39080
rect 449676 39040 449682 39052
rect 478230 39040 478236 39052
rect 478288 39040 478294 39092
rect 478598 39040 478604 39092
rect 478656 39080 478662 39092
rect 507210 39080 507216 39092
rect 478656 39052 507216 39080
rect 478656 39040 478662 39052
rect 507210 39040 507216 39052
rect 507268 39040 507274 39092
rect 507578 39040 507584 39092
rect 507636 39080 507642 39092
rect 536190 39080 536196 39092
rect 507636 39052 536196 39080
rect 507636 39040 507642 39052
rect 536190 39040 536196 39052
rect 536248 39040 536254 39092
rect 28902 38972 28908 39024
rect 28960 39012 28966 39024
rect 580166 39012 580172 39024
rect 28960 38984 580172 39012
rect 28960 38972 28966 38984
rect 580166 38972 580172 38984
rect 580224 38972 580230 39024
rect 8938 38156 8944 38208
rect 8996 38196 9002 38208
rect 22462 38196 22468 38208
rect 8996 38168 22468 38196
rect 8996 38156 9002 38168
rect 22462 38156 22468 38168
rect 22520 38156 22526 38208
rect 11698 38088 11704 38140
rect 11756 38128 11762 38140
rect 30190 38128 30196 38140
rect 11756 38100 30196 38128
rect 11756 38088 11762 38100
rect 30190 38088 30196 38100
rect 30248 38088 30254 38140
rect 4798 38020 4804 38072
rect 4856 38060 4862 38072
rect 19886 38060 19892 38072
rect 4856 38032 19892 38060
rect 4856 38020 4862 38032
rect 19886 38020 19892 38032
rect 19944 38020 19950 38072
rect 19978 38020 19984 38072
rect 20036 38060 20042 38072
rect 41782 38060 41788 38072
rect 20036 38032 41788 38060
rect 20036 38020 20042 38032
rect 41782 38020 41788 38032
rect 41840 38020 41846 38072
rect 3694 37952 3700 38004
rect 3752 37992 3758 38004
rect 38562 37992 38568 38004
rect 3752 37964 38568 37992
rect 3752 37952 3758 37964
rect 38562 37952 38568 37964
rect 38620 37952 38626 38004
rect 3786 37884 3792 37936
rect 3844 37924 3850 37936
rect 45002 37924 45008 37936
rect 3844 37896 45008 37924
rect 3844 37884 3850 37896
rect 45002 37884 45008 37896
rect 45060 37884 45066 37936
rect 29638 37340 29644 37392
rect 29696 37380 29702 37392
rect 33410 37380 33416 37392
rect 29696 37352 33416 37380
rect 29696 37340 29702 37352
rect 33410 37340 33416 37352
rect 33468 37340 33474 37392
rect 40034 37340 40040 37392
rect 40092 37380 40098 37392
rect 48222 37380 48228 37392
rect 40092 37352 48228 37380
rect 40092 37340 40098 37352
rect 48222 37340 48228 37352
rect 48280 37340 48286 37392
rect 61470 37380 61476 37392
rect 55186 37352 61476 37380
rect 36630 37272 36636 37324
rect 36688 37312 36694 37324
rect 55186 37312 55214 37352
rect 61470 37340 61476 37352
rect 61528 37340 61534 37392
rect 36688 37284 55214 37312
rect 36688 37272 36694 37284
rect 56594 37272 56600 37324
rect 56652 37312 56658 37324
rect 61378 37312 61384 37324
rect 56652 37284 61384 37312
rect 56652 37272 56658 37284
rect 61378 37272 61384 37284
rect 61436 37272 61442 37324
rect 9122 34416 9128 34468
rect 9180 34456 9186 34468
rect 12434 34456 12440 34468
rect 9180 34428 12440 34456
rect 9180 34416 9186 34428
rect 12434 34416 12440 34428
rect 12492 34416 12498 34468
rect 3326 31696 3332 31748
rect 3384 31736 3390 31748
rect 12434 31736 12440 31748
rect 3384 31708 12440 31736
rect 3384 31696 3390 31708
rect 12434 31696 12440 31708
rect 12492 31696 12498 31748
rect 63494 27344 63500 27396
rect 63552 27384 63558 27396
rect 65518 27384 65524 27396
rect 63552 27356 65524 27384
rect 63552 27344 63558 27356
rect 65518 27344 65524 27356
rect 65576 27344 65582 27396
rect 4890 23400 4896 23452
rect 4948 23440 4954 23452
rect 12434 23440 12440 23452
rect 4948 23412 12440 23440
rect 4948 23400 4954 23412
rect 12434 23400 12440 23412
rect 12492 23400 12498 23452
rect 7558 22040 7564 22092
rect 7616 22080 7622 22092
rect 12434 22080 12440 22092
rect 7616 22052 12440 22080
rect 7616 22040 7622 22052
rect 12434 22040 12440 22052
rect 12492 22040 12498 22092
rect 61470 20612 61476 20664
rect 61528 20652 61534 20664
rect 70394 20652 70400 20664
rect 61528 20624 70400 20652
rect 61528 20612 61534 20624
rect 70394 20612 70400 20624
rect 70452 20612 70458 20664
rect 9030 17892 9036 17944
rect 9088 17932 9094 17944
rect 12434 17932 12440 17944
rect 9088 17904 12440 17932
rect 9088 17892 9094 17904
rect 12434 17892 12440 17904
rect 12492 17892 12498 17944
rect 61378 17892 61384 17944
rect 61436 17932 61442 17944
rect 70394 17932 70400 17944
rect 61436 17904 70400 17932
rect 61436 17892 61442 17904
rect 70394 17892 70400 17904
rect 70452 17892 70458 17944
rect 3694 16532 3700 16584
rect 3752 16572 3758 16584
rect 63494 16572 63500 16584
rect 3752 16544 63500 16572
rect 3752 16532 3758 16544
rect 63494 16532 63500 16544
rect 63552 16532 63558 16584
rect 71682 16532 71688 16584
rect 71740 16572 71746 16584
rect 99834 16572 99840 16584
rect 71740 16544 99840 16572
rect 71740 16532 71746 16544
rect 99834 16532 99840 16544
rect 99892 16532 99898 16584
rect 100570 16532 100576 16584
rect 100628 16572 100634 16584
rect 128998 16572 129004 16584
rect 100628 16544 129004 16572
rect 100628 16532 100634 16544
rect 128998 16532 129004 16544
rect 129056 16532 129062 16584
rect 129550 16532 129556 16584
rect 129608 16572 129614 16584
rect 157978 16572 157984 16584
rect 129608 16544 157984 16572
rect 129608 16532 129614 16544
rect 157978 16532 157984 16544
rect 158036 16532 158042 16584
rect 158530 16532 158536 16584
rect 158588 16572 158594 16584
rect 186958 16572 186964 16584
rect 158588 16544 186964 16572
rect 158588 16532 158594 16544
rect 186958 16532 186964 16544
rect 187016 16532 187022 16584
rect 187326 16532 187332 16584
rect 187384 16572 187390 16584
rect 215754 16572 215760 16584
rect 187384 16544 215760 16572
rect 187384 16532 187390 16544
rect 215754 16532 215760 16544
rect 215812 16532 215818 16584
rect 216306 16532 216312 16584
rect 216364 16572 216370 16584
rect 245654 16572 245660 16584
rect 216364 16544 245660 16572
rect 216364 16532 216370 16544
rect 245654 16532 245660 16544
rect 245712 16532 245718 16584
rect 246850 16532 246856 16584
rect 246908 16572 246914 16584
rect 275278 16572 275284 16584
rect 246908 16544 275284 16572
rect 246908 16532 246914 16544
rect 275278 16532 275284 16544
rect 275336 16532 275342 16584
rect 275830 16532 275836 16584
rect 275888 16572 275894 16584
rect 304258 16572 304264 16584
rect 275888 16544 304264 16572
rect 275888 16532 275894 16544
rect 304258 16532 304264 16544
rect 304316 16532 304322 16584
rect 304626 16532 304632 16584
rect 304684 16572 304690 16584
rect 332594 16572 332600 16584
rect 304684 16544 332600 16572
rect 304684 16532 304690 16544
rect 332594 16532 332600 16544
rect 332652 16532 332658 16584
rect 333606 16532 333612 16584
rect 333664 16572 333670 16584
rect 361574 16572 361580 16584
rect 333664 16544 361580 16572
rect 333664 16532 333670 16544
rect 361574 16532 361580 16544
rect 361632 16532 361638 16584
rect 362586 16532 362592 16584
rect 362644 16572 362650 16584
rect 390554 16572 390560 16584
rect 362644 16544 390560 16572
rect 362644 16532 362650 16544
rect 390554 16532 390560 16544
rect 390612 16532 390618 16584
rect 391750 16532 391756 16584
rect 391808 16572 391814 16584
rect 420178 16572 420184 16584
rect 391808 16544 420184 16572
rect 391808 16532 391814 16544
rect 420178 16532 420184 16544
rect 420236 16532 420242 16584
rect 420730 16532 420736 16584
rect 420788 16572 420794 16584
rect 449158 16572 449164 16584
rect 420788 16544 449164 16572
rect 420788 16532 420794 16544
rect 449158 16532 449164 16544
rect 449216 16532 449222 16584
rect 449710 16532 449716 16584
rect 449768 16572 449774 16584
rect 478138 16572 478144 16584
rect 449768 16544 478144 16572
rect 449768 16532 449774 16544
rect 478138 16532 478144 16544
rect 478196 16532 478202 16584
rect 478506 16532 478512 16584
rect 478564 16572 478570 16584
rect 506474 16572 506480 16584
rect 478564 16544 506480 16572
rect 478564 16532 478570 16544
rect 506474 16532 506480 16544
rect 506532 16532 506538 16584
rect 507670 16532 507676 16584
rect 507728 16572 507734 16584
rect 536098 16572 536104 16584
rect 507728 16544 536104 16572
rect 507728 16532 507734 16544
rect 536098 16532 536104 16544
rect 536156 16532 536162 16584
rect 13630 16464 13636 16516
rect 13688 16504 13694 16516
rect 71130 16504 71136 16516
rect 13688 16476 71136 16504
rect 13688 16464 13694 16476
rect 71130 16464 71136 16476
rect 71188 16464 71194 16516
rect 71590 16464 71596 16516
rect 71648 16504 71654 16516
rect 100018 16504 100024 16516
rect 71648 16476 100024 16504
rect 71648 16464 71654 16476
rect 100018 16464 100024 16476
rect 100076 16464 100082 16516
rect 100662 16464 100668 16516
rect 100720 16504 100726 16516
rect 128814 16504 128820 16516
rect 100720 16476 128820 16504
rect 100720 16464 100726 16476
rect 128814 16464 128820 16476
rect 128872 16464 128878 16516
rect 129366 16464 129372 16516
rect 129424 16504 129430 16516
rect 157518 16504 157524 16516
rect 129424 16476 157524 16504
rect 129424 16464 129430 16476
rect 157518 16464 157524 16476
rect 157576 16464 157582 16516
rect 158346 16464 158352 16516
rect 158404 16504 158410 16516
rect 186774 16504 186780 16516
rect 158404 16476 186780 16504
rect 158404 16464 158410 16476
rect 186774 16464 186780 16476
rect 186832 16464 186838 16516
rect 187510 16464 187516 16516
rect 187568 16504 187574 16516
rect 215938 16504 215944 16516
rect 187568 16476 215944 16504
rect 187568 16464 187574 16476
rect 215938 16464 215944 16476
rect 215996 16464 216002 16516
rect 216490 16464 216496 16516
rect 216548 16504 216554 16516
rect 246298 16504 246304 16516
rect 216548 16476 246304 16504
rect 216548 16464 216554 16476
rect 246298 16464 246304 16476
rect 246356 16464 246362 16516
rect 246666 16464 246672 16516
rect 246724 16504 246730 16516
rect 274634 16504 274640 16516
rect 246724 16476 274640 16504
rect 246724 16464 246730 16476
rect 274634 16464 274640 16476
rect 274692 16464 274698 16516
rect 275646 16464 275652 16516
rect 275704 16504 275710 16516
rect 303614 16504 303620 16516
rect 275704 16476 303620 16504
rect 275704 16464 275710 16476
rect 303614 16464 303620 16476
rect 303672 16464 303678 16516
rect 304810 16464 304816 16516
rect 304868 16504 304874 16516
rect 333238 16504 333244 16516
rect 304868 16476 333244 16504
rect 304868 16464 304874 16476
rect 333238 16464 333244 16476
rect 333296 16464 333302 16516
rect 333790 16464 333796 16516
rect 333848 16504 333854 16516
rect 362218 16504 362224 16516
rect 333848 16476 362224 16504
rect 333848 16464 333854 16476
rect 362218 16464 362224 16476
rect 362276 16464 362282 16516
rect 362770 16464 362776 16516
rect 362828 16504 362834 16516
rect 391198 16504 391204 16516
rect 362828 16476 391204 16504
rect 362828 16464 362834 16476
rect 391198 16464 391204 16476
rect 391256 16464 391262 16516
rect 391566 16464 391572 16516
rect 391624 16504 391630 16516
rect 419534 16504 419540 16516
rect 391624 16476 419540 16504
rect 391624 16464 391630 16476
rect 419534 16464 419540 16476
rect 419592 16464 419598 16516
rect 420546 16464 420552 16516
rect 420604 16504 420610 16516
rect 448514 16504 448520 16516
rect 420604 16476 448520 16504
rect 420604 16464 420610 16476
rect 448514 16464 448520 16476
rect 448572 16464 448578 16516
rect 449526 16464 449532 16516
rect 449584 16504 449590 16516
rect 477494 16504 477500 16516
rect 449584 16476 477500 16504
rect 449584 16464 449590 16476
rect 477494 16464 477500 16476
rect 477552 16464 477558 16516
rect 478690 16464 478696 16516
rect 478748 16504 478754 16516
rect 507118 16504 507124 16516
rect 478748 16476 507124 16504
rect 478748 16464 478754 16476
rect 507118 16464 507124 16476
rect 507176 16464 507182 16516
rect 507486 16464 507492 16516
rect 507544 16504 507550 16516
rect 535454 16504 535460 16516
rect 507544 16476 535460 16504
rect 507544 16464 507550 16476
rect 535454 16464 535460 16476
rect 535512 16464 535518 16516
rect 38562 15104 38568 15156
rect 38620 15144 38626 15156
rect 71038 15144 71044 15156
rect 38620 15116 71044 15144
rect 38620 15104 38626 15116
rect 71038 15104 71044 15116
rect 71096 15104 71102 15156
rect 4062 13744 4068 13796
rect 4120 13784 4126 13796
rect 16022 13784 16028 13796
rect 4120 13756 16028 13784
rect 4120 13744 4126 13756
rect 16022 13744 16028 13756
rect 16080 13744 16086 13796
rect 17310 13744 17316 13796
rect 17368 13784 17374 13796
rect 580718 13784 580724 13796
rect 17368 13756 580724 13784
rect 17368 13744 17374 13756
rect 580718 13744 580724 13756
rect 580776 13744 580782 13796
rect 20530 13676 20536 13728
rect 20588 13716 20594 13728
rect 580810 13716 580816 13728
rect 20588 13688 580816 13716
rect 20588 13676 20594 13688
rect 580810 13676 580816 13688
rect 580868 13676 580874 13728
rect 3418 13608 3424 13660
rect 3476 13648 3482 13660
rect 30190 13648 30196 13660
rect 3476 13620 30196 13648
rect 3476 13608 3482 13620
rect 30190 13608 30196 13620
rect 30248 13608 30254 13660
rect 32122 13608 32128 13660
rect 32180 13648 32186 13660
rect 580902 13648 580908 13660
rect 32180 13620 580908 13648
rect 32180 13608 32186 13620
rect 580902 13608 580908 13620
rect 580960 13608 580966 13660
rect 6178 13540 6184 13592
rect 6236 13580 6242 13592
rect 28902 13580 28908 13592
rect 6236 13552 28908 13580
rect 6236 13540 6242 13552
rect 28902 13540 28908 13552
rect 28960 13540 28966 13592
rect 36630 13540 36636 13592
rect 36688 13580 36694 13592
rect 580534 13580 580540 13592
rect 36688 13552 580540 13580
rect 36688 13540 36694 13552
rect 580534 13540 580540 13552
rect 580592 13540 580598 13592
rect 3970 13472 3976 13524
rect 4028 13512 4034 13524
rect 25682 13512 25688 13524
rect 4028 13484 25688 13512
rect 4028 13472 4034 13484
rect 25682 13472 25688 13484
rect 25740 13472 25746 13524
rect 43070 13472 43076 13524
rect 43128 13512 43134 13524
rect 580626 13512 580632 13524
rect 43128 13484 580632 13512
rect 43128 13472 43134 13484
rect 580626 13472 580632 13484
rect 580684 13472 580690 13524
rect 3878 13404 3884 13456
rect 3936 13444 3942 13456
rect 22462 13444 22468 13456
rect 3936 13416 22468 13444
rect 3936 13404 3942 13416
rect 22462 13404 22468 13416
rect 22520 13404 22526 13456
rect 45002 13404 45008 13456
rect 45060 13444 45066 13456
rect 580350 13444 580356 13456
rect 45060 13416 580356 13444
rect 45060 13404 45066 13416
rect 580350 13404 580356 13416
rect 580408 13404 580414 13456
rect 3510 13336 3516 13388
rect 3568 13376 3574 13388
rect 54662 13376 54668 13388
rect 3568 13348 54668 13376
rect 3568 13336 3574 13348
rect 54662 13336 54668 13348
rect 54720 13336 54726 13388
rect 59814 13336 59820 13388
rect 59872 13376 59878 13388
rect 580442 13376 580448 13388
rect 59872 13348 580448 13376
rect 59872 13336 59878 13348
rect 580442 13336 580448 13348
rect 580500 13336 580506 13388
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 55950 13308 55956 13320
rect 6972 13280 55956 13308
rect 6972 13268 6978 13280
rect 55950 13268 55956 13280
rect 56008 13268 56014 13320
rect 61102 13268 61108 13320
rect 61160 13308 61166 13320
rect 580258 13308 580264 13320
rect 61160 13280 580264 13308
rect 61160 13268 61166 13280
rect 580258 13268 580264 13280
rect 580316 13268 580322 13320
rect 23750 13200 23756 13252
rect 23808 13240 23814 13252
rect 137002 13240 137008 13252
rect 23808 13212 137008 13240
rect 23808 13200 23814 13212
rect 137002 13200 137008 13212
rect 137060 13200 137066 13252
rect 39850 13132 39856 13184
rect 39908 13172 39914 13184
rect 71774 13172 71780 13184
rect 39908 13144 71780 13172
rect 39908 13132 39914 13144
rect 71774 13132 71780 13144
rect 71832 13132 71838 13184
rect 106 13064 112 13116
rect 164 13104 170 13116
rect 49510 13104 49516 13116
rect 164 13076 49516 13104
rect 164 13064 170 13076
rect 49510 13064 49516 13076
rect 49568 13064 49574 13116
rect 3602 12996 3608 13048
rect 3660 13036 3666 13048
rect 51442 13036 51448 13048
rect 3660 13008 51448 13036
rect 3660 12996 3666 13008
rect 51442 12996 51448 13008
rect 51500 12996 51506 13048
rect 64322 3544 64328 3596
rect 64380 3584 64386 3596
rect 125870 3584 125876 3596
rect 64380 3556 125876 3584
rect 64380 3544 64386 3556
rect 125870 3544 125876 3556
rect 125928 3544 125934 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 33134 3516 33140 3528
rect 1728 3488 33140 3516
rect 1728 3476 1734 3488
rect 33134 3476 33140 3488
rect 33192 3476 33198 3528
rect 64230 3476 64236 3528
rect 64288 3516 64294 3528
rect 126974 3516 126980 3528
rect 64288 3488 126980 3516
rect 64288 3476 64294 3488
rect 126974 3476 126980 3488
rect 127032 3476 127038 3528
rect 13722 3408 13728 3460
rect 13780 3448 13786 3460
rect 129366 3448 129372 3460
rect 13780 3420 129372 3448
rect 13780 3408 13786 3420
rect 129366 3408 129372 3420
rect 129424 3408 129430 3460
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 26240 700816 26292 700868
rect 105452 700816 105504 700868
rect 56600 700748 56652 700800
rect 202788 700748 202840 700800
rect 65524 700680 65576 700732
rect 267648 700680 267700 700732
rect 17960 700612 18012 700664
rect 235172 700612 235224 700664
rect 59360 700544 59412 700596
rect 332508 700544 332560 700596
rect 13728 700476 13780 700528
rect 300124 700476 300176 700528
rect 64144 700408 64196 700460
rect 364984 700408 365036 700460
rect 23480 700340 23532 700392
rect 462320 700340 462372 700392
rect 47032 700272 47084 700324
rect 494796 700272 494848 700324
rect 52460 696940 52512 696992
rect 580172 696940 580224 696992
rect 3424 657432 3476 657484
rect 8944 657432 8996 657484
rect 2780 632068 2832 632120
rect 4804 632068 4856 632120
rect 64236 590656 64288 590708
rect 580172 590656 580224 590708
rect 2964 579640 3016 579692
rect 6184 579640 6236 579692
rect 16580 563048 16632 563100
rect 580172 563048 580224 563100
rect 3424 553392 3476 553444
rect 11704 553392 11756 553444
rect 64328 536800 64380 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 7564 527144 7616 527196
rect 24860 510620 24912 510672
rect 580172 510620 580224 510672
rect 64420 470568 64472 470620
rect 579988 470568 580040 470620
rect 3148 448536 3200 448588
rect 19984 448536 20036 448588
rect 13636 430584 13688 430636
rect 579620 430584 579672 430636
rect 15200 404336 15252 404388
rect 580172 404336 580224 404388
rect 64512 378156 64564 378208
rect 580172 378156 580224 378208
rect 3332 357416 3384 357468
rect 61292 357416 61344 357468
rect 2780 345176 2832 345228
rect 4896 345176 4948 345228
rect 3332 292544 3384 292596
rect 9036 292544 9088 292596
rect 3148 253920 3200 253972
rect 29644 253920 29696 253972
rect 34520 231820 34572 231872
rect 579804 231820 579856 231872
rect 3332 201492 3384 201544
rect 61200 201492 61252 201544
rect 60832 191836 60884 191888
rect 580172 191836 580224 191888
rect 51080 151784 51132 151836
rect 579988 151784 580040 151836
rect 3332 136620 3384 136672
rect 11796 136620 11848 136672
rect 64604 111800 64656 111852
rect 579988 111800 580040 111852
rect 3240 44208 3292 44260
rect 9128 44208 9180 44260
rect 248512 44004 248564 44056
rect 249064 44004 249116 44056
rect 277492 44004 277544 44056
rect 306472 44004 306524 44056
rect 307024 44004 307076 44056
rect 333152 44004 333204 44056
rect 336004 44004 336056 44056
rect 362132 44004 362184 44056
rect 364984 44004 365036 44056
rect 391112 44004 391164 44056
rect 393964 44004 394016 44056
rect 420092 44004 420144 44056
rect 423036 44004 423088 44056
rect 451372 44004 451424 44056
rect 220176 43936 220228 43988
rect 220360 43936 220412 43988
rect 248420 43936 248472 43988
rect 249248 43936 249300 43988
rect 277400 43936 277452 43988
rect 278136 43936 278188 43988
rect 278044 43868 278096 43920
rect 304080 43936 304132 43988
rect 307116 43936 307168 43988
rect 335452 43936 335504 43988
rect 336096 43936 336148 43988
rect 364432 43936 364484 43988
rect 365076 43936 365128 43988
rect 393412 43936 393464 43988
rect 394056 43936 394108 43988
rect 422392 43936 422444 43988
rect 422944 43936 422996 43988
rect 449072 43936 449124 43988
rect 278320 43868 278372 43920
rect 306564 43868 306616 43920
rect 307208 43868 307260 43920
rect 335360 43868 335412 43920
rect 336188 43868 336240 43920
rect 364340 43868 364392 43920
rect 365168 43868 365220 43920
rect 393320 43868 393372 43920
rect 394148 43868 394200 43920
rect 422300 43868 422352 43920
rect 423128 43868 423180 43920
rect 451464 43868 451516 43920
rect 480352 44004 480404 44056
rect 509332 44004 509384 44056
rect 509976 44004 510028 44056
rect 538220 44004 538272 44056
rect 538864 44004 538916 44056
rect 565084 44004 565136 44056
rect 452016 43936 452068 43988
rect 480260 43936 480312 43988
rect 481088 43936 481140 43988
rect 452108 43868 452160 43920
rect 452200 43868 452252 43920
rect 480444 43868 480496 43920
rect 480996 43868 481048 43920
rect 509240 43936 509292 43988
rect 510068 43936 510120 43988
rect 538312 43936 538364 43988
rect 538956 43936 539008 43988
rect 567200 43936 567252 43988
rect 481272 43868 481324 43920
rect 509424 43868 509476 43920
rect 510160 43868 510212 43920
rect 538404 43868 538456 43920
rect 539048 43868 539100 43920
rect 567660 43868 567712 43920
rect 539140 43800 539192 43852
rect 567568 43800 567620 43852
rect 32128 40672 32180 40724
rect 219440 40672 219492 40724
rect 538128 40672 538180 40724
rect 567292 40672 567344 40724
rect 536564 39516 536616 39568
rect 567384 39516 567436 39568
rect 536748 39380 536800 39432
rect 567752 39380 567804 39432
rect 536656 39312 536708 39364
rect 567476 39312 567528 39364
rect 71412 39108 71464 39160
rect 100024 39108 100076 39160
rect 100392 39108 100444 39160
rect 129004 39108 129056 39160
rect 129648 39108 129700 39160
rect 157984 39108 158036 39160
rect 158628 39108 158680 39160
rect 186964 39108 187016 39160
rect 187608 39108 187660 39160
rect 215944 39108 215996 39160
rect 216588 39108 216640 39160
rect 246304 39108 246356 39160
rect 246948 39108 247000 39160
rect 275284 39108 275336 39160
rect 275928 39108 275980 39160
rect 304264 39108 304316 39160
rect 304908 39108 304960 39160
rect 333244 39108 333296 39160
rect 333888 39108 333940 39160
rect 362224 39108 362276 39160
rect 362868 39108 362920 39160
rect 391204 39108 391256 39160
rect 391848 39108 391900 39160
rect 420184 39108 420236 39160
rect 420828 39108 420880 39160
rect 449164 39108 449216 39160
rect 449808 39108 449860 39160
rect 478144 39108 478196 39160
rect 478788 39108 478840 39160
rect 507124 39108 507176 39160
rect 507768 39108 507820 39160
rect 536104 39108 536156 39160
rect 71504 39040 71556 39092
rect 100116 39040 100168 39092
rect 100484 39040 100536 39092
rect 129096 39040 129148 39092
rect 129464 39040 129516 39092
rect 158076 39040 158128 39092
rect 158444 39040 158496 39092
rect 187056 39040 187108 39092
rect 187424 39040 187476 39092
rect 216036 39040 216088 39092
rect 216404 39040 216456 39092
rect 246396 39040 246448 39092
rect 246764 39040 246816 39092
rect 275376 39040 275428 39092
rect 275744 39040 275796 39092
rect 304356 39040 304408 39092
rect 304724 39040 304776 39092
rect 333336 39040 333388 39092
rect 333704 39040 333756 39092
rect 362316 39040 362368 39092
rect 362684 39040 362736 39092
rect 391296 39040 391348 39092
rect 391664 39040 391716 39092
rect 420276 39040 420328 39092
rect 420644 39040 420696 39092
rect 449256 39040 449308 39092
rect 449624 39040 449676 39092
rect 478236 39040 478288 39092
rect 478604 39040 478656 39092
rect 507216 39040 507268 39092
rect 507584 39040 507636 39092
rect 536196 39040 536248 39092
rect 28908 38972 28960 39024
rect 580172 38972 580224 39024
rect 8944 38156 8996 38208
rect 22468 38156 22520 38208
rect 11704 38088 11756 38140
rect 30196 38088 30248 38140
rect 4804 38020 4856 38072
rect 19892 38020 19944 38072
rect 19984 38020 20036 38072
rect 41788 38020 41840 38072
rect 3700 37952 3752 38004
rect 38568 37952 38620 38004
rect 3792 37884 3844 37936
rect 45008 37884 45060 37936
rect 29644 37340 29696 37392
rect 33416 37340 33468 37392
rect 40040 37340 40092 37392
rect 48228 37340 48280 37392
rect 36636 37272 36688 37324
rect 61476 37340 61528 37392
rect 56600 37272 56652 37324
rect 61384 37272 61436 37324
rect 9128 34416 9180 34468
rect 12440 34416 12492 34468
rect 3332 31696 3384 31748
rect 12440 31696 12492 31748
rect 63500 27344 63552 27396
rect 65524 27344 65576 27396
rect 4896 23400 4948 23452
rect 12440 23400 12492 23452
rect 7564 22040 7616 22092
rect 12440 22040 12492 22092
rect 61476 20612 61528 20664
rect 70400 20612 70452 20664
rect 9036 17892 9088 17944
rect 12440 17892 12492 17944
rect 61384 17892 61436 17944
rect 70400 17892 70452 17944
rect 3700 16532 3752 16584
rect 63500 16532 63552 16584
rect 71688 16532 71740 16584
rect 99840 16532 99892 16584
rect 100576 16532 100628 16584
rect 129004 16532 129056 16584
rect 129556 16532 129608 16584
rect 157984 16532 158036 16584
rect 158536 16532 158588 16584
rect 186964 16532 187016 16584
rect 187332 16532 187384 16584
rect 215760 16532 215812 16584
rect 216312 16532 216364 16584
rect 245660 16532 245712 16584
rect 246856 16532 246908 16584
rect 275284 16532 275336 16584
rect 275836 16532 275888 16584
rect 304264 16532 304316 16584
rect 304632 16532 304684 16584
rect 332600 16532 332652 16584
rect 333612 16532 333664 16584
rect 361580 16532 361632 16584
rect 362592 16532 362644 16584
rect 390560 16532 390612 16584
rect 391756 16532 391808 16584
rect 420184 16532 420236 16584
rect 420736 16532 420788 16584
rect 449164 16532 449216 16584
rect 449716 16532 449768 16584
rect 478144 16532 478196 16584
rect 478512 16532 478564 16584
rect 506480 16532 506532 16584
rect 507676 16532 507728 16584
rect 536104 16532 536156 16584
rect 13636 16464 13688 16516
rect 71136 16464 71188 16516
rect 71596 16464 71648 16516
rect 100024 16464 100076 16516
rect 100668 16464 100720 16516
rect 128820 16464 128872 16516
rect 129372 16464 129424 16516
rect 157524 16464 157576 16516
rect 158352 16464 158404 16516
rect 186780 16464 186832 16516
rect 187516 16464 187568 16516
rect 215944 16464 215996 16516
rect 216496 16464 216548 16516
rect 246304 16464 246356 16516
rect 246672 16464 246724 16516
rect 274640 16464 274692 16516
rect 275652 16464 275704 16516
rect 303620 16464 303672 16516
rect 304816 16464 304868 16516
rect 333244 16464 333296 16516
rect 333796 16464 333848 16516
rect 362224 16464 362276 16516
rect 362776 16464 362828 16516
rect 391204 16464 391256 16516
rect 391572 16464 391624 16516
rect 419540 16464 419592 16516
rect 420552 16464 420604 16516
rect 448520 16464 448572 16516
rect 449532 16464 449584 16516
rect 477500 16464 477552 16516
rect 478696 16464 478748 16516
rect 507124 16464 507176 16516
rect 507492 16464 507544 16516
rect 535460 16464 535512 16516
rect 38568 15104 38620 15156
rect 71044 15104 71096 15156
rect 4068 13744 4120 13796
rect 16028 13744 16080 13796
rect 17316 13744 17368 13796
rect 580724 13744 580776 13796
rect 20536 13676 20588 13728
rect 580816 13676 580868 13728
rect 3424 13608 3476 13660
rect 30196 13608 30248 13660
rect 32128 13608 32180 13660
rect 580908 13608 580960 13660
rect 6184 13540 6236 13592
rect 28908 13540 28960 13592
rect 36636 13540 36688 13592
rect 580540 13540 580592 13592
rect 3976 13472 4028 13524
rect 25688 13472 25740 13524
rect 43076 13472 43128 13524
rect 580632 13472 580684 13524
rect 3884 13404 3936 13456
rect 22468 13404 22520 13456
rect 45008 13404 45060 13456
rect 580356 13404 580408 13456
rect 3516 13336 3568 13388
rect 54668 13336 54720 13388
rect 59820 13336 59872 13388
rect 580448 13336 580500 13388
rect 6920 13268 6972 13320
rect 55956 13268 56008 13320
rect 61108 13268 61160 13320
rect 580264 13268 580316 13320
rect 23756 13200 23808 13252
rect 137008 13200 137060 13252
rect 39856 13132 39908 13184
rect 71780 13132 71832 13184
rect 112 13064 164 13116
rect 49516 13064 49568 13116
rect 3608 12996 3660 13048
rect 51448 12996 51500 13048
rect 64328 3544 64380 3596
rect 125876 3544 125928 3596
rect 1676 3476 1728 3528
rect 33140 3476 33192 3528
rect 64236 3476 64288 3528
rect 126980 3476 127032 3528
rect 13728 3408 13780 3460
rect 129372 3408 129424 3460
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 657490 3464 658135
rect 3424 657484 3476 657490
rect 3424 657426 3476 657432
rect 2780 632120 2832 632126
rect 2778 632088 2780 632097
rect 4804 632120 4856 632126
rect 2832 632088 2834 632097
rect 4804 632062 4856 632068
rect 2778 632023 2834 632032
rect 2962 580000 3018 580009
rect 2962 579935 3018 579944
rect 2976 579698 3004 579935
rect 2964 579692 3016 579698
rect 2964 579634 3016 579640
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3344 357474 3372 358391
rect 3332 357468 3384 357474
rect 3332 357410 3384 357416
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 2792 345234 2820 345335
rect 2780 345228 2832 345234
rect 2780 345170 2832 345176
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3344 292602 3372 293111
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3160 253978 3188 254079
rect 3148 253972 3200 253978
rect 3148 253914 3200 253920
rect 3330 201920 3386 201929
rect 3330 201855 3386 201864
rect 3344 201550 3372 201855
rect 3332 201544 3384 201550
rect 3332 201486 3384 201492
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3344 136678 3372 136711
rect 3332 136672 3384 136678
rect 3332 136614 3384 136620
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 3238 45520 3294 45529
rect 3238 45455 3294 45464
rect 3252 44266 3280 45455
rect 3240 44260 3292 44266
rect 3240 44202 3292 44208
rect 3344 31754 3372 58511
rect 3332 31748 3384 31754
rect 3332 31690 3384 31696
rect 3436 13666 3464 410479
rect 3514 397488 3570 397497
rect 3514 397423 3570 397432
rect 3424 13660 3476 13666
rect 3424 13602 3476 13608
rect 3528 13394 3556 397423
rect 3606 306232 3662 306241
rect 3606 306167 3662 306176
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 112 13116 164 13122
rect 112 13058 164 13064
rect 124 354 152 13058
rect 3620 13054 3648 306167
rect 3698 241088 3754 241097
rect 3698 241023 3754 241032
rect 3712 38010 3740 241023
rect 3790 188864 3846 188873
rect 3790 188799 3846 188808
rect 3700 38004 3752 38010
rect 3700 37946 3752 37952
rect 3804 37942 3832 188799
rect 3882 149832 3938 149841
rect 3882 149767 3938 149776
rect 3792 37936 3844 37942
rect 3792 37878 3844 37884
rect 3698 19408 3754 19417
rect 3698 19343 3754 19352
rect 3712 16590 3740 19343
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3896 13462 3924 149767
rect 3974 97608 4030 97617
rect 3974 97543 4030 97552
rect 3988 13530 4016 97543
rect 4066 84688 4122 84697
rect 4066 84623 4122 84632
rect 4080 13802 4108 84623
rect 4816 38078 4844 632062
rect 6184 579692 6236 579698
rect 6184 579634 6236 579640
rect 4896 345228 4948 345234
rect 4896 345170 4948 345176
rect 4804 38072 4856 38078
rect 4804 38014 4856 38020
rect 4908 23458 4936 345170
rect 4896 23452 4948 23458
rect 4896 23394 4948 23400
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 6196 13598 6224 579634
rect 6184 13592 6236 13598
rect 6184 13534 6236 13540
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 3884 13456 3936 13462
rect 3884 13398 3936 13404
rect 6932 13326 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 26240 700868 26292 700874
rect 26240 700810 26292 700816
rect 17960 700664 18012 700670
rect 17960 700606 18012 700612
rect 13728 700528 13780 700534
rect 13728 700470 13780 700476
rect 8944 657484 8996 657490
rect 8944 657426 8996 657432
rect 7564 527196 7616 527202
rect 7564 527138 7616 527144
rect 7576 22098 7604 527138
rect 8956 38214 8984 657426
rect 11704 553444 11756 553450
rect 11704 553386 11756 553392
rect 9036 292596 9088 292602
rect 9036 292538 9088 292544
rect 8944 38208 8996 38214
rect 8944 38150 8996 38156
rect 7564 22092 7616 22098
rect 7564 22034 7616 22040
rect 9048 17950 9076 292538
rect 9128 44260 9180 44266
rect 9128 44202 9180 44208
rect 9140 34474 9168 44202
rect 11716 38146 11744 553386
rect 13636 430636 13688 430642
rect 13636 430578 13688 430584
rect 11796 136672 11848 136678
rect 11796 136614 11848 136620
rect 11704 38140 11756 38146
rect 11704 38082 11756 38088
rect 9128 34468 9180 34474
rect 9128 34410 9180 34416
rect 11808 19553 11836 136614
rect 13542 39400 13598 39409
rect 13542 39335 13598 39344
rect 12438 34504 12494 34513
rect 12438 34439 12440 34448
rect 12492 34439 12494 34448
rect 12440 34410 12492 34416
rect 12440 31748 12492 31754
rect 12440 31690 12492 31696
rect 12452 31113 12480 31690
rect 12438 31104 12494 31113
rect 12438 31039 12494 31048
rect 13556 27713 13584 39335
rect 13648 29753 13676 430578
rect 13740 33153 13768 700470
rect 16580 563100 16632 563106
rect 16580 563042 16632 563048
rect 15200 404388 15252 404394
rect 15200 404330 15252 404336
rect 15212 55214 15240 404330
rect 16592 55214 16620 563042
rect 17972 55214 18000 700606
rect 23480 700392 23532 700398
rect 23480 700334 23532 700340
rect 19984 448588 20036 448594
rect 19984 448530 20036 448536
rect 15212 55186 15608 55214
rect 16592 55186 16896 55214
rect 17972 55186 18920 55214
rect 15580 35986 15608 55186
rect 16868 35986 16896 55186
rect 18892 35986 18920 55186
rect 19996 38078 20024 448530
rect 22468 38208 22520 38214
rect 22468 38150 22520 38156
rect 19892 38072 19944 38078
rect 19892 38014 19944 38020
rect 19984 38072 20036 38078
rect 19984 38014 20036 38020
rect 19904 36122 19932 38014
rect 19904 36094 20208 36122
rect 20180 35986 20208 36094
rect 15580 35958 16054 35986
rect 16868 35958 17342 35986
rect 18892 35958 19274 35986
rect 20180 35958 20562 35986
rect 22480 35972 22508 38150
rect 23492 35986 23520 700334
rect 24860 510672 24912 510678
rect 24860 510614 24912 510620
rect 24872 55214 24900 510614
rect 26252 55214 26280 700810
rect 29644 253972 29696 253978
rect 29644 253914 29696 253920
rect 24872 55186 25360 55214
rect 26252 55186 26648 55214
rect 25332 35986 25360 55186
rect 26620 35986 26648 55186
rect 28908 39024 28960 39030
rect 28908 38966 28960 38972
rect 23492 35958 23782 35986
rect 25332 35958 25714 35986
rect 26620 35958 27002 35986
rect 28920 35972 28948 38966
rect 29656 37398 29684 253914
rect 34520 231872 34572 231878
rect 34520 231814 34572 231820
rect 34532 55214 34560 231814
rect 34532 55186 34928 55214
rect 32128 40724 32180 40730
rect 32128 40666 32180 40672
rect 30196 38140 30248 38146
rect 30196 38082 30248 38088
rect 29644 37392 29696 37398
rect 29644 37334 29696 37340
rect 30208 35972 30236 38082
rect 32140 35972 32168 40666
rect 33416 37392 33468 37398
rect 33416 37334 33468 37340
rect 33428 35972 33456 37334
rect 34900 35986 34928 55186
rect 38568 38004 38620 38010
rect 38568 37946 38620 37952
rect 36636 37324 36688 37330
rect 36636 37266 36688 37272
rect 34900 35958 35374 35986
rect 36648 35972 36676 37266
rect 38580 35972 38608 37946
rect 40052 37398 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137020 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 56600 700800 56652 700806
rect 56600 700742 56652 700748
rect 47032 700324 47084 700330
rect 47032 700266 47084 700272
rect 41788 38072 41840 38078
rect 41788 38014 41840 38020
rect 40040 37392 40092 37398
rect 40040 37334 40092 37340
rect 41800 35972 41828 38014
rect 45008 37936 45060 37942
rect 45008 37878 45060 37884
rect 45020 35972 45048 37878
rect 47044 35986 47072 700266
rect 52460 696992 52512 696998
rect 52460 696934 52512 696940
rect 51080 151836 51132 151842
rect 51080 151778 51132 151784
rect 48228 37392 48280 37398
rect 48228 37334 48280 37340
rect 46966 35958 47072 35986
rect 48240 35972 48268 37334
rect 51092 35986 51120 151778
rect 52472 55214 52500 696934
rect 56612 55214 56640 700742
rect 65524 700732 65576 700738
rect 65524 700674 65576 700680
rect 59360 700596 59412 700602
rect 59360 700538 59412 700544
rect 52472 55186 52960 55214
rect 56612 55186 57560 55214
rect 52932 35986 52960 55186
rect 54666 37904 54722 37913
rect 54666 37839 54722 37848
rect 51092 35958 51474 35986
rect 52932 35958 53406 35986
rect 54680 35972 54708 37839
rect 56600 37324 56652 37330
rect 56600 37266 56652 37272
rect 56612 35972 56640 37266
rect 57532 35986 57560 55186
rect 59372 35986 59400 700538
rect 64144 700460 64196 700466
rect 64144 700402 64196 700408
rect 61292 357468 61344 357474
rect 61292 357410 61344 357416
rect 61200 201544 61252 201550
rect 61200 201486 61252 201492
rect 60832 191888 60884 191894
rect 60832 191830 60884 191836
rect 60844 35986 60872 191830
rect 57532 35958 57914 35986
rect 59372 35958 59846 35986
rect 60844 35958 61134 35986
rect 39670 35320 39726 35329
rect 43442 35320 43498 35329
rect 39726 35278 39882 35306
rect 39670 35255 39726 35264
rect 50526 35320 50582 35329
rect 43498 35278 43746 35306
rect 50186 35278 50526 35306
rect 43442 35255 43498 35264
rect 50526 35255 50582 35264
rect 13726 33144 13782 33153
rect 13726 33079 13782 33088
rect 13634 29744 13690 29753
rect 13634 29679 13690 29688
rect 13542 27704 13598 27713
rect 13542 27639 13598 27648
rect 13634 26344 13690 26353
rect 13634 26279 13690 26288
rect 12440 23452 12492 23458
rect 12440 23394 12492 23400
rect 12452 22953 12480 23394
rect 12438 22944 12494 22953
rect 12438 22879 12494 22888
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12452 20913 12480 22034
rect 12438 20904 12494 20913
rect 12438 20839 12494 20848
rect 11794 19544 11850 19553
rect 11794 19479 11850 19488
rect 9036 17944 9088 17950
rect 9036 17886 9088 17892
rect 12440 17944 12492 17950
rect 12440 17886 12492 17892
rect 12452 17513 12480 17886
rect 12438 17504 12494 17513
rect 12438 17439 12494 17448
rect 13648 16522 13676 26279
rect 61212 26234 61240 201486
rect 61304 34377 61332 357410
rect 61476 37392 61528 37398
rect 61476 37334 61528 37340
rect 61384 37324 61436 37330
rect 61384 37266 61436 37272
rect 61290 34368 61346 34377
rect 61290 34303 61346 34312
rect 61212 26206 61332 26234
rect 13726 24168 13782 24177
rect 13726 24103 13782 24112
rect 13636 16516 13688 16522
rect 13636 16458 13688 16464
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 3608 13048 3660 13054
rect 3608 12990 3660 12996
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1688 480 1716 3470
rect 13740 3466 13768 24103
rect 61304 20641 61332 26206
rect 61290 20632 61346 20641
rect 61290 20567 61346 20576
rect 61396 17950 61424 37266
rect 61488 20670 61516 37334
rect 63500 27396 63552 27402
rect 63500 27338 63552 27344
rect 63512 27033 63540 27338
rect 63498 27024 63554 27033
rect 63498 26959 63554 26968
rect 64156 23633 64184 700402
rect 64236 590708 64288 590714
rect 64236 590650 64288 590656
rect 64248 31657 64276 590650
rect 64328 536852 64380 536858
rect 64328 536794 64380 536800
rect 64234 31648 64290 31657
rect 64234 31583 64290 31592
rect 64234 30288 64290 30297
rect 64234 30223 64290 30232
rect 64142 23624 64198 23633
rect 64142 23559 64198 23568
rect 63498 21448 63554 21457
rect 63498 21383 63554 21392
rect 61476 20664 61528 20670
rect 61476 20606 61528 20612
rect 61384 17944 61436 17950
rect 61384 17886 61436 17892
rect 63512 16590 63540 21383
rect 63500 16584 63552 16590
rect 46018 16552 46074 16561
rect 57610 16552 57666 16561
rect 46074 16510 46322 16538
rect 46018 16487 46074 16496
rect 57666 16510 57914 16538
rect 63500 16526 63552 16532
rect 57610 16487 57666 16496
rect 16040 13802 16068 16116
rect 17328 13802 17356 16116
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 17316 13796 17368 13802
rect 17316 13738 17368 13744
rect 19260 13025 19288 16116
rect 20548 13734 20576 16116
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 22480 13462 22508 16116
rect 22468 13456 22520 13462
rect 22468 13398 22520 13404
rect 23768 13258 23796 16116
rect 25700 13530 25728 16116
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 26988 13297 27016 16116
rect 28920 13598 28948 16116
rect 30208 13666 30236 16116
rect 32140 13666 32168 16116
rect 33152 16102 33442 16130
rect 30196 13660 30248 13666
rect 30196 13602 30248 13608
rect 32128 13660 32180 13666
rect 32128 13602 32180 13608
rect 28908 13592 28960 13598
rect 28908 13534 28960 13540
rect 26974 13288 27030 13297
rect 23756 13252 23808 13258
rect 26974 13223 27030 13232
rect 23756 13194 23808 13200
rect 19246 13016 19302 13025
rect 19246 12951 19302 12960
rect 33152 3534 33180 16102
rect 35360 13569 35388 16116
rect 36648 13598 36676 16116
rect 38580 15162 38608 16116
rect 38568 15156 38620 15162
rect 38568 15098 38620 15104
rect 36636 13592 36688 13598
rect 35346 13560 35402 13569
rect 36636 13534 36688 13540
rect 35346 13495 35402 13504
rect 39868 13190 39896 16116
rect 41800 13433 41828 16116
rect 43088 13530 43116 16116
rect 43076 13524 43128 13530
rect 43076 13466 43128 13472
rect 45020 13462 45048 16116
rect 45008 13456 45060 13462
rect 41786 13424 41842 13433
rect 45008 13398 45060 13404
rect 41786 13359 41842 13368
rect 39856 13184 39908 13190
rect 48240 13161 48268 16116
rect 39856 13126 39908 13132
rect 48226 13152 48282 13161
rect 49528 13122 49556 16116
rect 48226 13087 48282 13096
rect 49516 13116 49568 13122
rect 49516 13058 49568 13064
rect 51460 13054 51488 16116
rect 52748 13569 52776 16116
rect 52734 13560 52790 13569
rect 52734 13495 52790 13504
rect 54680 13394 54708 16116
rect 54668 13388 54720 13394
rect 54668 13330 54720 13336
rect 55968 13326 55996 16116
rect 59832 13394 59860 16116
rect 59820 13388 59872 13394
rect 59820 13330 59872 13336
rect 61120 13326 61148 16116
rect 55956 13320 56008 13326
rect 55956 13262 56008 13268
rect 61108 13320 61160 13326
rect 61108 13262 61160 13268
rect 51448 13048 51500 13054
rect 51448 12990 51500 12996
rect 64248 3534 64276 30223
rect 64340 28393 64368 536794
rect 64420 470620 64472 470626
rect 64420 470562 64472 470568
rect 64326 28384 64382 28393
rect 64326 28319 64382 28328
rect 64326 24984 64382 24993
rect 64326 24919 64382 24928
rect 64340 3602 64368 24919
rect 64432 18193 64460 470562
rect 64512 378208 64564 378214
rect 64512 378150 64564 378156
rect 64524 35193 64552 378150
rect 64604 111852 64656 111858
rect 64604 111794 64656 111800
rect 64510 35184 64566 35193
rect 64510 35119 64566 35128
rect 64418 18184 64474 18193
rect 64418 18119 64474 18128
rect 64616 16833 64644 111794
rect 65536 27402 65564 700674
rect 71412 39160 71464 39166
rect 71412 39102 71464 39108
rect 71424 32473 71452 39102
rect 71504 39092 71556 39098
rect 71504 39034 71556 39040
rect 71410 32464 71466 32473
rect 71410 32399 71466 32408
rect 71516 29481 71544 39034
rect 71686 38448 71742 38457
rect 71686 38383 71742 38392
rect 71594 35456 71650 35465
rect 71594 35391 71650 35400
rect 71502 29472 71558 29481
rect 71502 29407 71558 29416
rect 65524 27396 65576 27402
rect 65524 27338 65576 27344
rect 71042 26480 71098 26489
rect 71042 26415 71098 26424
rect 70400 20664 70452 20670
rect 70400 20606 70452 20612
rect 70412 20505 70440 20606
rect 70398 20496 70454 20505
rect 70398 20431 70454 20440
rect 70400 17944 70452 17950
rect 70400 17886 70452 17892
rect 70412 17513 70440 17886
rect 70398 17504 70454 17513
rect 70398 17439 70454 17448
rect 64602 16824 64658 16833
rect 64602 16759 64658 16768
rect 71056 15162 71084 26415
rect 71134 23488 71190 23497
rect 71134 23423 71190 23432
rect 71148 16522 71176 23423
rect 71608 16522 71636 35391
rect 71700 16590 71728 38383
rect 71688 16584 71740 16590
rect 71688 16526 71740 16532
rect 71136 16516 71188 16522
rect 71136 16458 71188 16464
rect 71596 16516 71648 16522
rect 71596 16458 71648 16464
rect 71044 15156 71096 15162
rect 71044 15098 71096 15104
rect 71792 13190 71820 702986
rect 105464 700874 105492 703520
rect 105452 700868 105504 700874
rect 105452 700810 105504 700816
rect 100024 39160 100076 39166
rect 100024 39102 100076 39108
rect 100392 39160 100444 39166
rect 100392 39102 100444 39108
rect 129004 39160 129056 39166
rect 129004 39102 129056 39108
rect 129648 39160 129700 39166
rect 129648 39102 129700 39108
rect 100036 23497 100064 39102
rect 100116 39092 100168 39098
rect 100116 39034 100168 39040
rect 100128 26489 100156 39034
rect 100404 32473 100432 39102
rect 100484 39092 100536 39098
rect 100484 39034 100536 39040
rect 100390 32464 100446 32473
rect 100390 32399 100446 32408
rect 100496 29481 100524 39034
rect 100666 38448 100722 38457
rect 100666 38383 100722 38392
rect 100574 35456 100630 35465
rect 100574 35391 100630 35400
rect 100482 29472 100538 29481
rect 100482 29407 100538 29416
rect 100114 26480 100170 26489
rect 100114 26415 100170 26424
rect 100022 23488 100078 23497
rect 100022 23423 100078 23432
rect 100022 20496 100078 20505
rect 100022 20431 100078 20440
rect 99838 17504 99894 17513
rect 99838 17439 99894 17448
rect 99852 16590 99880 17439
rect 99840 16584 99892 16590
rect 99840 16526 99892 16532
rect 100036 16522 100064 20431
rect 100588 16590 100616 35391
rect 100576 16584 100628 16590
rect 100576 16526 100628 16532
rect 100680 16522 100708 38383
rect 129016 23497 129044 39102
rect 129096 39092 129148 39098
rect 129096 39034 129148 39040
rect 129464 39092 129516 39098
rect 129464 39034 129516 39040
rect 129108 26489 129136 39034
rect 129370 38448 129426 38457
rect 129370 38383 129426 38392
rect 129094 26480 129150 26489
rect 129094 26415 129150 26424
rect 129002 23488 129058 23497
rect 129002 23423 129058 23432
rect 129002 20496 129058 20505
rect 129002 20431 129058 20440
rect 128818 17504 128874 17513
rect 128818 17439 128874 17448
rect 128832 16522 128860 17439
rect 129016 16590 129044 20431
rect 129004 16584 129056 16590
rect 129004 16526 129056 16532
rect 129384 16522 129412 38383
rect 129476 29481 129504 39034
rect 129554 35456 129610 35465
rect 129554 35391 129610 35400
rect 129462 29472 129518 29481
rect 129462 29407 129518 29416
rect 129568 16590 129596 35391
rect 129660 32473 129688 39102
rect 129646 32464 129702 32473
rect 129646 32399 129702 32408
rect 129556 16584 129608 16590
rect 129556 16526 129608 16532
rect 100024 16516 100076 16522
rect 100024 16458 100076 16464
rect 100668 16516 100720 16522
rect 100668 16458 100720 16464
rect 128820 16516 128872 16522
rect 128820 16458 128872 16464
rect 129372 16516 129424 16522
rect 129372 16458 129424 16464
rect 137020 13258 137048 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 170324 699825 170352 703520
rect 202800 700806 202828 703520
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 235184 700670 235212 703520
rect 267660 700738 267688 703520
rect 267648 700732 267700 700738
rect 267648 700674 267700 700680
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 300136 700534 300164 703520
rect 332520 700602 332548 703520
rect 332508 700596 332560 700602
rect 332508 700538 332560 700544
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 364996 700466 365024 703520
rect 364984 700460 365036 700466
rect 364984 700402 365036 700408
rect 397472 699825 397500 703520
rect 429856 699825 429884 703520
rect 462332 700398 462360 703520
rect 462320 700392 462372 700398
rect 462320 700334 462372 700340
rect 494808 700330 494836 703520
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 527192 699825 527220 703520
rect 559668 699825 559696 703520
rect 170310 699816 170366 699825
rect 170310 699751 170366 699760
rect 397458 699816 397514 699825
rect 397458 699751 397514 699760
rect 429842 699816 429898 699825
rect 429842 699751 429898 699760
rect 527178 699816 527234 699825
rect 527178 699751 527234 699760
rect 559654 699816 559710 699825
rect 559654 699751 559710 699760
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 590714 580212 590951
rect 580172 590708 580224 590714
rect 580172 590650 580224 590656
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563106 580212 564295
rect 580172 563100 580224 563106
rect 580172 563042 580224 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 579618 431624 579674 431633
rect 579618 431559 579674 431568
rect 579632 430642 579660 431559
rect 579620 430636 579672 430642
rect 579620 430578 579672 430584
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579802 232384 579858 232393
rect 579802 232319 579858 232328
rect 579816 231878 579844 232319
rect 579804 231872 579856 231878
rect 579804 231814 579856 231820
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191894 580212 192471
rect 580172 191888 580224 191894
rect 580172 191830 580224 191836
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 579986 112840 580042 112849
rect 579986 112775 580042 112784
rect 580000 111858 580028 112775
rect 579988 111852 580040 111858
rect 579988 111794 580040 111800
rect 451922 65648 451978 65657
rect 451922 65583 451978 65592
rect 480902 65648 480958 65657
rect 480902 65583 480958 65592
rect 509882 65648 509938 65657
rect 509882 65583 509938 65592
rect 538862 65648 538918 65657
rect 538862 65583 538918 65592
rect 567198 65648 567254 65657
rect 567198 65583 567254 65592
rect 220082 65104 220138 65113
rect 220082 65039 220138 65048
rect 219438 47152 219494 47161
rect 219438 47087 219494 47096
rect 217138 44160 217194 44169
rect 217138 44095 217194 44104
rect 217152 39409 217180 44095
rect 219452 40730 219480 47087
rect 220096 43353 220124 65039
rect 249154 62656 249210 62665
rect 249154 62591 249210 62600
rect 278042 62656 278098 62665
rect 278042 62591 278098 62600
rect 307022 62656 307078 62665
rect 307022 62591 307078 62600
rect 336002 62656 336058 62665
rect 336002 62591 336058 62600
rect 364982 62656 365038 62665
rect 364982 62591 365038 62600
rect 393962 62656 394018 62665
rect 393962 62591 394018 62600
rect 422942 62656 422998 62665
rect 422942 62591 422998 62600
rect 220266 62248 220322 62257
rect 220266 62183 220322 62192
rect 220174 59392 220230 59401
rect 220174 59327 220230 59336
rect 220188 43994 220216 59327
rect 220176 43988 220228 43994
rect 220176 43930 220228 43936
rect 220280 43625 220308 62183
rect 249062 59664 249118 59673
rect 249062 59599 249118 59608
rect 220358 56808 220414 56817
rect 220358 56743 220414 56752
rect 220372 43994 220400 56743
rect 248418 53680 248474 53689
rect 248418 53615 248474 53624
rect 246118 47152 246174 47161
rect 245948 47110 246118 47138
rect 220360 43988 220412 43994
rect 220360 43930 220412 43936
rect 245948 43625 245976 47110
rect 246118 47087 246174 47096
rect 248432 43994 248460 53615
rect 248510 50688 248566 50697
rect 248510 50623 248566 50632
rect 248524 44062 248552 50623
rect 249076 44062 249104 59599
rect 248512 44056 248564 44062
rect 248512 43998 248564 44004
rect 249064 44056 249116 44062
rect 249064 43998 249116 44004
rect 248420 43988 248472 43994
rect 248420 43930 248472 43936
rect 249168 43625 249196 62591
rect 249246 56672 249302 56681
rect 249246 56607 249302 56616
rect 249260 43994 249288 56607
rect 277398 53680 277454 53689
rect 277398 53615 277454 53624
rect 275098 47152 275154 47161
rect 275098 47087 275154 47096
rect 249248 43988 249300 43994
rect 249248 43930 249300 43936
rect 220266 43616 220322 43625
rect 220266 43551 220322 43560
rect 245934 43616 245990 43625
rect 245934 43551 245990 43560
rect 249154 43616 249210 43625
rect 249154 43551 249210 43560
rect 275006 43616 275062 43625
rect 275112 43602 275140 47087
rect 277412 43994 277440 53615
rect 277490 50688 277546 50697
rect 277490 50623 277546 50632
rect 277504 44062 277532 50623
rect 277492 44056 277544 44062
rect 277492 43998 277544 44004
rect 277400 43988 277452 43994
rect 277400 43930 277452 43936
rect 278056 43926 278084 62591
rect 278134 59664 278190 59673
rect 278134 59599 278190 59608
rect 278148 43994 278176 59599
rect 278226 56672 278282 56681
rect 278226 56607 278282 56616
rect 278240 55214 278268 56607
rect 278240 55186 278360 55214
rect 278136 43988 278188 43994
rect 278136 43930 278188 43936
rect 278332 43926 278360 55186
rect 306562 53680 306618 53689
rect 306562 53615 306618 53624
rect 306470 50688 306526 50697
rect 306470 50623 306526 50632
rect 304078 47152 304134 47161
rect 304078 47087 304134 47096
rect 304092 43994 304120 47087
rect 306484 44062 306512 50623
rect 306472 44056 306524 44062
rect 306472 43998 306524 44004
rect 304080 43988 304132 43994
rect 304080 43930 304132 43936
rect 306576 43926 306604 53615
rect 307036 44062 307064 62591
rect 307114 59664 307170 59673
rect 307114 59599 307170 59608
rect 307024 44056 307076 44062
rect 307024 43998 307076 44004
rect 307128 43994 307156 59599
rect 307206 56672 307262 56681
rect 307206 56607 307262 56616
rect 307116 43988 307168 43994
rect 307116 43930 307168 43936
rect 307220 43926 307248 56607
rect 335358 53680 335414 53689
rect 335358 53615 335414 53624
rect 333150 47152 333206 47161
rect 333150 47087 333206 47096
rect 333164 44062 333192 47087
rect 333152 44056 333204 44062
rect 333152 43998 333204 44004
rect 335372 43926 335400 53615
rect 335450 50688 335506 50697
rect 335450 50623 335506 50632
rect 335464 43994 335492 50623
rect 336016 44062 336044 62591
rect 336094 59664 336150 59673
rect 336094 59599 336150 59608
rect 336004 44056 336056 44062
rect 336004 43998 336056 44004
rect 336108 43994 336136 59599
rect 336186 56672 336242 56681
rect 336186 56607 336242 56616
rect 335452 43988 335504 43994
rect 335452 43930 335504 43936
rect 336096 43988 336148 43994
rect 336096 43930 336148 43936
rect 336200 43926 336228 56607
rect 364338 53680 364394 53689
rect 364338 53615 364394 53624
rect 362130 47152 362186 47161
rect 362130 47087 362186 47096
rect 362144 44062 362172 47087
rect 362132 44056 362184 44062
rect 362132 43998 362184 44004
rect 364352 43926 364380 53615
rect 364430 50688 364486 50697
rect 364430 50623 364486 50632
rect 364444 43994 364472 50623
rect 364996 44062 365024 62591
rect 365074 59664 365130 59673
rect 365074 59599 365130 59608
rect 364984 44056 365036 44062
rect 364984 43998 365036 44004
rect 365088 43994 365116 59599
rect 365166 56672 365222 56681
rect 365166 56607 365222 56616
rect 364432 43988 364484 43994
rect 364432 43930 364484 43936
rect 365076 43988 365128 43994
rect 365076 43930 365128 43936
rect 365180 43926 365208 56607
rect 393318 53680 393374 53689
rect 393318 53615 393374 53624
rect 391110 47152 391166 47161
rect 391110 47087 391166 47096
rect 391124 44062 391152 47087
rect 391112 44056 391164 44062
rect 391112 43998 391164 44004
rect 393332 43926 393360 53615
rect 393410 50688 393466 50697
rect 393410 50623 393466 50632
rect 393424 43994 393452 50623
rect 393976 44062 394004 62591
rect 394054 59664 394110 59673
rect 394054 59599 394110 59608
rect 393964 44056 394016 44062
rect 393964 43998 394016 44004
rect 394068 43994 394096 59599
rect 394146 56672 394202 56681
rect 394146 56607 394202 56616
rect 393412 43988 393464 43994
rect 393412 43930 393464 43936
rect 394056 43988 394108 43994
rect 394056 43930 394108 43936
rect 394160 43926 394188 56607
rect 422298 53680 422354 53689
rect 422298 53615 422354 53624
rect 420090 47152 420146 47161
rect 420090 47087 420146 47096
rect 420104 44062 420132 47087
rect 420092 44056 420144 44062
rect 420092 43998 420144 44004
rect 422312 43926 422340 53615
rect 422390 50688 422446 50697
rect 422390 50623 422446 50632
rect 422404 43994 422432 50623
rect 422956 43994 422984 62591
rect 423034 59664 423090 59673
rect 423034 59599 423090 59608
rect 423048 44062 423076 59599
rect 423126 56672 423182 56681
rect 423126 56607 423182 56616
rect 423036 44056 423088 44062
rect 423036 43998 423088 44004
rect 422392 43988 422444 43994
rect 422392 43930 422444 43936
rect 422944 43988 422996 43994
rect 422944 43930 422996 43936
rect 423140 43926 423168 56607
rect 451462 53680 451518 53689
rect 451462 53615 451518 53624
rect 451370 50688 451426 50697
rect 451370 50623 451426 50632
rect 449070 47152 449126 47161
rect 449070 47087 449126 47096
rect 449084 43994 449112 47087
rect 451384 44062 451412 50623
rect 451372 44056 451424 44062
rect 451372 43998 451424 44004
rect 449072 43988 449124 43994
rect 449072 43930 449124 43936
rect 451476 43926 451504 53615
rect 278044 43920 278096 43926
rect 278044 43862 278096 43868
rect 278320 43920 278372 43926
rect 278320 43862 278372 43868
rect 306564 43920 306616 43926
rect 306564 43862 306616 43868
rect 307208 43920 307260 43926
rect 307208 43862 307260 43868
rect 335360 43920 335412 43926
rect 335360 43862 335412 43868
rect 336188 43920 336240 43926
rect 336188 43862 336240 43868
rect 364340 43920 364392 43926
rect 364340 43862 364392 43868
rect 365168 43920 365220 43926
rect 365168 43862 365220 43868
rect 393320 43920 393372 43926
rect 393320 43862 393372 43868
rect 394148 43920 394200 43926
rect 394148 43862 394200 43868
rect 422300 43920 422352 43926
rect 422300 43862 422352 43868
rect 423128 43920 423180 43926
rect 423128 43862 423180 43868
rect 451464 43920 451516 43926
rect 451464 43862 451516 43868
rect 451936 43625 451964 65583
rect 452014 62656 452070 62665
rect 452014 62591 452070 62600
rect 452028 43994 452056 62591
rect 452106 59664 452162 59673
rect 452106 59599 452162 59608
rect 452016 43988 452068 43994
rect 452016 43930 452068 43936
rect 452120 43926 452148 59599
rect 452198 56672 452254 56681
rect 452198 56607 452254 56616
rect 452212 43926 452240 56607
rect 480442 53680 480498 53689
rect 480442 53615 480498 53624
rect 480350 50688 480406 50697
rect 480350 50623 480406 50632
rect 480258 47696 480314 47705
rect 480258 47631 480314 47640
rect 480272 43994 480300 47631
rect 480364 44062 480392 50623
rect 480352 44056 480404 44062
rect 480352 43998 480404 44004
rect 480260 43988 480312 43994
rect 480260 43930 480312 43936
rect 480456 43926 480484 53615
rect 452108 43920 452160 43926
rect 452108 43862 452160 43868
rect 452200 43920 452252 43926
rect 452200 43862 452252 43868
rect 480444 43920 480496 43926
rect 480444 43862 480496 43868
rect 480916 43625 480944 65583
rect 480994 62656 481050 62665
rect 480994 62591 481050 62600
rect 481008 43926 481036 62591
rect 481086 59664 481142 59673
rect 481086 59599 481142 59608
rect 481100 43994 481128 59599
rect 481178 56672 481234 56681
rect 481178 56607 481234 56616
rect 481192 55214 481220 56607
rect 481192 55186 481312 55214
rect 481088 43988 481140 43994
rect 481088 43930 481140 43936
rect 481284 43926 481312 55186
rect 509422 53680 509478 53689
rect 509422 53615 509478 53624
rect 509330 50688 509386 50697
rect 509330 50623 509386 50632
rect 509238 47696 509294 47705
rect 509238 47631 509294 47640
rect 509252 43994 509280 47631
rect 509344 44062 509372 50623
rect 509332 44056 509384 44062
rect 509332 43998 509384 44004
rect 509240 43988 509292 43994
rect 509240 43930 509292 43936
rect 509436 43926 509464 53615
rect 480996 43920 481048 43926
rect 480996 43862 481048 43868
rect 481272 43920 481324 43926
rect 481272 43862 481324 43868
rect 509424 43920 509476 43926
rect 509424 43862 509476 43868
rect 509896 43625 509924 65583
rect 509974 62656 510030 62665
rect 509974 62591 510030 62600
rect 509988 44062 510016 62591
rect 510066 59664 510122 59673
rect 510066 59599 510122 59608
rect 509976 44056 510028 44062
rect 509976 43998 510028 44004
rect 510080 43994 510108 59599
rect 510158 56672 510214 56681
rect 510158 56607 510214 56616
rect 510068 43988 510120 43994
rect 510068 43930 510120 43936
rect 510172 43926 510200 56607
rect 538402 53680 538458 53689
rect 538402 53615 538458 53624
rect 538310 50688 538366 50697
rect 538310 50623 538366 50632
rect 538218 47696 538274 47705
rect 538218 47631 538274 47640
rect 538232 44062 538260 47631
rect 538220 44056 538272 44062
rect 538220 43998 538272 44004
rect 538324 43994 538352 50623
rect 538312 43988 538364 43994
rect 538312 43930 538364 43936
rect 538416 43926 538444 53615
rect 538876 44062 538904 65583
rect 538954 62656 539010 62665
rect 538954 62591 539010 62600
rect 538864 44056 538916 44062
rect 538864 43998 538916 44004
rect 538968 43994 538996 62591
rect 539046 59664 539102 59673
rect 539046 59599 539102 59608
rect 538956 43988 539008 43994
rect 538956 43930 539008 43936
rect 539060 43926 539088 59599
rect 539138 56672 539194 56681
rect 539138 56607 539194 56616
rect 510160 43920 510212 43926
rect 510160 43862 510212 43868
rect 538404 43920 538456 43926
rect 538404 43862 538456 43868
rect 539048 43920 539100 43926
rect 539048 43862 539100 43868
rect 539152 43858 539180 56607
rect 567212 50810 567240 65583
rect 567290 62656 567346 62665
rect 567290 62591 567346 62600
rect 567304 50946 567332 62591
rect 567382 59664 567438 59673
rect 567382 59599 567438 59608
rect 567396 51082 567424 59599
rect 567474 56672 567530 56681
rect 567474 56607 567530 56616
rect 567488 55214 567516 56607
rect 567488 55186 567792 55214
rect 567566 53680 567622 53689
rect 567566 53615 567622 53624
rect 567396 51054 567516 51082
rect 567304 50918 567424 50946
rect 567212 50782 567332 50810
rect 567198 47696 567254 47705
rect 567198 47631 567254 47640
rect 565082 44160 565138 44169
rect 565082 44095 565138 44104
rect 565096 44062 565124 44095
rect 565084 44056 565136 44062
rect 565084 43998 565136 44004
rect 567212 43994 567240 47631
rect 567200 43988 567252 43994
rect 567200 43930 567252 43936
rect 539140 43852 539192 43858
rect 539140 43794 539192 43800
rect 275062 43574 275140 43602
rect 451922 43616 451978 43625
rect 275006 43551 275062 43560
rect 451922 43551 451978 43560
rect 480902 43616 480958 43625
rect 480902 43551 480958 43560
rect 509882 43616 509938 43625
rect 509882 43551 509938 43560
rect 220082 43344 220138 43353
rect 220082 43279 220138 43288
rect 567304 40730 567332 50782
rect 219440 40724 219492 40730
rect 219440 40666 219492 40672
rect 538128 40724 538180 40730
rect 538128 40666 538180 40672
rect 567292 40724 567344 40730
rect 567292 40666 567344 40672
rect 536564 39568 536616 39574
rect 536564 39510 536616 39516
rect 217138 39400 217194 39409
rect 217138 39335 217194 39344
rect 157984 39160 158036 39166
rect 157984 39102 158036 39108
rect 158628 39160 158680 39166
rect 158628 39102 158680 39108
rect 186964 39160 187016 39166
rect 186964 39102 187016 39108
rect 187608 39160 187660 39166
rect 187608 39102 187660 39108
rect 215944 39160 215996 39166
rect 215944 39102 215996 39108
rect 216588 39160 216640 39166
rect 216588 39102 216640 39108
rect 246304 39160 246356 39166
rect 246304 39102 246356 39108
rect 246948 39160 247000 39166
rect 246948 39102 247000 39108
rect 275284 39160 275336 39166
rect 275284 39102 275336 39108
rect 275928 39160 275980 39166
rect 275928 39102 275980 39108
rect 304264 39160 304316 39166
rect 304264 39102 304316 39108
rect 304908 39160 304960 39166
rect 304908 39102 304960 39108
rect 333244 39160 333296 39166
rect 333244 39102 333296 39108
rect 333888 39160 333940 39166
rect 333888 39102 333940 39108
rect 362224 39160 362276 39166
rect 362224 39102 362276 39108
rect 362868 39160 362920 39166
rect 362868 39102 362920 39108
rect 391204 39160 391256 39166
rect 391204 39102 391256 39108
rect 391848 39160 391900 39166
rect 391848 39102 391900 39108
rect 420184 39160 420236 39166
rect 420184 39102 420236 39108
rect 420828 39160 420880 39166
rect 420828 39102 420880 39108
rect 449164 39160 449216 39166
rect 449164 39102 449216 39108
rect 449808 39160 449860 39166
rect 449808 39102 449860 39108
rect 478144 39160 478196 39166
rect 478144 39102 478196 39108
rect 478788 39160 478840 39166
rect 478788 39102 478840 39108
rect 507124 39160 507176 39166
rect 507124 39102 507176 39108
rect 507768 39160 507820 39166
rect 507768 39102 507820 39108
rect 536104 39160 536156 39166
rect 536104 39102 536156 39108
rect 157996 23497 158024 39102
rect 158076 39092 158128 39098
rect 158076 39034 158128 39040
rect 158444 39092 158496 39098
rect 158444 39034 158496 39040
rect 158088 26489 158116 39034
rect 158350 38448 158406 38457
rect 158350 38383 158406 38392
rect 158074 26480 158130 26489
rect 158074 26415 158130 26424
rect 157982 23488 158038 23497
rect 157982 23423 158038 23432
rect 157982 20496 158038 20505
rect 157982 20431 158038 20440
rect 157522 17504 157578 17513
rect 157522 17439 157578 17448
rect 157536 16522 157564 17439
rect 157996 16590 158024 20431
rect 157984 16584 158036 16590
rect 157984 16526 158036 16532
rect 158364 16522 158392 38383
rect 158456 29481 158484 39034
rect 158534 35456 158590 35465
rect 158534 35391 158590 35400
rect 158442 29472 158498 29481
rect 158442 29407 158498 29416
rect 158548 16590 158576 35391
rect 158640 32473 158668 39102
rect 158626 32464 158682 32473
rect 158626 32399 158682 32408
rect 186976 23497 187004 39102
rect 187056 39092 187108 39098
rect 187056 39034 187108 39040
rect 187424 39092 187476 39098
rect 187424 39034 187476 39040
rect 187068 26489 187096 39034
rect 187330 38448 187386 38457
rect 187330 38383 187386 38392
rect 187054 26480 187110 26489
rect 187054 26415 187110 26424
rect 186962 23488 187018 23497
rect 186962 23423 187018 23432
rect 186962 20496 187018 20505
rect 186962 20431 187018 20440
rect 186778 17504 186834 17513
rect 186778 17439 186834 17448
rect 158536 16584 158588 16590
rect 158536 16526 158588 16532
rect 186792 16522 186820 17439
rect 186976 16590 187004 20431
rect 187344 16590 187372 38383
rect 187436 29481 187464 39034
rect 187514 35456 187570 35465
rect 187514 35391 187570 35400
rect 187422 29472 187478 29481
rect 187422 29407 187478 29416
rect 186964 16584 187016 16590
rect 186964 16526 187016 16532
rect 187332 16584 187384 16590
rect 187332 16526 187384 16532
rect 187528 16522 187556 35391
rect 187620 32473 187648 39102
rect 187606 32464 187662 32473
rect 187606 32399 187662 32408
rect 215956 23497 215984 39102
rect 216036 39092 216088 39098
rect 216036 39034 216088 39040
rect 216404 39092 216456 39098
rect 216404 39034 216456 39040
rect 216048 26489 216076 39034
rect 216310 38448 216366 38457
rect 216310 38383 216366 38392
rect 216034 26480 216090 26489
rect 216034 26415 216090 26424
rect 215942 23488 215998 23497
rect 215942 23423 215998 23432
rect 215942 20496 215998 20505
rect 215942 20431 215998 20440
rect 215758 17504 215814 17513
rect 215758 17439 215814 17448
rect 215772 16590 215800 17439
rect 215760 16584 215812 16590
rect 215760 16526 215812 16532
rect 215956 16522 215984 20431
rect 216324 16590 216352 38383
rect 216416 29481 216444 39034
rect 216494 35456 216550 35465
rect 216494 35391 216550 35400
rect 216402 29472 216458 29481
rect 216402 29407 216458 29416
rect 216312 16584 216364 16590
rect 216312 16526 216364 16532
rect 216508 16522 216536 35391
rect 216600 32473 216628 39102
rect 216586 32464 216642 32473
rect 216586 32399 216642 32408
rect 246316 23497 246344 39102
rect 246396 39092 246448 39098
rect 246396 39034 246448 39040
rect 246764 39092 246816 39098
rect 246764 39034 246816 39040
rect 246408 26489 246436 39034
rect 246670 38448 246726 38457
rect 246670 38383 246726 38392
rect 246394 26480 246450 26489
rect 246394 26415 246450 26424
rect 246302 23488 246358 23497
rect 246302 23423 246358 23432
rect 246302 20496 246358 20505
rect 246302 20431 246358 20440
rect 245658 17504 245714 17513
rect 245658 17439 245714 17448
rect 245672 16590 245700 17439
rect 245660 16584 245712 16590
rect 245660 16526 245712 16532
rect 246316 16522 246344 20431
rect 246684 16522 246712 38383
rect 246776 29481 246804 39034
rect 246854 35456 246910 35465
rect 246854 35391 246910 35400
rect 246762 29472 246818 29481
rect 246762 29407 246818 29416
rect 246868 16590 246896 35391
rect 246960 32473 246988 39102
rect 246946 32464 247002 32473
rect 246946 32399 247002 32408
rect 275296 23497 275324 39102
rect 275376 39092 275428 39098
rect 275376 39034 275428 39040
rect 275744 39092 275796 39098
rect 275744 39034 275796 39040
rect 275388 26489 275416 39034
rect 275650 38448 275706 38457
rect 275650 38383 275706 38392
rect 275374 26480 275430 26489
rect 275374 26415 275430 26424
rect 275282 23488 275338 23497
rect 275282 23423 275338 23432
rect 275282 20496 275338 20505
rect 275282 20431 275338 20440
rect 274638 17504 274694 17513
rect 274638 17439 274694 17448
rect 246856 16584 246908 16590
rect 246856 16526 246908 16532
rect 274652 16522 274680 17439
rect 275296 16590 275324 20431
rect 275284 16584 275336 16590
rect 275284 16526 275336 16532
rect 275664 16522 275692 38383
rect 275756 29481 275784 39034
rect 275834 35456 275890 35465
rect 275834 35391 275890 35400
rect 275742 29472 275798 29481
rect 275742 29407 275798 29416
rect 275848 16590 275876 35391
rect 275940 32473 275968 39102
rect 275926 32464 275982 32473
rect 275926 32399 275982 32408
rect 304276 23497 304304 39102
rect 304356 39092 304408 39098
rect 304356 39034 304408 39040
rect 304724 39092 304776 39098
rect 304724 39034 304776 39040
rect 304368 26489 304396 39034
rect 304630 38448 304686 38457
rect 304630 38383 304686 38392
rect 304354 26480 304410 26489
rect 304354 26415 304410 26424
rect 304262 23488 304318 23497
rect 304262 23423 304318 23432
rect 304262 20496 304318 20505
rect 304262 20431 304318 20440
rect 303618 17504 303674 17513
rect 303618 17439 303674 17448
rect 275836 16584 275888 16590
rect 275836 16526 275888 16532
rect 303632 16522 303660 17439
rect 304276 16590 304304 20431
rect 304644 16590 304672 38383
rect 304736 29481 304764 39034
rect 304814 35456 304870 35465
rect 304814 35391 304870 35400
rect 304722 29472 304778 29481
rect 304722 29407 304778 29416
rect 304264 16584 304316 16590
rect 304264 16526 304316 16532
rect 304632 16584 304684 16590
rect 304632 16526 304684 16532
rect 304828 16522 304856 35391
rect 304920 32473 304948 39102
rect 304906 32464 304962 32473
rect 304906 32399 304962 32408
rect 333256 23497 333284 39102
rect 333336 39092 333388 39098
rect 333336 39034 333388 39040
rect 333704 39092 333756 39098
rect 333704 39034 333756 39040
rect 333348 26489 333376 39034
rect 333610 38448 333666 38457
rect 333610 38383 333666 38392
rect 333334 26480 333390 26489
rect 333334 26415 333390 26424
rect 333242 23488 333298 23497
rect 333242 23423 333298 23432
rect 333242 20496 333298 20505
rect 333242 20431 333298 20440
rect 332598 17504 332654 17513
rect 332598 17439 332654 17448
rect 332612 16590 332640 17439
rect 332600 16584 332652 16590
rect 332600 16526 332652 16532
rect 333256 16522 333284 20431
rect 333624 16590 333652 38383
rect 333716 29481 333744 39034
rect 333794 35456 333850 35465
rect 333794 35391 333850 35400
rect 333702 29472 333758 29481
rect 333702 29407 333758 29416
rect 333612 16584 333664 16590
rect 333612 16526 333664 16532
rect 333808 16522 333836 35391
rect 333900 32473 333928 39102
rect 333886 32464 333942 32473
rect 333886 32399 333942 32408
rect 362236 23497 362264 39102
rect 362316 39092 362368 39098
rect 362316 39034 362368 39040
rect 362684 39092 362736 39098
rect 362684 39034 362736 39040
rect 362328 26489 362356 39034
rect 362590 38448 362646 38457
rect 362590 38383 362646 38392
rect 362314 26480 362370 26489
rect 362314 26415 362370 26424
rect 362222 23488 362278 23497
rect 362222 23423 362278 23432
rect 362222 20496 362278 20505
rect 362222 20431 362278 20440
rect 361578 17504 361634 17513
rect 361578 17439 361634 17448
rect 361592 16590 361620 17439
rect 361580 16584 361632 16590
rect 361580 16526 361632 16532
rect 362236 16522 362264 20431
rect 362604 16590 362632 38383
rect 362696 29481 362724 39034
rect 362774 35456 362830 35465
rect 362774 35391 362830 35400
rect 362682 29472 362738 29481
rect 362682 29407 362738 29416
rect 362592 16584 362644 16590
rect 362592 16526 362644 16532
rect 362788 16522 362816 35391
rect 362880 32473 362908 39102
rect 362866 32464 362922 32473
rect 362866 32399 362922 32408
rect 391216 23497 391244 39102
rect 391296 39092 391348 39098
rect 391296 39034 391348 39040
rect 391664 39092 391716 39098
rect 391664 39034 391716 39040
rect 391308 26489 391336 39034
rect 391570 38448 391626 38457
rect 391570 38383 391626 38392
rect 391294 26480 391350 26489
rect 391294 26415 391350 26424
rect 391202 23488 391258 23497
rect 391202 23423 391258 23432
rect 391202 20496 391258 20505
rect 391202 20431 391258 20440
rect 390558 17504 390614 17513
rect 390558 17439 390614 17448
rect 390572 16590 390600 17439
rect 390560 16584 390612 16590
rect 390560 16526 390612 16532
rect 391216 16522 391244 20431
rect 391584 16522 391612 38383
rect 391676 29481 391704 39034
rect 391754 35456 391810 35465
rect 391754 35391 391810 35400
rect 391662 29472 391718 29481
rect 391662 29407 391718 29416
rect 391768 16590 391796 35391
rect 391860 32473 391888 39102
rect 391846 32464 391902 32473
rect 391846 32399 391902 32408
rect 420196 23497 420224 39102
rect 420276 39092 420328 39098
rect 420276 39034 420328 39040
rect 420644 39092 420696 39098
rect 420644 39034 420696 39040
rect 420288 26489 420316 39034
rect 420550 38448 420606 38457
rect 420550 38383 420606 38392
rect 420274 26480 420330 26489
rect 420274 26415 420330 26424
rect 420182 23488 420238 23497
rect 420182 23423 420238 23432
rect 420182 20496 420238 20505
rect 420182 20431 420238 20440
rect 419538 17504 419594 17513
rect 419538 17439 419594 17448
rect 391756 16584 391808 16590
rect 391756 16526 391808 16532
rect 419552 16522 419580 17439
rect 420196 16590 420224 20431
rect 420184 16584 420236 16590
rect 420184 16526 420236 16532
rect 420564 16522 420592 38383
rect 420656 29481 420684 39034
rect 420734 35456 420790 35465
rect 420734 35391 420790 35400
rect 420642 29472 420698 29481
rect 420642 29407 420698 29416
rect 420748 16590 420776 35391
rect 420840 32473 420868 39102
rect 420826 32464 420882 32473
rect 420826 32399 420882 32408
rect 449176 23497 449204 39102
rect 449256 39092 449308 39098
rect 449256 39034 449308 39040
rect 449624 39092 449676 39098
rect 449624 39034 449676 39040
rect 449268 26489 449296 39034
rect 449530 38448 449586 38457
rect 449530 38383 449586 38392
rect 449254 26480 449310 26489
rect 449254 26415 449310 26424
rect 449162 23488 449218 23497
rect 449162 23423 449218 23432
rect 449162 20496 449218 20505
rect 449162 20431 449218 20440
rect 448518 17504 448574 17513
rect 448518 17439 448574 17448
rect 420736 16584 420788 16590
rect 420736 16526 420788 16532
rect 448532 16522 448560 17439
rect 449176 16590 449204 20431
rect 449164 16584 449216 16590
rect 449164 16526 449216 16532
rect 449544 16522 449572 38383
rect 449636 29481 449664 39034
rect 449714 35456 449770 35465
rect 449714 35391 449770 35400
rect 449622 29472 449678 29481
rect 449622 29407 449678 29416
rect 449728 16590 449756 35391
rect 449820 32473 449848 39102
rect 449806 32464 449862 32473
rect 449806 32399 449862 32408
rect 478156 23497 478184 39102
rect 478236 39092 478288 39098
rect 478236 39034 478288 39040
rect 478604 39092 478656 39098
rect 478604 39034 478656 39040
rect 478248 26489 478276 39034
rect 478510 38448 478566 38457
rect 478510 38383 478566 38392
rect 478234 26480 478290 26489
rect 478234 26415 478290 26424
rect 478142 23488 478198 23497
rect 478142 23423 478198 23432
rect 478142 20496 478198 20505
rect 478142 20431 478198 20440
rect 477498 17504 477554 17513
rect 477498 17439 477554 17448
rect 449716 16584 449768 16590
rect 449716 16526 449768 16532
rect 477512 16522 477540 17439
rect 478156 16590 478184 20431
rect 478524 16590 478552 38383
rect 478616 29481 478644 39034
rect 478694 35456 478750 35465
rect 478694 35391 478750 35400
rect 478602 29472 478658 29481
rect 478602 29407 478658 29416
rect 478144 16584 478196 16590
rect 478144 16526 478196 16532
rect 478512 16584 478564 16590
rect 478512 16526 478564 16532
rect 478708 16522 478736 35391
rect 478800 32473 478828 39102
rect 478786 32464 478842 32473
rect 478786 32399 478842 32408
rect 507136 24041 507164 39102
rect 507216 39092 507268 39098
rect 507216 39034 507268 39040
rect 507584 39092 507636 39098
rect 507584 39034 507636 39040
rect 507228 27033 507256 39034
rect 507490 37904 507546 37913
rect 507490 37839 507546 37848
rect 507214 27024 507270 27033
rect 507214 26959 507270 26968
rect 507122 24032 507178 24041
rect 507122 23967 507178 23976
rect 507122 19952 507178 19961
rect 507122 19887 507178 19896
rect 506478 17096 506534 17105
rect 506478 17031 506534 17040
rect 506492 16590 506520 17031
rect 506480 16584 506532 16590
rect 506480 16526 506532 16532
rect 507136 16522 507164 19887
rect 507504 16522 507532 37839
rect 507596 30025 507624 39034
rect 507674 34912 507730 34921
rect 507674 34847 507730 34856
rect 507582 30016 507638 30025
rect 507582 29951 507638 29960
rect 507688 16590 507716 34847
rect 507780 33017 507808 39102
rect 507766 33008 507822 33017
rect 507766 32943 507822 32952
rect 536116 23497 536144 39102
rect 536196 39092 536248 39098
rect 536196 39034 536248 39040
rect 536208 26489 536236 39034
rect 536576 35465 536604 39510
rect 536748 39432 536800 39438
rect 536748 39374 536800 39380
rect 536656 39364 536708 39370
rect 536656 39306 536708 39312
rect 536562 35456 536618 35465
rect 536562 35391 536618 35400
rect 536668 32473 536696 39306
rect 536654 32464 536710 32473
rect 536654 32399 536710 32408
rect 536760 29481 536788 39374
rect 538140 38593 538168 40666
rect 567396 39574 567424 50918
rect 567384 39568 567436 39574
rect 567384 39510 567436 39516
rect 567488 39370 567516 51054
rect 567580 43858 567608 53615
rect 567658 50688 567714 50697
rect 567658 50623 567714 50632
rect 567672 43926 567700 50623
rect 567660 43920 567712 43926
rect 567660 43862 567712 43868
rect 567568 43852 567620 43858
rect 567568 43794 567620 43800
rect 567764 39438 567792 55186
rect 567752 39432 567804 39438
rect 567752 39374 567804 39380
rect 567476 39364 567528 39370
rect 567476 39306 567528 39312
rect 580172 39024 580224 39030
rect 580172 38966 580224 38972
rect 538126 38584 538182 38593
rect 538126 38519 538182 38528
rect 580184 33153 580212 38966
rect 580170 33144 580226 33153
rect 580170 33079 580226 33088
rect 536746 29472 536802 29481
rect 536746 29407 536802 29416
rect 536194 26480 536250 26489
rect 536194 26415 536250 26424
rect 536102 23488 536158 23497
rect 536102 23423 536158 23432
rect 536102 20496 536158 20505
rect 536102 20431 536158 20440
rect 535458 17504 535514 17513
rect 535458 17439 535514 17448
rect 507676 16584 507728 16590
rect 507676 16526 507728 16532
rect 535472 16522 535500 17439
rect 536116 16590 536144 20431
rect 536104 16584 536156 16590
rect 536104 16526 536156 16532
rect 157524 16516 157576 16522
rect 157524 16458 157576 16464
rect 158352 16516 158404 16522
rect 158352 16458 158404 16464
rect 186780 16516 186832 16522
rect 186780 16458 186832 16464
rect 187516 16516 187568 16522
rect 187516 16458 187568 16464
rect 215944 16516 215996 16522
rect 215944 16458 215996 16464
rect 216496 16516 216548 16522
rect 216496 16458 216548 16464
rect 246304 16516 246356 16522
rect 246304 16458 246356 16464
rect 246672 16516 246724 16522
rect 246672 16458 246724 16464
rect 274640 16516 274692 16522
rect 274640 16458 274692 16464
rect 275652 16516 275704 16522
rect 275652 16458 275704 16464
rect 303620 16516 303672 16522
rect 303620 16458 303672 16464
rect 304816 16516 304868 16522
rect 304816 16458 304868 16464
rect 333244 16516 333296 16522
rect 333244 16458 333296 16464
rect 333796 16516 333848 16522
rect 333796 16458 333848 16464
rect 362224 16516 362276 16522
rect 362224 16458 362276 16464
rect 362776 16516 362828 16522
rect 362776 16458 362828 16464
rect 391204 16516 391256 16522
rect 391204 16458 391256 16464
rect 391572 16516 391624 16522
rect 391572 16458 391624 16464
rect 419540 16516 419592 16522
rect 419540 16458 419592 16464
rect 420552 16516 420604 16522
rect 420552 16458 420604 16464
rect 448520 16516 448572 16522
rect 448520 16458 448572 16464
rect 449532 16516 449584 16522
rect 449532 16458 449584 16464
rect 477500 16516 477552 16522
rect 477500 16458 477552 16464
rect 478696 16516 478748 16522
rect 478696 16458 478748 16464
rect 507124 16516 507176 16522
rect 507124 16458 507176 16464
rect 507492 16516 507544 16522
rect 507492 16458 507544 16464
rect 535460 16516 535512 16522
rect 535460 16458 535512 16464
rect 580276 13326 580304 670647
rect 580354 644056 580410 644065
rect 580354 643991 580410 644000
rect 580368 13462 580396 643991
rect 580446 617536 580502 617545
rect 580446 617471 580502 617480
rect 580356 13456 580408 13462
rect 580356 13398 580408 13404
rect 580460 13394 580488 617471
rect 580538 484664 580594 484673
rect 580538 484599 580594 484608
rect 580552 13598 580580 484599
rect 580630 351928 580686 351937
rect 580630 351863 580686 351872
rect 580540 13592 580592 13598
rect 580540 13534 580592 13540
rect 580644 13530 580672 351863
rect 580722 325272 580778 325281
rect 580722 325207 580778 325216
rect 580736 13802 580764 325207
rect 580814 272232 580870 272241
rect 580814 272167 580870 272176
rect 580724 13796 580776 13802
rect 580724 13738 580776 13744
rect 580828 13734 580856 272167
rect 580906 72992 580962 73001
rect 580906 72927 580962 72936
rect 580816 13728 580868 13734
rect 580816 13670 580868 13676
rect 580920 13666 580948 72927
rect 580908 13660 580960 13666
rect 580908 13602 580960 13608
rect 580632 13524 580684 13530
rect 580632 13466 580684 13472
rect 580448 13388 580500 13394
rect 580448 13330 580500 13336
rect 580264 13320 580316 13326
rect 580264 13262 580316 13268
rect 137008 13252 137060 13258
rect 137008 13194 137060 13200
rect 71780 13184 71832 13190
rect 71780 13126 71832 13132
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 33140 3528 33192 3534
rect 33140 3470 33192 3476
rect 64236 3528 64288 3534
rect 64236 3470 64288 3476
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 125888 480 125916 3538
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 132958 3496 133014 3505
rect 126992 480 127020 3470
rect 129372 3460 129424 3466
rect 132958 3431 133014 3440
rect 129372 3402 129424 3408
rect 129384 480 129412 3402
rect 132972 480 133000 3431
rect 136454 3360 136510 3369
rect 136454 3295 136510 3304
rect 136468 480 136496 3295
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 658144 3478 658200
rect 2778 632068 2780 632088
rect 2780 632068 2832 632088
rect 2832 632068 2834 632088
rect 2778 632032 2834 632068
rect 2962 579944 3018 580000
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3146 449520 3202 449576
rect 3422 410488 3478 410544
rect 3330 358400 3386 358456
rect 2778 345344 2834 345400
rect 3330 293120 3386 293176
rect 3146 254088 3202 254144
rect 3330 201864 3386 201920
rect 3330 136720 3386 136776
rect 3330 58520 3386 58576
rect 3238 45464 3294 45520
rect 3514 397432 3570 397488
rect 3606 306176 3662 306232
rect 3698 241032 3754 241088
rect 3790 188808 3846 188864
rect 3882 149776 3938 149832
rect 3698 19352 3754 19408
rect 3974 97552 4030 97608
rect 4066 84632 4122 84688
rect 13542 39344 13598 39400
rect 12438 34468 12494 34504
rect 12438 34448 12440 34468
rect 12440 34448 12492 34468
rect 12492 34448 12494 34468
rect 12438 31048 12494 31104
rect 54666 37848 54722 37904
rect 39670 35264 39726 35320
rect 43442 35264 43498 35320
rect 50526 35264 50582 35320
rect 13726 33088 13782 33144
rect 13634 29688 13690 29744
rect 13542 27648 13598 27704
rect 13634 26288 13690 26344
rect 12438 22888 12494 22944
rect 12438 20848 12494 20904
rect 11794 19488 11850 19544
rect 12438 17448 12494 17504
rect 61290 34312 61346 34368
rect 13726 24112 13782 24168
rect 61290 20576 61346 20632
rect 63498 26968 63554 27024
rect 64234 31592 64290 31648
rect 64234 30232 64290 30288
rect 64142 23568 64198 23624
rect 63498 21392 63554 21448
rect 46018 16496 46074 16552
rect 57610 16496 57666 16552
rect 26974 13232 27030 13288
rect 19246 12960 19302 13016
rect 35346 13504 35402 13560
rect 41786 13368 41842 13424
rect 48226 13096 48282 13152
rect 52734 13504 52790 13560
rect 64326 28328 64382 28384
rect 64326 24928 64382 24984
rect 64510 35128 64566 35184
rect 64418 18128 64474 18184
rect 71410 32408 71466 32464
rect 71686 38392 71742 38448
rect 71594 35400 71650 35456
rect 71502 29416 71558 29472
rect 71042 26424 71098 26480
rect 70398 20440 70454 20496
rect 70398 17448 70454 17504
rect 64602 16768 64658 16824
rect 71134 23432 71190 23488
rect 100390 32408 100446 32464
rect 100666 38392 100722 38448
rect 100574 35400 100630 35456
rect 100482 29416 100538 29472
rect 100114 26424 100170 26480
rect 100022 23432 100078 23488
rect 100022 20440 100078 20496
rect 99838 17448 99894 17504
rect 129370 38392 129426 38448
rect 129094 26424 129150 26480
rect 129002 23432 129058 23488
rect 129002 20440 129058 20496
rect 128818 17448 128874 17504
rect 129554 35400 129610 35456
rect 129462 29416 129518 29472
rect 129646 32408 129702 32464
rect 170310 699760 170366 699816
rect 397458 699760 397514 699816
rect 429842 699760 429898 699816
rect 527178 699760 527234 699816
rect 559654 699760 559710 699816
rect 580170 697176 580226 697232
rect 580262 670656 580318 670712
rect 580170 590960 580226 591016
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 580170 511264 580226 511320
rect 579986 471416 580042 471472
rect 579618 431568 579674 431624
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579802 232328 579858 232384
rect 580170 192480 580226 192536
rect 579986 152632 580042 152688
rect 579986 112784 580042 112840
rect 451922 65592 451978 65648
rect 480902 65592 480958 65648
rect 509882 65592 509938 65648
rect 538862 65592 538918 65648
rect 567198 65592 567254 65648
rect 220082 65048 220138 65104
rect 219438 47096 219494 47152
rect 217138 44104 217194 44160
rect 249154 62600 249210 62656
rect 278042 62600 278098 62656
rect 307022 62600 307078 62656
rect 336002 62600 336058 62656
rect 364982 62600 365038 62656
rect 393962 62600 394018 62656
rect 422942 62600 422998 62656
rect 220266 62192 220322 62248
rect 220174 59336 220230 59392
rect 249062 59608 249118 59664
rect 220358 56752 220414 56808
rect 248418 53624 248474 53680
rect 246118 47096 246174 47152
rect 248510 50632 248566 50688
rect 249246 56616 249302 56672
rect 277398 53624 277454 53680
rect 275098 47096 275154 47152
rect 220266 43560 220322 43616
rect 245934 43560 245990 43616
rect 249154 43560 249210 43616
rect 275006 43560 275062 43616
rect 277490 50632 277546 50688
rect 278134 59608 278190 59664
rect 278226 56616 278282 56672
rect 306562 53624 306618 53680
rect 306470 50632 306526 50688
rect 304078 47096 304134 47152
rect 307114 59608 307170 59664
rect 307206 56616 307262 56672
rect 335358 53624 335414 53680
rect 333150 47096 333206 47152
rect 335450 50632 335506 50688
rect 336094 59608 336150 59664
rect 336186 56616 336242 56672
rect 364338 53624 364394 53680
rect 362130 47096 362186 47152
rect 364430 50632 364486 50688
rect 365074 59608 365130 59664
rect 365166 56616 365222 56672
rect 393318 53624 393374 53680
rect 391110 47096 391166 47152
rect 393410 50632 393466 50688
rect 394054 59608 394110 59664
rect 394146 56616 394202 56672
rect 422298 53624 422354 53680
rect 420090 47096 420146 47152
rect 422390 50632 422446 50688
rect 423034 59608 423090 59664
rect 423126 56616 423182 56672
rect 451462 53624 451518 53680
rect 451370 50632 451426 50688
rect 449070 47096 449126 47152
rect 452014 62600 452070 62656
rect 452106 59608 452162 59664
rect 452198 56616 452254 56672
rect 480442 53624 480498 53680
rect 480350 50632 480406 50688
rect 480258 47640 480314 47696
rect 480994 62600 481050 62656
rect 481086 59608 481142 59664
rect 481178 56616 481234 56672
rect 509422 53624 509478 53680
rect 509330 50632 509386 50688
rect 509238 47640 509294 47696
rect 509974 62600 510030 62656
rect 510066 59608 510122 59664
rect 510158 56616 510214 56672
rect 538402 53624 538458 53680
rect 538310 50632 538366 50688
rect 538218 47640 538274 47696
rect 538954 62600 539010 62656
rect 539046 59608 539102 59664
rect 539138 56616 539194 56672
rect 567290 62600 567346 62656
rect 567382 59608 567438 59664
rect 567474 56616 567530 56672
rect 567566 53624 567622 53680
rect 567198 47640 567254 47696
rect 565082 44104 565138 44160
rect 451922 43560 451978 43616
rect 480902 43560 480958 43616
rect 509882 43560 509938 43616
rect 220082 43288 220138 43344
rect 217138 39344 217194 39400
rect 158350 38392 158406 38448
rect 158074 26424 158130 26480
rect 157982 23432 158038 23488
rect 157982 20440 158038 20496
rect 157522 17448 157578 17504
rect 158534 35400 158590 35456
rect 158442 29416 158498 29472
rect 158626 32408 158682 32464
rect 187330 38392 187386 38448
rect 187054 26424 187110 26480
rect 186962 23432 187018 23488
rect 186962 20440 187018 20496
rect 186778 17448 186834 17504
rect 187514 35400 187570 35456
rect 187422 29416 187478 29472
rect 187606 32408 187662 32464
rect 216310 38392 216366 38448
rect 216034 26424 216090 26480
rect 215942 23432 215998 23488
rect 215942 20440 215998 20496
rect 215758 17448 215814 17504
rect 216494 35400 216550 35456
rect 216402 29416 216458 29472
rect 216586 32408 216642 32464
rect 246670 38392 246726 38448
rect 246394 26424 246450 26480
rect 246302 23432 246358 23488
rect 246302 20440 246358 20496
rect 245658 17448 245714 17504
rect 246854 35400 246910 35456
rect 246762 29416 246818 29472
rect 246946 32408 247002 32464
rect 275650 38392 275706 38448
rect 275374 26424 275430 26480
rect 275282 23432 275338 23488
rect 275282 20440 275338 20496
rect 274638 17448 274694 17504
rect 275834 35400 275890 35456
rect 275742 29416 275798 29472
rect 275926 32408 275982 32464
rect 304630 38392 304686 38448
rect 304354 26424 304410 26480
rect 304262 23432 304318 23488
rect 304262 20440 304318 20496
rect 303618 17448 303674 17504
rect 304814 35400 304870 35456
rect 304722 29416 304778 29472
rect 304906 32408 304962 32464
rect 333610 38392 333666 38448
rect 333334 26424 333390 26480
rect 333242 23432 333298 23488
rect 333242 20440 333298 20496
rect 332598 17448 332654 17504
rect 333794 35400 333850 35456
rect 333702 29416 333758 29472
rect 333886 32408 333942 32464
rect 362590 38392 362646 38448
rect 362314 26424 362370 26480
rect 362222 23432 362278 23488
rect 362222 20440 362278 20496
rect 361578 17448 361634 17504
rect 362774 35400 362830 35456
rect 362682 29416 362738 29472
rect 362866 32408 362922 32464
rect 391570 38392 391626 38448
rect 391294 26424 391350 26480
rect 391202 23432 391258 23488
rect 391202 20440 391258 20496
rect 390558 17448 390614 17504
rect 391754 35400 391810 35456
rect 391662 29416 391718 29472
rect 391846 32408 391902 32464
rect 420550 38392 420606 38448
rect 420274 26424 420330 26480
rect 420182 23432 420238 23488
rect 420182 20440 420238 20496
rect 419538 17448 419594 17504
rect 420734 35400 420790 35456
rect 420642 29416 420698 29472
rect 420826 32408 420882 32464
rect 449530 38392 449586 38448
rect 449254 26424 449310 26480
rect 449162 23432 449218 23488
rect 449162 20440 449218 20496
rect 448518 17448 448574 17504
rect 449714 35400 449770 35456
rect 449622 29416 449678 29472
rect 449806 32408 449862 32464
rect 478510 38392 478566 38448
rect 478234 26424 478290 26480
rect 478142 23432 478198 23488
rect 478142 20440 478198 20496
rect 477498 17448 477554 17504
rect 478694 35400 478750 35456
rect 478602 29416 478658 29472
rect 478786 32408 478842 32464
rect 507490 37848 507546 37904
rect 507214 26968 507270 27024
rect 507122 23976 507178 24032
rect 507122 19896 507178 19952
rect 506478 17040 506534 17096
rect 507674 34856 507730 34912
rect 507582 29960 507638 30016
rect 507766 32952 507822 33008
rect 536562 35400 536618 35456
rect 536654 32408 536710 32464
rect 567658 50632 567714 50688
rect 538126 38528 538182 38584
rect 580170 33088 580226 33144
rect 536746 29416 536802 29472
rect 536194 26424 536250 26480
rect 536102 23432 536158 23488
rect 536102 20440 536158 20496
rect 535458 17448 535514 17504
rect 580354 644000 580410 644056
rect 580446 617480 580502 617536
rect 580538 484608 580594 484664
rect 580630 351872 580686 351928
rect 580722 325216 580778 325272
rect 580814 272176 580870 272232
rect 580906 72936 580962 72992
rect 132958 3440 133014 3496
rect 136454 3304 136510 3360
<< metal3 >>
rect 169702 699756 169708 699820
rect 169772 699818 169778 699820
rect 170305 699818 170371 699821
rect 169772 699816 170371 699818
rect 169772 699760 170310 699816
rect 170366 699760 170371 699816
rect 169772 699758 170371 699760
rect 169772 699756 169778 699758
rect 170305 699755 170371 699758
rect 397453 699818 397519 699821
rect 397678 699818 397684 699820
rect 397453 699816 397684 699818
rect 397453 699760 397458 699816
rect 397514 699760 397684 699816
rect 397453 699758 397684 699760
rect 397453 699755 397519 699758
rect 397678 699756 397684 699758
rect 397748 699756 397754 699820
rect 429326 699756 429332 699820
rect 429396 699818 429402 699820
rect 429837 699818 429903 699821
rect 429396 699816 429903 699818
rect 429396 699760 429842 699816
rect 429898 699760 429903 699816
rect 429396 699758 429903 699760
rect 429396 699756 429402 699758
rect 429837 699755 429903 699758
rect 527173 699818 527239 699821
rect 527398 699818 527404 699820
rect 527173 699816 527404 699818
rect 527173 699760 527178 699816
rect 527234 699760 527404 699816
rect 527173 699758 527404 699760
rect 527173 699755 527239 699758
rect 527398 699756 527404 699758
rect 527468 699756 527474 699820
rect 558862 699756 558868 699820
rect 558932 699818 558938 699820
rect 559649 699818 559715 699821
rect 558932 699816 559715 699818
rect 558932 699760 559654 699816
rect 559710 699760 559715 699816
rect 558932 699758 559715 699760
rect 558932 699756 558938 699758
rect 559649 699755 559715 699758
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3366 684314 3372 684316
rect -960 684254 3372 684314
rect -960 684164 480 684254
rect 3366 684252 3372 684254
rect 3436 684252 3442 684316
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580349 644058 580415 644061
rect 583520 644058 584960 644148
rect 580349 644056 584960 644058
rect 580349 644000 580354 644056
rect 580410 644000 584960 644056
rect 580349 643998 584960 644000
rect 580349 643995 580415 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 580441 617538 580507 617541
rect 583520 617538 584960 617628
rect 580441 617536 584960 617538
rect 580441 617480 580446 617536
rect 580502 617480 584960 617536
rect 580441 617478 584960 617480
rect 580441 617475 580507 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3550 606114 3556 606116
rect -960 606054 3556 606114
rect -960 605964 480 606054
rect 3550 606052 3556 606054
rect 3620 606052 3626 606116
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 2957 580002 3023 580005
rect -960 580000 3023 580002
rect -960 579944 2962 580000
rect 3018 579944 3023 580000
rect -960 579942 3023 579944
rect -960 579852 480 579942
rect 2957 579939 3023 579942
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect -960 501742 674 501802
rect -960 501666 480 501742
rect 614 501666 674 501742
rect -960 501652 674 501666
rect 246 501606 674 501652
rect 246 501122 306 501606
rect 246 501062 6930 501122
rect 6870 500986 6930 501062
rect 45318 500986 45324 500988
rect 6870 500926 45324 500986
rect 45318 500924 45324 500926
rect 45388 500924 45394 500988
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580533 484666 580599 484669
rect 583520 484666 584960 484756
rect 580533 484664 584960 484666
rect 580533 484608 580538 484664
rect 580594 484608 584960 484664
rect 580533 484606 584960 484608
rect 580533 484603 580599 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect -960 475630 674 475690
rect -960 475554 480 475630
rect 614 475554 674 475630
rect -960 475540 674 475554
rect 246 475494 674 475540
rect 246 475010 306 475494
rect 246 474950 6930 475010
rect 6870 474874 6930 474950
rect 54334 474874 54340 474876
rect 6870 474814 54340 474874
rect 54334 474812 54340 474814
rect 54404 474812 54410 474876
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579613 431626 579679 431629
rect 583520 431626 584960 431716
rect 579613 431624 584960 431626
rect 579613 431568 579618 431624
rect 579674 431568 584960 431624
rect 579613 431566 584960 431568
rect 579613 431563 579679 431566
rect 583520 431476 584960 431566
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 580625 351930 580691 351933
rect 583520 351930 584960 352020
rect 580625 351928 584960 351930
rect 580625 351872 580630 351928
rect 580686 351872 584960 351928
rect 580625 351870 584960 351872
rect 580625 351867 580691 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580717 325274 580783 325277
rect 583520 325274 584960 325364
rect 580717 325272 584960 325274
rect 580717 325216 580722 325272
rect 580778 325216 584960 325272
rect 580717 325214 584960 325216
rect 580717 325211 580783 325214
rect 583520 325124 584960 325214
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306234 480 306324
rect 3601 306234 3667 306237
rect -960 306232 3667 306234
rect -960 306176 3606 306232
rect 3662 306176 3667 306232
rect -960 306174 3667 306176
rect -960 306084 480 306174
rect 3601 306171 3667 306174
rect 583520 298604 584960 298844
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580809 272234 580875 272237
rect 583520 272234 584960 272324
rect 580809 272232 584960 272234
rect 580809 272176 580814 272232
rect 580870 272176 584960 272232
rect 580809 272174 584960 272176
rect 580809 272171 580875 272174
rect 583520 272084 584960 272174
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 583520 245428 584960 245668
rect -960 241090 480 241180
rect 3693 241090 3759 241093
rect -960 241088 3759 241090
rect -960 241032 3698 241088
rect 3754 241032 3759 241088
rect -960 241030 3759 241032
rect -960 240940 480 241030
rect 3693 241027 3759 241030
rect 579797 232386 579863 232389
rect 583520 232386 584960 232476
rect 579797 232384 584960 232386
rect 579797 232328 579802 232384
rect 579858 232328 584960 232384
rect 579797 232326 584960 232328
rect 579797 232323 579863 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201922 480 202012
rect 3325 201922 3391 201925
rect -960 201920 3391 201922
rect -960 201864 3330 201920
rect 3386 201864 3391 201920
rect -960 201862 3391 201864
rect -960 201772 480 201862
rect 3325 201859 3391 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3785 188866 3851 188869
rect -960 188864 3851 188866
rect -960 188808 3790 188864
rect 3846 188808 3851 188864
rect -960 188806 3851 188808
rect -960 188716 480 188806
rect 3785 188803 3851 188806
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3877 149834 3943 149837
rect -960 149832 3943 149834
rect -960 149776 3882 149832
rect 3938 149776 3943 149832
rect -960 149774 3943 149776
rect -960 149684 480 149774
rect 3877 149771 3943 149774
rect 583520 139212 584960 139452
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 579981 112842 580047 112845
rect 583520 112842 584960 112932
rect 579981 112840 584960 112842
rect 579981 112784 579986 112840
rect 580042 112784 584960 112840
rect 579981 112782 584960 112784
rect 579981 112779 580047 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 3969 97610 4035 97613
rect -960 97608 4035 97610
rect -960 97552 3974 97608
rect 4030 97552 4035 97608
rect -960 97550 4035 97552
rect -960 97460 480 97550
rect 3969 97547 4035 97550
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 4061 84690 4127 84693
rect -960 84688 4127 84690
rect -960 84632 4066 84688
rect 4122 84632 4127 84688
rect -960 84630 4127 84632
rect -960 84540 480 84630
rect 4061 84627 4127 84630
rect 580901 72994 580967 72997
rect 583520 72994 584960 73084
rect 580901 72992 584960 72994
rect 580901 72936 580906 72992
rect 580962 72936 584960 72992
rect 580901 72934 584960 72936
rect 580901 72931 580967 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 265758 66406 269866 66466
rect 207828 66270 211876 66330
rect 236900 66270 240948 66330
rect 265758 66300 265818 66406
rect 269806 66300 269866 66406
rect 410934 66406 415042 66466
rect 294860 66270 298908 66330
rect 323932 66270 327980 66330
rect 352820 66270 356868 66330
rect 381892 66270 385940 66330
rect 410934 66300 410994 66406
rect 414982 66300 415042 66406
rect 439852 66270 443900 66330
rect 468924 66270 472972 66330
rect 497812 66270 501860 66330
rect 526884 66270 530932 66330
rect 555956 66270 560004 66330
rect 249006 65650 249012 65652
rect 217734 65106 217794 65620
rect 246652 65590 249012 65650
rect 249006 65588 249012 65590
rect 249076 65588 249082 65652
rect 277894 65650 277900 65652
rect 275724 65590 277900 65650
rect 277894 65588 277900 65590
rect 277964 65588 277970 65652
rect 306966 65650 306972 65652
rect 304612 65590 306972 65650
rect 306966 65588 306972 65590
rect 307036 65588 307042 65652
rect 335854 65650 335860 65652
rect 333684 65590 335860 65650
rect 335854 65588 335860 65590
rect 335924 65588 335930 65652
rect 364926 65650 364932 65652
rect 362756 65590 364932 65650
rect 364926 65588 364932 65590
rect 364996 65588 365002 65652
rect 393814 65650 393820 65652
rect 391644 65590 393820 65650
rect 393814 65588 393820 65590
rect 393884 65588 393890 65652
rect 422886 65650 422892 65652
rect 420716 65590 422892 65650
rect 422886 65588 422892 65590
rect 422956 65588 422962 65652
rect 451917 65650 451983 65653
rect 480897 65650 480963 65653
rect 509877 65650 509943 65653
rect 538857 65650 538923 65653
rect 567193 65650 567259 65653
rect 449604 65648 451983 65650
rect 449604 65592 451922 65648
rect 451978 65592 451983 65648
rect 449604 65590 451983 65592
rect 478676 65648 480963 65650
rect 478676 65592 480902 65648
rect 480958 65592 480963 65648
rect 478676 65590 480963 65592
rect 507748 65648 509943 65650
rect 507748 65592 509882 65648
rect 509938 65592 509943 65648
rect 507748 65590 509943 65592
rect 536636 65648 538923 65650
rect 536636 65592 538862 65648
rect 538918 65592 538923 65648
rect 536636 65590 538923 65592
rect 565708 65648 567259 65650
rect 565708 65592 567198 65648
rect 567254 65592 567259 65648
rect 565708 65590 567259 65592
rect 451917 65587 451983 65590
rect 480897 65587 480963 65590
rect 509877 65587 509943 65590
rect 538857 65587 538923 65590
rect 567193 65587 567259 65590
rect 220077 65106 220143 65109
rect 217734 65104 220143 65106
rect 217734 65048 220082 65104
rect 220138 65048 220143 65104
rect 217734 65046 220143 65048
rect 220077 65043 220143 65046
rect 207828 64774 211876 64834
rect 236900 64774 240948 64834
rect 265758 64698 265818 64804
rect 269806 64698 269866 64804
rect 294860 64774 298908 64834
rect 323932 64774 327980 64834
rect 352820 64774 356868 64834
rect 381892 64774 385940 64834
rect 265758 64638 269866 64698
rect 410934 64698 410994 64804
rect 414982 64698 415042 64804
rect 439852 64774 443900 64834
rect 468924 64774 472972 64834
rect 497812 64774 501860 64834
rect 526884 64774 530932 64834
rect 555956 64774 560004 64834
rect 410934 64638 415042 64698
rect 265758 63414 269866 63474
rect 207828 63278 211876 63338
rect 236900 63278 240948 63338
rect 265758 63308 265818 63414
rect 269806 63308 269866 63414
rect 410934 63414 415042 63474
rect 294860 63278 298908 63338
rect 323932 63278 327980 63338
rect 352820 63278 356868 63338
rect 381892 63278 385940 63338
rect 410934 63308 410994 63414
rect 414982 63308 415042 63414
rect 439852 63278 443900 63338
rect 468924 63278 472972 63338
rect 497812 63278 501860 63338
rect 526884 63278 530932 63338
rect 555956 63278 560004 63338
rect 249149 62658 249215 62661
rect 278037 62658 278103 62661
rect 307017 62658 307083 62661
rect 335997 62658 336063 62661
rect 364977 62658 365043 62661
rect 393957 62658 394023 62661
rect 422937 62658 423003 62661
rect 452009 62658 452075 62661
rect 480989 62658 481055 62661
rect 509969 62658 510035 62661
rect 538949 62658 539015 62661
rect 567285 62658 567351 62661
rect 246652 62656 249215 62658
rect 217734 62250 217794 62628
rect 246652 62600 249154 62656
rect 249210 62600 249215 62656
rect 246652 62598 249215 62600
rect 275724 62656 278103 62658
rect 275724 62600 278042 62656
rect 278098 62600 278103 62656
rect 275724 62598 278103 62600
rect 304612 62656 307083 62658
rect 304612 62600 307022 62656
rect 307078 62600 307083 62656
rect 304612 62598 307083 62600
rect 333684 62656 336063 62658
rect 333684 62600 336002 62656
rect 336058 62600 336063 62656
rect 333684 62598 336063 62600
rect 362756 62656 365043 62658
rect 362756 62600 364982 62656
rect 365038 62600 365043 62656
rect 362756 62598 365043 62600
rect 391644 62656 394023 62658
rect 391644 62600 393962 62656
rect 394018 62600 394023 62656
rect 391644 62598 394023 62600
rect 420716 62656 423003 62658
rect 420716 62600 422942 62656
rect 422998 62600 423003 62656
rect 420716 62598 423003 62600
rect 449604 62656 452075 62658
rect 449604 62600 452014 62656
rect 452070 62600 452075 62656
rect 449604 62598 452075 62600
rect 478676 62656 481055 62658
rect 478676 62600 480994 62656
rect 481050 62600 481055 62656
rect 478676 62598 481055 62600
rect 507748 62656 510035 62658
rect 507748 62600 509974 62656
rect 510030 62600 510035 62656
rect 507748 62598 510035 62600
rect 536636 62656 539015 62658
rect 536636 62600 538954 62656
rect 539010 62600 539015 62656
rect 536636 62598 539015 62600
rect 565708 62656 567351 62658
rect 565708 62600 567290 62656
rect 567346 62600 567351 62656
rect 565708 62598 567351 62600
rect 249149 62595 249215 62598
rect 278037 62595 278103 62598
rect 307017 62595 307083 62598
rect 335997 62595 336063 62598
rect 364977 62595 365043 62598
rect 393957 62595 394023 62598
rect 422937 62595 423003 62598
rect 452009 62595 452075 62598
rect 480989 62595 481055 62598
rect 509969 62595 510035 62598
rect 538949 62595 539015 62598
rect 567285 62595 567351 62598
rect 220261 62250 220327 62253
rect 217734 62248 220327 62250
rect 217734 62192 220266 62248
rect 220322 62192 220327 62248
rect 217734 62190 220327 62192
rect 220261 62187 220327 62190
rect 265758 61918 269866 61978
rect 207828 61782 211876 61842
rect 236900 61782 240948 61842
rect 265758 61812 265818 61918
rect 269806 61812 269866 61918
rect 410934 61918 415042 61978
rect 294860 61782 298908 61842
rect 323932 61782 327980 61842
rect 352820 61782 356868 61842
rect 381892 61782 385940 61842
rect 410934 61812 410994 61918
rect 414982 61812 415042 61918
rect 439852 61782 443900 61842
rect 468924 61782 472972 61842
rect 497812 61782 501860 61842
rect 526884 61782 530932 61842
rect 555956 61782 560004 61842
rect 265758 60422 269866 60482
rect 207828 60286 211876 60346
rect 236900 60286 240948 60346
rect 265758 60316 265818 60422
rect 269806 60316 269866 60422
rect 410934 60422 415042 60482
rect 294860 60286 298908 60346
rect 323932 60286 327980 60346
rect 352820 60286 356868 60346
rect 381892 60286 385940 60346
rect 410934 60316 410994 60422
rect 414982 60316 415042 60422
rect 439852 60286 443900 60346
rect 468924 60286 472972 60346
rect 497812 60286 501860 60346
rect 526884 60286 530932 60346
rect 555956 60286 560004 60346
rect 249057 59666 249123 59669
rect 278129 59666 278195 59669
rect 307109 59666 307175 59669
rect 336089 59666 336155 59669
rect 365069 59666 365135 59669
rect 394049 59666 394115 59669
rect 423029 59666 423095 59669
rect 452101 59666 452167 59669
rect 481081 59666 481147 59669
rect 510061 59666 510127 59669
rect 539041 59666 539107 59669
rect 567377 59666 567443 59669
rect 246652 59664 249123 59666
rect 217734 59394 217794 59636
rect 246652 59608 249062 59664
rect 249118 59608 249123 59664
rect 246652 59606 249123 59608
rect 275724 59664 278195 59666
rect 275724 59608 278134 59664
rect 278190 59608 278195 59664
rect 275724 59606 278195 59608
rect 304612 59664 307175 59666
rect 304612 59608 307114 59664
rect 307170 59608 307175 59664
rect 304612 59606 307175 59608
rect 333684 59664 336155 59666
rect 333684 59608 336094 59664
rect 336150 59608 336155 59664
rect 333684 59606 336155 59608
rect 362756 59664 365135 59666
rect 362756 59608 365074 59664
rect 365130 59608 365135 59664
rect 362756 59606 365135 59608
rect 391644 59664 394115 59666
rect 391644 59608 394054 59664
rect 394110 59608 394115 59664
rect 391644 59606 394115 59608
rect 420716 59664 423095 59666
rect 420716 59608 423034 59664
rect 423090 59608 423095 59664
rect 420716 59606 423095 59608
rect 449604 59664 452167 59666
rect 449604 59608 452106 59664
rect 452162 59608 452167 59664
rect 449604 59606 452167 59608
rect 478676 59664 481147 59666
rect 478676 59608 481086 59664
rect 481142 59608 481147 59664
rect 478676 59606 481147 59608
rect 507748 59664 510127 59666
rect 507748 59608 510066 59664
rect 510122 59608 510127 59664
rect 507748 59606 510127 59608
rect 536636 59664 539107 59666
rect 536636 59608 539046 59664
rect 539102 59608 539107 59664
rect 536636 59606 539107 59608
rect 565708 59664 567443 59666
rect 565708 59608 567382 59664
rect 567438 59608 567443 59664
rect 565708 59606 567443 59608
rect 249057 59603 249123 59606
rect 278129 59603 278195 59606
rect 307109 59603 307175 59606
rect 336089 59603 336155 59606
rect 365069 59603 365135 59606
rect 394049 59603 394115 59606
rect 423029 59603 423095 59606
rect 452101 59603 452167 59606
rect 481081 59603 481147 59606
rect 510061 59603 510127 59606
rect 539041 59603 539107 59606
rect 567377 59603 567443 59606
rect 583520 59516 584960 59756
rect 220169 59394 220235 59397
rect 217734 59392 220235 59394
rect 217734 59336 220174 59392
rect 220230 59336 220235 59392
rect 217734 59334 220235 59336
rect 220169 59331 220235 59334
rect 265758 58926 269866 58986
rect 207828 58790 211876 58850
rect 236900 58790 240948 58850
rect 265758 58820 265818 58926
rect 269806 58820 269866 58926
rect 410934 58926 415042 58986
rect 294860 58790 298908 58850
rect 323932 58790 327980 58850
rect 352820 58790 356868 58850
rect 381892 58790 385940 58850
rect 410934 58820 410994 58926
rect 414982 58820 415042 58926
rect 439852 58790 443900 58850
rect 468924 58790 472972 58850
rect 497812 58790 501860 58850
rect 526884 58790 530932 58850
rect 555956 58790 560004 58850
rect -960 58578 480 58668
rect 3325 58578 3391 58581
rect -960 58576 3391 58578
rect -960 58520 3330 58576
rect 3386 58520 3391 58576
rect -960 58518 3391 58520
rect -960 58428 480 58518
rect 3325 58515 3391 58518
rect 265758 57430 269866 57490
rect 207828 57294 211876 57354
rect 236900 57294 240948 57354
rect 265758 57324 265818 57430
rect 269806 57324 269866 57430
rect 410934 57430 415042 57490
rect 294860 57294 298908 57354
rect 323932 57294 327980 57354
rect 352820 57294 356868 57354
rect 381892 57294 385940 57354
rect 410934 57324 410994 57430
rect 414982 57324 415042 57430
rect 439852 57294 443900 57354
rect 468924 57294 472972 57354
rect 497812 57294 501860 57354
rect 526884 57294 530932 57354
rect 555956 57294 560004 57354
rect 220353 56810 220419 56813
rect 217734 56808 220419 56810
rect 217734 56752 220358 56808
rect 220414 56752 220419 56808
rect 217734 56750 220419 56752
rect 217734 56644 217794 56750
rect 220353 56747 220419 56750
rect 249241 56674 249307 56677
rect 278221 56674 278287 56677
rect 307201 56674 307267 56677
rect 336181 56674 336247 56677
rect 365161 56674 365227 56677
rect 394141 56674 394207 56677
rect 423121 56674 423187 56677
rect 452193 56674 452259 56677
rect 481173 56674 481239 56677
rect 510153 56674 510219 56677
rect 539133 56674 539199 56677
rect 567469 56674 567535 56677
rect 246652 56672 249307 56674
rect 246652 56616 249246 56672
rect 249302 56616 249307 56672
rect 246652 56614 249307 56616
rect 275724 56672 278287 56674
rect 275724 56616 278226 56672
rect 278282 56616 278287 56672
rect 275724 56614 278287 56616
rect 304612 56672 307267 56674
rect 304612 56616 307206 56672
rect 307262 56616 307267 56672
rect 304612 56614 307267 56616
rect 333684 56672 336247 56674
rect 333684 56616 336186 56672
rect 336242 56616 336247 56672
rect 333684 56614 336247 56616
rect 362756 56672 365227 56674
rect 362756 56616 365166 56672
rect 365222 56616 365227 56672
rect 362756 56614 365227 56616
rect 391644 56672 394207 56674
rect 391644 56616 394146 56672
rect 394202 56616 394207 56672
rect 391644 56614 394207 56616
rect 420716 56672 423187 56674
rect 420716 56616 423126 56672
rect 423182 56616 423187 56672
rect 420716 56614 423187 56616
rect 449604 56672 452259 56674
rect 449604 56616 452198 56672
rect 452254 56616 452259 56672
rect 449604 56614 452259 56616
rect 478676 56672 481239 56674
rect 478676 56616 481178 56672
rect 481234 56616 481239 56672
rect 478676 56614 481239 56616
rect 507748 56672 510219 56674
rect 507748 56616 510158 56672
rect 510214 56616 510219 56672
rect 507748 56614 510219 56616
rect 536636 56672 539199 56674
rect 536636 56616 539138 56672
rect 539194 56616 539199 56672
rect 536636 56614 539199 56616
rect 565708 56672 567535 56674
rect 565708 56616 567474 56672
rect 567530 56616 567535 56672
rect 565708 56614 567535 56616
rect 249241 56611 249307 56614
rect 278221 56611 278287 56614
rect 307201 56611 307267 56614
rect 336181 56611 336247 56614
rect 365161 56611 365227 56614
rect 394141 56611 394207 56614
rect 423121 56611 423187 56614
rect 452193 56611 452259 56614
rect 481173 56611 481239 56614
rect 510153 56611 510219 56614
rect 539133 56611 539199 56614
rect 567469 56611 567535 56614
rect 265758 55934 269866 55994
rect 207828 55798 211876 55858
rect 236900 55798 240948 55858
rect 265758 55828 265818 55934
rect 269806 55828 269866 55934
rect 410934 55934 415042 55994
rect 294860 55798 298908 55858
rect 323932 55798 327980 55858
rect 352820 55798 356868 55858
rect 381892 55798 385940 55858
rect 410934 55828 410994 55934
rect 414982 55828 415042 55934
rect 439852 55798 443900 55858
rect 468924 55798 472972 55858
rect 497812 55798 501860 55858
rect 526884 55798 530932 55858
rect 555956 55798 560004 55858
rect 265758 54438 269866 54498
rect 207828 54302 211876 54362
rect 236900 54302 240948 54362
rect 265758 54332 265818 54438
rect 269806 54332 269866 54438
rect 410934 54438 415042 54498
rect 294860 54302 298908 54362
rect 323932 54302 327980 54362
rect 352820 54302 356868 54362
rect 381892 54302 385940 54362
rect 410934 54332 410994 54438
rect 414982 54332 415042 54438
rect 439852 54302 443900 54362
rect 468924 54302 472972 54362
rect 497812 54302 501860 54362
rect 526884 54302 530932 54362
rect 555956 54302 560004 54362
rect 248413 53682 248479 53685
rect 277393 53682 277459 53685
rect 306557 53682 306623 53685
rect 335353 53682 335419 53685
rect 364333 53682 364399 53685
rect 393313 53682 393379 53685
rect 422293 53682 422359 53685
rect 451457 53682 451523 53685
rect 480437 53682 480503 53685
rect 509417 53682 509483 53685
rect 538397 53682 538463 53685
rect 567561 53682 567627 53685
rect 246652 53680 248479 53682
rect 246652 53624 248418 53680
rect 248474 53624 248479 53680
rect 246652 53622 248479 53624
rect 275724 53680 277459 53682
rect 275724 53624 277398 53680
rect 277454 53624 277459 53680
rect 275724 53622 277459 53624
rect 304612 53680 306623 53682
rect 304612 53624 306562 53680
rect 306618 53624 306623 53680
rect 304612 53622 306623 53624
rect 333684 53680 335419 53682
rect 333684 53624 335358 53680
rect 335414 53624 335419 53680
rect 333684 53622 335419 53624
rect 362756 53680 364399 53682
rect 362756 53624 364338 53680
rect 364394 53624 364399 53680
rect 362756 53622 364399 53624
rect 391644 53680 393379 53682
rect 391644 53624 393318 53680
rect 393374 53624 393379 53680
rect 391644 53622 393379 53624
rect 420716 53680 422359 53682
rect 420716 53624 422298 53680
rect 422354 53624 422359 53680
rect 420716 53622 422359 53624
rect 449604 53680 451523 53682
rect 449604 53624 451462 53680
rect 451518 53624 451523 53680
rect 449604 53622 451523 53624
rect 478676 53680 480503 53682
rect 478676 53624 480442 53680
rect 480498 53624 480503 53680
rect 478676 53622 480503 53624
rect 507748 53680 509483 53682
rect 507748 53624 509422 53680
rect 509478 53624 509483 53680
rect 507748 53622 509483 53624
rect 536636 53680 538463 53682
rect 536636 53624 538402 53680
rect 538458 53624 538463 53680
rect 536636 53622 538463 53624
rect 565708 53680 567627 53682
rect 565708 53624 567566 53680
rect 567622 53624 567627 53680
rect 565708 53622 567627 53624
rect 248413 53619 248479 53622
rect 277393 53619 277459 53622
rect 306557 53619 306623 53622
rect 335353 53619 335419 53622
rect 364333 53619 364399 53622
rect 393313 53619 393379 53622
rect 422293 53619 422359 53622
rect 451457 53619 451523 53622
rect 480437 53619 480503 53622
rect 509417 53619 509483 53622
rect 538397 53619 538463 53622
rect 567561 53619 567627 53622
rect 265758 52942 269866 53002
rect 207828 52806 211876 52866
rect 236900 52806 240948 52866
rect 265758 52836 265818 52942
rect 269806 52836 269866 52942
rect 410934 52942 415042 53002
rect 294860 52806 298908 52866
rect 323932 52806 327980 52866
rect 352820 52806 356868 52866
rect 381892 52806 385940 52866
rect 410934 52836 410994 52942
rect 414982 52836 415042 52942
rect 439852 52806 443900 52866
rect 468924 52806 472972 52866
rect 497812 52806 501860 52866
rect 526884 52806 530932 52866
rect 555956 52806 560004 52866
rect 265758 51446 269866 51506
rect 207828 51310 211876 51370
rect 236900 51310 240948 51370
rect 265758 51340 265818 51446
rect 269806 51340 269866 51446
rect 410934 51446 415042 51506
rect 294860 51310 298908 51370
rect 323932 51310 327980 51370
rect 352820 51310 356868 51370
rect 381892 51310 385940 51370
rect 410934 51340 410994 51446
rect 414982 51340 415042 51446
rect 439852 51310 443900 51370
rect 468924 51310 472972 51370
rect 497812 51310 501860 51370
rect 526884 51310 530932 51370
rect 555956 51310 560004 51370
rect 248505 50690 248571 50693
rect 277485 50690 277551 50693
rect 306465 50690 306531 50693
rect 335445 50690 335511 50693
rect 364425 50690 364491 50693
rect 393405 50690 393471 50693
rect 422385 50690 422451 50693
rect 451365 50690 451431 50693
rect 480345 50690 480411 50693
rect 509325 50690 509391 50693
rect 538305 50690 538371 50693
rect 567653 50690 567719 50693
rect 246652 50688 248571 50690
rect 246652 50632 248510 50688
rect 248566 50632 248571 50688
rect 246652 50630 248571 50632
rect 275724 50688 277551 50690
rect 275724 50632 277490 50688
rect 277546 50632 277551 50688
rect 275724 50630 277551 50632
rect 304612 50688 306531 50690
rect 304612 50632 306470 50688
rect 306526 50632 306531 50688
rect 304612 50630 306531 50632
rect 333684 50688 335511 50690
rect 333684 50632 335450 50688
rect 335506 50632 335511 50688
rect 333684 50630 335511 50632
rect 362756 50688 364491 50690
rect 362756 50632 364430 50688
rect 364486 50632 364491 50688
rect 362756 50630 364491 50632
rect 391644 50688 393471 50690
rect 391644 50632 393410 50688
rect 393466 50632 393471 50688
rect 391644 50630 393471 50632
rect 420716 50688 422451 50690
rect 420716 50632 422390 50688
rect 422446 50632 422451 50688
rect 420716 50630 422451 50632
rect 449604 50688 451431 50690
rect 449604 50632 451370 50688
rect 451426 50632 451431 50688
rect 449604 50630 451431 50632
rect 478676 50688 480411 50690
rect 478676 50632 480350 50688
rect 480406 50632 480411 50688
rect 478676 50630 480411 50632
rect 507748 50688 509391 50690
rect 507748 50632 509330 50688
rect 509386 50632 509391 50688
rect 507748 50630 509391 50632
rect 536636 50688 538371 50690
rect 536636 50632 538310 50688
rect 538366 50632 538371 50688
rect 536636 50630 538371 50632
rect 565708 50688 567719 50690
rect 565708 50632 567658 50688
rect 567714 50632 567719 50688
rect 565708 50630 567719 50632
rect 248505 50627 248571 50630
rect 277485 50627 277551 50630
rect 306465 50627 306531 50630
rect 335445 50627 335511 50630
rect 364425 50627 364491 50630
rect 393405 50627 393471 50630
rect 422385 50627 422451 50630
rect 451365 50627 451431 50630
rect 480345 50627 480411 50630
rect 509325 50627 509391 50630
rect 538305 50627 538371 50630
rect 567653 50627 567719 50630
rect 265758 49950 269866 50010
rect 207828 49814 211876 49874
rect 236900 49814 240948 49874
rect 265758 49844 265818 49950
rect 269806 49844 269866 49950
rect 410934 49950 415042 50010
rect 294860 49814 298908 49874
rect 323932 49814 327980 49874
rect 352820 49814 356868 49874
rect 381892 49814 385940 49874
rect 410934 49844 410994 49950
rect 414982 49844 415042 49950
rect 439852 49814 443900 49874
rect 468924 49814 472972 49874
rect 497812 49814 501860 49874
rect 526884 49814 530932 49874
rect 555956 49814 560004 49874
rect 265758 48454 269866 48514
rect 207828 48318 211876 48378
rect 236900 48318 240948 48378
rect 265758 48348 265818 48454
rect 269806 48348 269866 48454
rect 410934 48454 415042 48514
rect 294860 48318 298908 48378
rect 323932 48318 327980 48378
rect 352820 48318 356868 48378
rect 381892 48318 385940 48378
rect 410934 48348 410994 48454
rect 414982 48348 415042 48454
rect 439852 48318 443900 48378
rect 468924 48318 472972 48378
rect 497812 48318 501860 48378
rect 526884 48318 530932 48378
rect 555956 48318 560004 48378
rect 480253 47698 480319 47701
rect 509233 47698 509299 47701
rect 538213 47698 538279 47701
rect 567193 47698 567259 47701
rect 478676 47696 480319 47698
rect 217734 47154 217794 47668
rect 246070 47157 246130 47668
rect 275142 47157 275202 47668
rect 219433 47154 219499 47157
rect 217734 47152 219499 47154
rect 217734 47096 219438 47152
rect 219494 47096 219499 47152
rect 217734 47094 219499 47096
rect 246070 47152 246179 47157
rect 246070 47096 246118 47152
rect 246174 47096 246179 47152
rect 246070 47094 246179 47096
rect 219433 47091 219499 47094
rect 246113 47091 246179 47094
rect 275093 47152 275202 47157
rect 275093 47096 275098 47152
rect 275154 47096 275202 47152
rect 275093 47094 275202 47096
rect 304073 47154 304139 47157
rect 304214 47154 304274 47668
rect 304073 47152 304274 47154
rect 304073 47096 304078 47152
rect 304134 47096 304274 47152
rect 304073 47094 304274 47096
rect 333102 47157 333162 47668
rect 362174 47157 362234 47668
rect 333102 47152 333211 47157
rect 333102 47096 333150 47152
rect 333206 47096 333211 47152
rect 333102 47094 333211 47096
rect 275093 47091 275159 47094
rect 304073 47091 304139 47094
rect 333145 47091 333211 47094
rect 362125 47152 362234 47157
rect 362125 47096 362130 47152
rect 362186 47096 362234 47152
rect 362125 47094 362234 47096
rect 391062 47157 391122 47668
rect 420134 47157 420194 47668
rect 391062 47152 391171 47157
rect 391062 47096 391110 47152
rect 391166 47096 391171 47152
rect 391062 47094 391171 47096
rect 362125 47091 362191 47094
rect 391105 47091 391171 47094
rect 420085 47152 420194 47157
rect 420085 47096 420090 47152
rect 420146 47096 420194 47152
rect 420085 47094 420194 47096
rect 449065 47154 449131 47157
rect 449206 47154 449266 47668
rect 478676 47640 480258 47696
rect 480314 47640 480319 47696
rect 478676 47638 480319 47640
rect 507748 47696 509299 47698
rect 507748 47640 509238 47696
rect 509294 47640 509299 47696
rect 507748 47638 509299 47640
rect 536636 47696 538279 47698
rect 536636 47640 538218 47696
rect 538274 47640 538279 47696
rect 536636 47638 538279 47640
rect 565708 47696 567259 47698
rect 565708 47640 567198 47696
rect 567254 47640 567259 47696
rect 565708 47638 567259 47640
rect 480253 47635 480319 47638
rect 509233 47635 509299 47638
rect 538213 47635 538279 47638
rect 567193 47635 567259 47638
rect 449065 47152 449266 47154
rect 449065 47096 449070 47152
rect 449126 47096 449266 47152
rect 449065 47094 449266 47096
rect 420085 47091 420151 47094
rect 449065 47091 449131 47094
rect 207828 46822 211876 46882
rect 236900 46822 240948 46882
rect 265758 46746 265818 46852
rect 269806 46746 269866 46852
rect 294860 46822 298908 46882
rect 323932 46822 327980 46882
rect 352820 46822 356868 46882
rect 381892 46822 385940 46882
rect 265758 46686 269866 46746
rect 410934 46746 410994 46852
rect 414982 46746 415042 46852
rect 439852 46822 443900 46882
rect 468924 46822 472972 46882
rect 497812 46822 501860 46882
rect 526884 46822 530932 46882
rect 555956 46822 560004 46882
rect 410934 46686 415042 46746
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 3233 45522 3299 45525
rect -960 45520 3299 45522
rect -960 45464 3238 45520
rect 3294 45464 3299 45520
rect -960 45462 3299 45464
rect -960 45372 480 45462
rect 3233 45459 3299 45462
rect 265758 45462 269866 45522
rect 207828 45326 211876 45386
rect 236900 45326 240948 45386
rect 265758 45356 265818 45462
rect 269806 45356 269866 45462
rect 410934 45462 415042 45522
rect 294860 45326 298908 45386
rect 323932 45326 327980 45386
rect 352820 45326 356868 45386
rect 381892 45326 385940 45386
rect 410934 45356 410994 45462
rect 414982 45356 415042 45462
rect 439852 45326 443900 45386
rect 468924 45326 472972 45386
rect 497812 45326 501860 45386
rect 526884 45326 530932 45386
rect 555956 45326 560004 45386
rect 217182 44165 217242 44676
rect 217133 44160 217242 44165
rect 217133 44104 217138 44160
rect 217194 44104 217242 44160
rect 217133 44102 217242 44104
rect 217133 44099 217199 44102
rect 207828 43830 211876 43890
rect 236900 43830 240948 43890
rect 220261 43618 220327 43621
rect 245929 43618 245995 43621
rect 220261 43616 245995 43618
rect 220261 43560 220266 43616
rect 220322 43560 245934 43616
rect 245990 43560 245995 43616
rect 220261 43558 245995 43560
rect 220261 43555 220327 43558
rect 245929 43555 245995 43558
rect 220077 43346 220143 43349
rect 246070 43346 246130 44676
rect 265758 43966 269866 44026
rect 265758 43860 265818 43966
rect 269806 43860 269866 43966
rect 249149 43618 249215 43621
rect 275001 43618 275067 43621
rect 249149 43616 275067 43618
rect 249149 43560 249154 43616
rect 249210 43560 275006 43616
rect 275062 43560 275067 43616
rect 249149 43558 275067 43560
rect 249149 43555 249215 43558
rect 275001 43555 275067 43558
rect 220077 43344 246130 43346
rect 220077 43288 220082 43344
rect 220138 43288 246130 43344
rect 220077 43286 246130 43288
rect 220077 43283 220143 43286
rect 249006 43284 249012 43348
rect 249076 43346 249082 43348
rect 275142 43346 275202 44676
rect 294860 43830 298908 43890
rect 277894 43556 277900 43620
rect 277964 43618 277970 43620
rect 304214 43618 304274 44676
rect 323932 43830 327980 43890
rect 277964 43558 304274 43618
rect 277964 43556 277970 43558
rect 306966 43556 306972 43620
rect 307036 43618 307042 43620
rect 333102 43618 333162 44676
rect 352820 43830 356868 43890
rect 307036 43558 333162 43618
rect 307036 43556 307042 43558
rect 335854 43556 335860 43620
rect 335924 43618 335930 43620
rect 362174 43618 362234 44676
rect 381892 43830 385940 43890
rect 335924 43558 362234 43618
rect 335924 43556 335930 43558
rect 364926 43556 364932 43620
rect 364996 43618 365002 43620
rect 391062 43618 391122 44676
rect 410934 43966 415042 44026
rect 410934 43860 410994 43966
rect 414982 43860 415042 43966
rect 364996 43558 391122 43618
rect 364996 43556 365002 43558
rect 393814 43556 393820 43620
rect 393884 43618 393890 43620
rect 420134 43618 420194 44676
rect 439852 43830 443900 43890
rect 393884 43558 420194 43618
rect 393884 43556 393890 43558
rect 422886 43556 422892 43620
rect 422956 43618 422962 43620
rect 449206 43618 449266 44676
rect 468924 43830 472972 43890
rect 422956 43558 449266 43618
rect 451917 43618 451983 43621
rect 478094 43618 478154 44676
rect 497812 43830 501860 43890
rect 451917 43616 478154 43618
rect 451917 43560 451922 43616
rect 451978 43560 478154 43616
rect 451917 43558 478154 43560
rect 480897 43618 480963 43621
rect 507166 43618 507226 44676
rect 526884 43830 530932 43890
rect 480897 43616 507226 43618
rect 480897 43560 480902 43616
rect 480958 43560 507226 43616
rect 480897 43558 507226 43560
rect 509877 43618 509943 43621
rect 536238 43618 536298 44676
rect 565126 44165 565186 44676
rect 565077 44160 565186 44165
rect 565077 44104 565082 44160
rect 565138 44104 565186 44160
rect 565077 44102 565186 44104
rect 565077 44099 565143 44102
rect 555956 43830 560004 43890
rect 509877 43616 536298 43618
rect 509877 43560 509882 43616
rect 509938 43560 536298 43616
rect 509877 43558 536298 43560
rect 422956 43556 422962 43558
rect 451917 43555 451983 43558
rect 480897 43555 480963 43558
rect 509877 43555 509943 43558
rect 249076 43286 275202 43346
rect 249076 43284 249082 43286
rect 13537 39402 13603 39405
rect 217133 39402 217199 39405
rect 13537 39400 217199 39402
rect 13537 39344 13542 39400
rect 13598 39344 217138 39400
rect 217194 39344 217199 39400
rect 13537 39342 217199 39344
rect 13537 39339 13603 39342
rect 217133 39339 217199 39342
rect 456934 39342 458282 39402
rect 79918 39130 79978 39236
rect 81206 39130 81266 39236
rect 108836 39206 110308 39266
rect 137908 39206 139380 39266
rect 166796 39206 168268 39266
rect 195868 39206 197340 39266
rect 224940 39206 226412 39266
rect 253828 39206 255300 39266
rect 282900 39206 284372 39266
rect 311788 39206 313260 39266
rect 340860 39206 342332 39266
rect 369932 39206 371404 39266
rect 398820 39206 400292 39266
rect 427892 39206 429364 39266
rect 456934 39236 456994 39342
rect 458222 39236 458282 39342
rect 485852 39206 487324 39266
rect 514924 39206 516396 39266
rect 543812 39206 545284 39266
rect 79918 39070 81266 39130
rect 538121 38586 538187 38589
rect 538078 38584 538187 38586
rect 538078 38528 538126 38584
rect 538182 38528 538187 38584
rect 538078 38523 538187 38528
rect 71681 38450 71747 38453
rect 100661 38450 100727 38453
rect 129365 38450 129431 38453
rect 158345 38450 158411 38453
rect 187325 38450 187391 38453
rect 216305 38450 216371 38453
rect 246665 38450 246731 38453
rect 275645 38450 275711 38453
rect 304625 38450 304691 38453
rect 333605 38450 333671 38453
rect 362585 38450 362651 38453
rect 391565 38450 391631 38453
rect 420545 38450 420611 38453
rect 449525 38450 449591 38453
rect 478505 38450 478571 38453
rect 71681 38448 74060 38450
rect 71681 38392 71686 38448
rect 71742 38392 74060 38448
rect 71681 38390 74060 38392
rect 100661 38448 103132 38450
rect 100661 38392 100666 38448
rect 100722 38392 103132 38448
rect 100661 38390 103132 38392
rect 129365 38448 132204 38450
rect 129365 38392 129370 38448
rect 129426 38392 132204 38448
rect 129365 38390 132204 38392
rect 158345 38448 161092 38450
rect 158345 38392 158350 38448
rect 158406 38392 161092 38448
rect 158345 38390 161092 38392
rect 187325 38448 190164 38450
rect 187325 38392 187330 38448
rect 187386 38392 190164 38448
rect 187325 38390 190164 38392
rect 216305 38448 219052 38450
rect 216305 38392 216310 38448
rect 216366 38392 219052 38448
rect 216305 38390 219052 38392
rect 246665 38448 248124 38450
rect 246665 38392 246670 38448
rect 246726 38392 248124 38448
rect 246665 38390 248124 38392
rect 275645 38448 277196 38450
rect 275645 38392 275650 38448
rect 275706 38392 277196 38448
rect 275645 38390 277196 38392
rect 304625 38448 306084 38450
rect 304625 38392 304630 38448
rect 304686 38392 306084 38448
rect 304625 38390 306084 38392
rect 333605 38448 335156 38450
rect 333605 38392 333610 38448
rect 333666 38392 335156 38448
rect 333605 38390 335156 38392
rect 362585 38448 364044 38450
rect 362585 38392 362590 38448
rect 362646 38392 364044 38448
rect 362585 38390 364044 38392
rect 391565 38448 393116 38450
rect 391565 38392 391570 38448
rect 391626 38392 393116 38448
rect 391565 38390 393116 38392
rect 420545 38448 422188 38450
rect 420545 38392 420550 38448
rect 420606 38392 422188 38448
rect 420545 38390 422188 38392
rect 449525 38448 451076 38450
rect 449525 38392 449530 38448
rect 449586 38392 451076 38448
rect 449525 38390 451076 38392
rect 478505 38448 480148 38450
rect 478505 38392 478510 38448
rect 478566 38392 480148 38448
rect 538078 38420 538138 38523
rect 478505 38390 480148 38392
rect 71681 38387 71747 38390
rect 100661 38387 100727 38390
rect 129365 38387 129431 38390
rect 158345 38387 158411 38390
rect 187325 38387 187391 38390
rect 216305 38387 216371 38390
rect 246665 38387 246731 38390
rect 275645 38387 275711 38390
rect 304625 38387 304691 38390
rect 333605 38387 333671 38390
rect 362585 38387 362651 38390
rect 391565 38387 391631 38390
rect 420545 38387 420611 38390
rect 449525 38387 449591 38390
rect 478505 38387 478571 38390
rect 3366 37844 3372 37908
rect 3436 37906 3442 37908
rect 54661 37906 54727 37909
rect 507485 37906 507551 37909
rect 509006 37906 509066 38420
rect 3436 37904 54727 37906
rect 3436 37848 54666 37904
rect 54722 37848 54727 37904
rect 3436 37846 54727 37848
rect 3436 37844 3442 37846
rect 54661 37843 54727 37846
rect 79918 37846 81266 37906
rect 79918 37740 79978 37846
rect 81206 37740 81266 37846
rect 456934 37846 458282 37906
rect 108836 37710 110308 37770
rect 137908 37710 139380 37770
rect 166796 37710 168268 37770
rect 195868 37710 197340 37770
rect 224940 37710 226412 37770
rect 253828 37710 255300 37770
rect 282900 37710 284372 37770
rect 311788 37710 313260 37770
rect 340860 37710 342332 37770
rect 369932 37710 371404 37770
rect 398820 37710 400292 37770
rect 427892 37710 429364 37770
rect 456934 37740 456994 37846
rect 458222 37740 458282 37846
rect 507485 37904 509066 37906
rect 507485 37848 507490 37904
rect 507546 37848 509066 37904
rect 507485 37846 509066 37848
rect 507485 37843 507551 37846
rect 485852 37710 487324 37770
rect 514924 37710 516396 37770
rect 543812 37710 545284 37770
rect 79918 36350 81266 36410
rect 79918 36244 79978 36350
rect 81206 36244 81266 36350
rect 456934 36350 458282 36410
rect 108836 36214 110308 36274
rect 137908 36214 139380 36274
rect 166796 36214 168268 36274
rect 195868 36214 197340 36274
rect 224940 36214 226412 36274
rect 253828 36214 255300 36274
rect 282900 36214 284372 36274
rect 311788 36214 313260 36274
rect 340860 36214 342332 36274
rect 369932 36214 371404 36274
rect 398820 36214 400292 36274
rect 427892 36214 429364 36274
rect 456934 36244 456994 36350
rect 458222 36244 458282 36350
rect 485852 36214 487324 36274
rect 514924 36214 516396 36274
rect 543812 36214 545284 36274
rect 71589 35458 71655 35461
rect 100569 35458 100635 35461
rect 129549 35458 129615 35461
rect 158529 35458 158595 35461
rect 187509 35458 187575 35461
rect 216489 35458 216555 35461
rect 246849 35458 246915 35461
rect 275829 35458 275895 35461
rect 304809 35458 304875 35461
rect 333789 35458 333855 35461
rect 362769 35458 362835 35461
rect 391749 35458 391815 35461
rect 420729 35458 420795 35461
rect 449709 35458 449775 35461
rect 478689 35458 478755 35461
rect 536557 35458 536623 35461
rect 71589 35456 74060 35458
rect 71589 35400 71594 35456
rect 71650 35400 74060 35456
rect 71589 35398 74060 35400
rect 100569 35456 103132 35458
rect 100569 35400 100574 35456
rect 100630 35400 103132 35456
rect 100569 35398 103132 35400
rect 129549 35456 132204 35458
rect 129549 35400 129554 35456
rect 129610 35400 132204 35456
rect 129549 35398 132204 35400
rect 158529 35456 161092 35458
rect 158529 35400 158534 35456
rect 158590 35400 161092 35456
rect 158529 35398 161092 35400
rect 187509 35456 190164 35458
rect 187509 35400 187514 35456
rect 187570 35400 190164 35456
rect 187509 35398 190164 35400
rect 216489 35456 219052 35458
rect 216489 35400 216494 35456
rect 216550 35400 219052 35456
rect 216489 35398 219052 35400
rect 246849 35456 248124 35458
rect 246849 35400 246854 35456
rect 246910 35400 248124 35456
rect 246849 35398 248124 35400
rect 275829 35456 277196 35458
rect 275829 35400 275834 35456
rect 275890 35400 277196 35456
rect 275829 35398 277196 35400
rect 304809 35456 306084 35458
rect 304809 35400 304814 35456
rect 304870 35400 306084 35456
rect 304809 35398 306084 35400
rect 333789 35456 335156 35458
rect 333789 35400 333794 35456
rect 333850 35400 335156 35456
rect 333789 35398 335156 35400
rect 362769 35456 364044 35458
rect 362769 35400 362774 35456
rect 362830 35400 364044 35456
rect 362769 35398 364044 35400
rect 391749 35456 393116 35458
rect 391749 35400 391754 35456
rect 391810 35400 393116 35456
rect 391749 35398 393116 35400
rect 420729 35456 422188 35458
rect 420729 35400 420734 35456
rect 420790 35400 422188 35456
rect 420729 35398 422188 35400
rect 449709 35456 451076 35458
rect 449709 35400 449714 35456
rect 449770 35400 451076 35456
rect 449709 35398 451076 35400
rect 478689 35456 480148 35458
rect 478689 35400 478694 35456
rect 478750 35400 480148 35456
rect 536557 35456 538108 35458
rect 478689 35398 480148 35400
rect 71589 35395 71655 35398
rect 100569 35395 100635 35398
rect 129549 35395 129615 35398
rect 158529 35395 158595 35398
rect 187509 35395 187575 35398
rect 216489 35395 216555 35398
rect 246849 35395 246915 35398
rect 275829 35395 275895 35398
rect 304809 35395 304875 35398
rect 333789 35395 333855 35398
rect 362769 35395 362835 35398
rect 391749 35395 391815 35398
rect 420729 35395 420795 35398
rect 449709 35395 449775 35398
rect 478689 35395 478755 35398
rect 39665 35322 39731 35325
rect 39798 35322 39804 35324
rect 39665 35320 39804 35322
rect 39665 35264 39670 35320
rect 39726 35264 39804 35320
rect 39665 35262 39804 35264
rect 39665 35259 39731 35262
rect 39798 35260 39804 35262
rect 39868 35260 39874 35324
rect 42742 35260 42748 35324
rect 42812 35322 42818 35324
rect 43437 35322 43503 35325
rect 42812 35320 43503 35322
rect 42812 35264 43442 35320
rect 43498 35264 43503 35320
rect 42812 35262 43503 35264
rect 42812 35260 42818 35262
rect 43437 35259 43503 35262
rect 50521 35322 50587 35325
rect 50838 35322 50844 35324
rect 50521 35320 50844 35322
rect 50521 35264 50526 35320
rect 50582 35264 50844 35320
rect 50521 35262 50844 35264
rect 50521 35259 50587 35262
rect 50838 35260 50844 35262
rect 50908 35260 50914 35324
rect 64505 35186 64571 35189
rect 61916 35184 64571 35186
rect 61916 35128 64510 35184
rect 64566 35128 64571 35184
rect 61916 35126 64571 35128
rect 64505 35123 64571 35126
rect 507669 34914 507735 34917
rect 509006 34914 509066 35428
rect 536557 35400 536562 35456
rect 536618 35400 538108 35456
rect 536557 35398 538108 35400
rect 536557 35395 536623 35398
rect 79918 34854 81266 34914
rect 79918 34748 79978 34854
rect 81206 34748 81266 34854
rect 456934 34854 458282 34914
rect 108836 34718 110308 34778
rect 137908 34718 139380 34778
rect 166796 34718 168268 34778
rect 195868 34718 197340 34778
rect 224940 34718 226412 34778
rect 253828 34718 255300 34778
rect 282900 34718 284372 34778
rect 311788 34718 313260 34778
rect 340860 34718 342332 34778
rect 369932 34718 371404 34778
rect 398820 34718 400292 34778
rect 427892 34718 429364 34778
rect 456934 34748 456994 34854
rect 458222 34748 458282 34854
rect 507669 34912 509066 34914
rect 507669 34856 507674 34912
rect 507730 34856 509066 34912
rect 507669 34854 509066 34856
rect 507669 34851 507735 34854
rect 485852 34718 487324 34778
rect 514924 34718 516396 34778
rect 543812 34718 545284 34778
rect 12433 34506 12499 34509
rect 12433 34504 16100 34506
rect 12433 34448 12438 34504
rect 12494 34448 16100 34504
rect 12433 34446 16100 34448
rect 12433 34443 12499 34446
rect 61285 34370 61351 34373
rect 61285 34368 61394 34370
rect 61285 34312 61290 34368
rect 61346 34312 61394 34368
rect 61285 34307 61394 34312
rect 61334 33796 61394 34307
rect 79918 33358 81266 33418
rect 79918 33252 79978 33358
rect 81206 33252 81266 33358
rect 456934 33358 458282 33418
rect 108836 33222 110308 33282
rect 137908 33222 139380 33282
rect 166796 33222 168268 33282
rect 195868 33222 197340 33282
rect 224940 33222 226412 33282
rect 253828 33222 255300 33282
rect 282900 33222 284372 33282
rect 311788 33222 313260 33282
rect 340860 33222 342332 33282
rect 369932 33222 371404 33282
rect 398820 33222 400292 33282
rect 427892 33222 429364 33282
rect 456934 33252 456994 33358
rect 458222 33252 458282 33358
rect 485852 33222 487324 33282
rect 514924 33222 516396 33282
rect 543812 33222 545284 33282
rect 13721 33146 13787 33149
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 13721 33144 16100 33146
rect 13721 33088 13726 33144
rect 13782 33088 16100 33144
rect 13721 33086 16100 33088
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 13721 33083 13787 33086
rect 580165 33083 580231 33086
rect 507761 33010 507827 33013
rect 507761 33008 509066 33010
rect 507761 32952 507766 33008
rect 507822 32952 509066 33008
rect 583520 32996 584960 33086
rect 507761 32950 509066 32952
rect 507761 32947 507827 32950
rect -960 32316 480 32556
rect 71405 32466 71471 32469
rect 100385 32466 100451 32469
rect 129641 32466 129707 32469
rect 158621 32466 158687 32469
rect 187601 32466 187667 32469
rect 216581 32466 216647 32469
rect 246941 32466 247007 32469
rect 275921 32466 275987 32469
rect 304901 32466 304967 32469
rect 333881 32466 333947 32469
rect 362861 32466 362927 32469
rect 391841 32466 391907 32469
rect 420821 32466 420887 32469
rect 449801 32466 449867 32469
rect 478781 32466 478847 32469
rect 71405 32464 74060 32466
rect 71405 32408 71410 32464
rect 71466 32408 74060 32464
rect 71405 32406 74060 32408
rect 100385 32464 103132 32466
rect 100385 32408 100390 32464
rect 100446 32408 103132 32464
rect 100385 32406 103132 32408
rect 129641 32464 132204 32466
rect 129641 32408 129646 32464
rect 129702 32408 132204 32464
rect 129641 32406 132204 32408
rect 158621 32464 161092 32466
rect 158621 32408 158626 32464
rect 158682 32408 161092 32464
rect 158621 32406 161092 32408
rect 187601 32464 190164 32466
rect 187601 32408 187606 32464
rect 187662 32408 190164 32464
rect 187601 32406 190164 32408
rect 216581 32464 219052 32466
rect 216581 32408 216586 32464
rect 216642 32408 219052 32464
rect 216581 32406 219052 32408
rect 246941 32464 248124 32466
rect 246941 32408 246946 32464
rect 247002 32408 248124 32464
rect 246941 32406 248124 32408
rect 275921 32464 277196 32466
rect 275921 32408 275926 32464
rect 275982 32408 277196 32464
rect 275921 32406 277196 32408
rect 304901 32464 306084 32466
rect 304901 32408 304906 32464
rect 304962 32408 306084 32464
rect 304901 32406 306084 32408
rect 333881 32464 335156 32466
rect 333881 32408 333886 32464
rect 333942 32408 335156 32464
rect 333881 32406 335156 32408
rect 362861 32464 364044 32466
rect 362861 32408 362866 32464
rect 362922 32408 364044 32464
rect 362861 32406 364044 32408
rect 391841 32464 393116 32466
rect 391841 32408 391846 32464
rect 391902 32408 393116 32464
rect 391841 32406 393116 32408
rect 420821 32464 422188 32466
rect 420821 32408 420826 32464
rect 420882 32408 422188 32464
rect 420821 32406 422188 32408
rect 449801 32464 451076 32466
rect 449801 32408 449806 32464
rect 449862 32408 451076 32464
rect 449801 32406 451076 32408
rect 478781 32464 480148 32466
rect 478781 32408 478786 32464
rect 478842 32408 480148 32464
rect 509006 32436 509066 32950
rect 536649 32466 536715 32469
rect 536649 32464 538108 32466
rect 478781 32406 480148 32408
rect 536649 32408 536654 32464
rect 536710 32408 538108 32464
rect 536649 32406 538108 32408
rect 71405 32403 71471 32406
rect 100385 32403 100451 32406
rect 129641 32403 129707 32406
rect 158621 32403 158687 32406
rect 187601 32403 187667 32406
rect 216581 32403 216647 32406
rect 246941 32403 247007 32406
rect 275921 32403 275987 32406
rect 304901 32403 304967 32406
rect 333881 32403 333947 32406
rect 362861 32403 362927 32406
rect 391841 32403 391907 32406
rect 420821 32403 420887 32406
rect 449801 32403 449867 32406
rect 478781 32403 478847 32406
rect 536649 32403 536715 32406
rect 79918 31862 81266 31922
rect 79918 31756 79978 31862
rect 81206 31756 81266 31862
rect 456934 31862 458282 31922
rect 108836 31726 110308 31786
rect 137908 31726 139380 31786
rect 166796 31726 168268 31786
rect 195868 31726 197340 31786
rect 224940 31726 226412 31786
rect 253828 31726 255300 31786
rect 282900 31726 284372 31786
rect 311788 31726 313260 31786
rect 340860 31726 342332 31786
rect 369932 31726 371404 31786
rect 398820 31726 400292 31786
rect 427892 31726 429364 31786
rect 456934 31756 456994 31862
rect 458222 31756 458282 31862
rect 485852 31726 487324 31786
rect 514924 31726 516396 31786
rect 543812 31726 545284 31786
rect 64229 31650 64295 31653
rect 61916 31648 64295 31650
rect 61916 31592 64234 31648
rect 64290 31592 64295 31648
rect 61916 31590 64295 31592
rect 64229 31587 64295 31590
rect 12433 31106 12499 31109
rect 12433 31104 16100 31106
rect 12433 31048 12438 31104
rect 12494 31048 16100 31104
rect 12433 31046 16100 31048
rect 12433 31043 12499 31046
rect 64229 30290 64295 30293
rect 61916 30288 64295 30290
rect 61916 30232 64234 30288
rect 64290 30232 64295 30288
rect 61916 30230 64295 30232
rect 64229 30227 64295 30230
rect 79918 30154 79978 30260
rect 81206 30154 81266 30260
rect 108836 30230 110308 30290
rect 137908 30230 139380 30290
rect 166796 30230 168268 30290
rect 195868 30230 197340 30290
rect 224940 30230 226412 30290
rect 253828 30230 255300 30290
rect 282900 30230 284372 30290
rect 311788 30230 313260 30290
rect 340860 30230 342332 30290
rect 369932 30230 371404 30290
rect 398820 30230 400292 30290
rect 427892 30230 429364 30290
rect 79918 30094 81266 30154
rect 456934 30154 456994 30260
rect 458222 30154 458282 30260
rect 485852 30230 487324 30290
rect 514924 30230 516396 30290
rect 543812 30230 545284 30290
rect 456934 30094 458282 30154
rect 507577 30018 507643 30021
rect 507577 30016 509066 30018
rect 507577 29960 507582 30016
rect 507638 29960 509066 30016
rect 507577 29958 509066 29960
rect 507577 29955 507643 29958
rect 13629 29746 13695 29749
rect 13629 29744 16100 29746
rect 13629 29688 13634 29744
rect 13690 29688 16100 29744
rect 13629 29686 16100 29688
rect 13629 29683 13695 29686
rect 71497 29474 71563 29477
rect 100477 29474 100543 29477
rect 129457 29474 129523 29477
rect 158437 29474 158503 29477
rect 187417 29474 187483 29477
rect 216397 29474 216463 29477
rect 246757 29474 246823 29477
rect 275737 29474 275803 29477
rect 304717 29474 304783 29477
rect 333697 29474 333763 29477
rect 362677 29474 362743 29477
rect 391657 29474 391723 29477
rect 420637 29474 420703 29477
rect 449617 29474 449683 29477
rect 478597 29474 478663 29477
rect 71497 29472 74060 29474
rect 71497 29416 71502 29472
rect 71558 29416 74060 29472
rect 71497 29414 74060 29416
rect 100477 29472 103132 29474
rect 100477 29416 100482 29472
rect 100538 29416 103132 29472
rect 100477 29414 103132 29416
rect 129457 29472 132204 29474
rect 129457 29416 129462 29472
rect 129518 29416 132204 29472
rect 129457 29414 132204 29416
rect 158437 29472 161092 29474
rect 158437 29416 158442 29472
rect 158498 29416 161092 29472
rect 158437 29414 161092 29416
rect 187417 29472 190164 29474
rect 187417 29416 187422 29472
rect 187478 29416 190164 29472
rect 187417 29414 190164 29416
rect 216397 29472 219052 29474
rect 216397 29416 216402 29472
rect 216458 29416 219052 29472
rect 216397 29414 219052 29416
rect 246757 29472 248124 29474
rect 246757 29416 246762 29472
rect 246818 29416 248124 29472
rect 246757 29414 248124 29416
rect 275737 29472 277196 29474
rect 275737 29416 275742 29472
rect 275798 29416 277196 29472
rect 275737 29414 277196 29416
rect 304717 29472 306084 29474
rect 304717 29416 304722 29472
rect 304778 29416 306084 29472
rect 304717 29414 306084 29416
rect 333697 29472 335156 29474
rect 333697 29416 333702 29472
rect 333758 29416 335156 29472
rect 333697 29414 335156 29416
rect 362677 29472 364044 29474
rect 362677 29416 362682 29472
rect 362738 29416 364044 29472
rect 362677 29414 364044 29416
rect 391657 29472 393116 29474
rect 391657 29416 391662 29472
rect 391718 29416 393116 29472
rect 391657 29414 393116 29416
rect 420637 29472 422188 29474
rect 420637 29416 420642 29472
rect 420698 29416 422188 29472
rect 420637 29414 422188 29416
rect 449617 29472 451076 29474
rect 449617 29416 449622 29472
rect 449678 29416 451076 29472
rect 449617 29414 451076 29416
rect 478597 29472 480148 29474
rect 478597 29416 478602 29472
rect 478658 29416 480148 29472
rect 509006 29444 509066 29958
rect 536741 29474 536807 29477
rect 536741 29472 538108 29474
rect 478597 29414 480148 29416
rect 536741 29416 536746 29472
rect 536802 29416 538108 29472
rect 536741 29414 538108 29416
rect 71497 29411 71563 29414
rect 100477 29411 100543 29414
rect 129457 29411 129523 29414
rect 158437 29411 158503 29414
rect 187417 29411 187483 29414
rect 216397 29411 216463 29414
rect 246757 29411 246823 29414
rect 275737 29411 275803 29414
rect 304717 29411 304783 29414
rect 333697 29411 333763 29414
rect 362677 29411 362743 29414
rect 391657 29411 391723 29414
rect 420637 29411 420703 29414
rect 449617 29411 449683 29414
rect 478597 29411 478663 29414
rect 536741 29411 536807 29414
rect 79918 28870 81266 28930
rect 79918 28764 79978 28870
rect 81206 28764 81266 28870
rect 456934 28870 458282 28930
rect 108836 28734 110308 28794
rect 137908 28734 139380 28794
rect 166796 28734 168268 28794
rect 195868 28734 197340 28794
rect 224940 28734 226412 28794
rect 253828 28734 255300 28794
rect 282900 28734 284372 28794
rect 311788 28734 313260 28794
rect 340860 28734 342332 28794
rect 369932 28734 371404 28794
rect 398820 28734 400292 28794
rect 427892 28734 429364 28794
rect 456934 28764 456994 28870
rect 458222 28764 458282 28870
rect 485852 28734 487324 28794
rect 514924 28734 516396 28794
rect 543812 28734 545284 28794
rect 64321 28386 64387 28389
rect 61916 28384 64387 28386
rect 61916 28328 64326 28384
rect 64382 28328 64387 28384
rect 61916 28326 64387 28328
rect 64321 28323 64387 28326
rect 13537 27706 13603 27709
rect 13537 27704 16100 27706
rect 13537 27648 13542 27704
rect 13598 27648 16100 27704
rect 13537 27646 16100 27648
rect 13537 27643 13603 27646
rect 79918 27374 81266 27434
rect 79918 27268 79978 27374
rect 81206 27268 81266 27374
rect 456934 27374 458282 27434
rect 108836 27238 110308 27298
rect 137908 27238 139380 27298
rect 166796 27238 168268 27298
rect 195868 27238 197340 27298
rect 224940 27238 226412 27298
rect 253828 27238 255300 27298
rect 282900 27238 284372 27298
rect 311788 27238 313260 27298
rect 340860 27238 342332 27298
rect 369932 27238 371404 27298
rect 398820 27238 400292 27298
rect 427892 27238 429364 27298
rect 456934 27268 456994 27374
rect 458222 27268 458282 27374
rect 485852 27238 487324 27298
rect 514924 27238 516396 27298
rect 543812 27238 545284 27298
rect 63493 27026 63559 27029
rect 61916 27024 63559 27026
rect 61916 26968 63498 27024
rect 63554 26968 63559 27024
rect 61916 26966 63559 26968
rect 63493 26963 63559 26966
rect 507209 27026 507275 27029
rect 507209 27024 509066 27026
rect 507209 26968 507214 27024
rect 507270 26968 509066 27024
rect 507209 26966 509066 26968
rect 507209 26963 507275 26966
rect 71037 26482 71103 26485
rect 100109 26482 100175 26485
rect 129089 26482 129155 26485
rect 158069 26482 158135 26485
rect 187049 26482 187115 26485
rect 216029 26482 216095 26485
rect 246389 26482 246455 26485
rect 275369 26482 275435 26485
rect 304349 26482 304415 26485
rect 333329 26482 333395 26485
rect 362309 26482 362375 26485
rect 391289 26482 391355 26485
rect 420269 26482 420335 26485
rect 449249 26482 449315 26485
rect 478229 26482 478295 26485
rect 71037 26480 74060 26482
rect 71037 26424 71042 26480
rect 71098 26424 74060 26480
rect 71037 26422 74060 26424
rect 100109 26480 103132 26482
rect 100109 26424 100114 26480
rect 100170 26424 103132 26480
rect 100109 26422 103132 26424
rect 129089 26480 132204 26482
rect 129089 26424 129094 26480
rect 129150 26424 132204 26480
rect 129089 26422 132204 26424
rect 158069 26480 161092 26482
rect 158069 26424 158074 26480
rect 158130 26424 161092 26480
rect 158069 26422 161092 26424
rect 187049 26480 190164 26482
rect 187049 26424 187054 26480
rect 187110 26424 190164 26480
rect 187049 26422 190164 26424
rect 216029 26480 219052 26482
rect 216029 26424 216034 26480
rect 216090 26424 219052 26480
rect 216029 26422 219052 26424
rect 246389 26480 248124 26482
rect 246389 26424 246394 26480
rect 246450 26424 248124 26480
rect 246389 26422 248124 26424
rect 275369 26480 277196 26482
rect 275369 26424 275374 26480
rect 275430 26424 277196 26480
rect 275369 26422 277196 26424
rect 304349 26480 306084 26482
rect 304349 26424 304354 26480
rect 304410 26424 306084 26480
rect 304349 26422 306084 26424
rect 333329 26480 335156 26482
rect 333329 26424 333334 26480
rect 333390 26424 335156 26480
rect 333329 26422 335156 26424
rect 362309 26480 364044 26482
rect 362309 26424 362314 26480
rect 362370 26424 364044 26480
rect 362309 26422 364044 26424
rect 391289 26480 393116 26482
rect 391289 26424 391294 26480
rect 391350 26424 393116 26480
rect 391289 26422 393116 26424
rect 420269 26480 422188 26482
rect 420269 26424 420274 26480
rect 420330 26424 422188 26480
rect 420269 26422 422188 26424
rect 449249 26480 451076 26482
rect 449249 26424 449254 26480
rect 449310 26424 451076 26480
rect 449249 26422 451076 26424
rect 478229 26480 480148 26482
rect 478229 26424 478234 26480
rect 478290 26424 480148 26480
rect 509006 26452 509066 26966
rect 536189 26482 536255 26485
rect 536189 26480 538108 26482
rect 478229 26422 480148 26424
rect 536189 26424 536194 26480
rect 536250 26424 538108 26480
rect 536189 26422 538108 26424
rect 71037 26419 71103 26422
rect 100109 26419 100175 26422
rect 129089 26419 129155 26422
rect 158069 26419 158135 26422
rect 187049 26419 187115 26422
rect 216029 26419 216095 26422
rect 246389 26419 246455 26422
rect 275369 26419 275435 26422
rect 304349 26419 304415 26422
rect 333329 26419 333395 26422
rect 362309 26419 362375 26422
rect 391289 26419 391355 26422
rect 420269 26419 420335 26422
rect 449249 26419 449315 26422
rect 478229 26419 478295 26422
rect 536189 26419 536255 26422
rect 13629 26346 13695 26349
rect 13629 26344 16100 26346
rect 13629 26288 13634 26344
rect 13690 26288 16100 26344
rect 13629 26286 16100 26288
rect 13629 26283 13695 26286
rect 79918 25878 81266 25938
rect 79918 25772 79978 25878
rect 81206 25772 81266 25878
rect 456934 25878 458282 25938
rect 108836 25742 110308 25802
rect 137908 25742 139380 25802
rect 166796 25742 168268 25802
rect 195868 25742 197340 25802
rect 224940 25742 226412 25802
rect 253828 25742 255300 25802
rect 282900 25742 284372 25802
rect 311788 25742 313260 25802
rect 340860 25742 342332 25802
rect 369932 25742 371404 25802
rect 398820 25742 400292 25802
rect 427892 25742 429364 25802
rect 456934 25772 456994 25878
rect 458222 25772 458282 25878
rect 485852 25742 487324 25802
rect 514924 25742 516396 25802
rect 543812 25742 545284 25802
rect 64321 24986 64387 24989
rect 61916 24984 64387 24986
rect 61916 24928 64326 24984
rect 64382 24928 64387 24984
rect 61916 24926 64387 24928
rect 64321 24923 64387 24926
rect 79918 24382 81266 24442
rect 79918 24276 79978 24382
rect 81206 24276 81266 24382
rect 456934 24382 458282 24442
rect 108836 24246 110308 24306
rect 137908 24246 139380 24306
rect 166796 24246 168268 24306
rect 195868 24246 197340 24306
rect 224940 24246 226412 24306
rect 253828 24246 255300 24306
rect 282900 24246 284372 24306
rect 311788 24246 313260 24306
rect 340860 24246 342332 24306
rect 369932 24246 371404 24306
rect 398820 24246 400292 24306
rect 427892 24246 429364 24306
rect 456934 24276 456994 24382
rect 458222 24276 458282 24382
rect 485852 24246 487324 24306
rect 514924 24246 516396 24306
rect 543812 24246 545284 24306
rect 13721 24170 13787 24173
rect 13721 24168 16100 24170
rect 13721 24112 13726 24168
rect 13782 24112 16100 24168
rect 13721 24110 16100 24112
rect 13721 24107 13787 24110
rect 507117 24034 507183 24037
rect 507117 24032 509066 24034
rect 507117 23976 507122 24032
rect 507178 23976 509066 24032
rect 507117 23974 509066 23976
rect 507117 23971 507183 23974
rect 64137 23626 64203 23629
rect 61916 23624 64203 23626
rect 61916 23568 64142 23624
rect 64198 23568 64203 23624
rect 61916 23566 64203 23568
rect 64137 23563 64203 23566
rect 71129 23490 71195 23493
rect 100017 23490 100083 23493
rect 128997 23490 129063 23493
rect 157977 23490 158043 23493
rect 186957 23490 187023 23493
rect 215937 23490 216003 23493
rect 246297 23490 246363 23493
rect 275277 23490 275343 23493
rect 304257 23490 304323 23493
rect 333237 23490 333303 23493
rect 362217 23490 362283 23493
rect 391197 23490 391263 23493
rect 420177 23490 420243 23493
rect 449157 23490 449223 23493
rect 478137 23490 478203 23493
rect 71129 23488 74060 23490
rect 71129 23432 71134 23488
rect 71190 23432 74060 23488
rect 71129 23430 74060 23432
rect 100017 23488 103132 23490
rect 100017 23432 100022 23488
rect 100078 23432 103132 23488
rect 100017 23430 103132 23432
rect 128997 23488 132204 23490
rect 128997 23432 129002 23488
rect 129058 23432 132204 23488
rect 128997 23430 132204 23432
rect 157977 23488 161092 23490
rect 157977 23432 157982 23488
rect 158038 23432 161092 23488
rect 157977 23430 161092 23432
rect 186957 23488 190164 23490
rect 186957 23432 186962 23488
rect 187018 23432 190164 23488
rect 186957 23430 190164 23432
rect 215937 23488 219052 23490
rect 215937 23432 215942 23488
rect 215998 23432 219052 23488
rect 215937 23430 219052 23432
rect 246297 23488 248124 23490
rect 246297 23432 246302 23488
rect 246358 23432 248124 23488
rect 246297 23430 248124 23432
rect 275277 23488 277196 23490
rect 275277 23432 275282 23488
rect 275338 23432 277196 23488
rect 275277 23430 277196 23432
rect 304257 23488 306084 23490
rect 304257 23432 304262 23488
rect 304318 23432 306084 23488
rect 304257 23430 306084 23432
rect 333237 23488 335156 23490
rect 333237 23432 333242 23488
rect 333298 23432 335156 23488
rect 333237 23430 335156 23432
rect 362217 23488 364044 23490
rect 362217 23432 362222 23488
rect 362278 23432 364044 23488
rect 362217 23430 364044 23432
rect 391197 23488 393116 23490
rect 391197 23432 391202 23488
rect 391258 23432 393116 23488
rect 391197 23430 393116 23432
rect 420177 23488 422188 23490
rect 420177 23432 420182 23488
rect 420238 23432 422188 23488
rect 420177 23430 422188 23432
rect 449157 23488 451076 23490
rect 449157 23432 449162 23488
rect 449218 23432 451076 23488
rect 449157 23430 451076 23432
rect 478137 23488 480148 23490
rect 478137 23432 478142 23488
rect 478198 23432 480148 23488
rect 509006 23460 509066 23974
rect 536097 23490 536163 23493
rect 536097 23488 538108 23490
rect 478137 23430 480148 23432
rect 536097 23432 536102 23488
rect 536158 23432 538108 23488
rect 536097 23430 538108 23432
rect 71129 23427 71195 23430
rect 100017 23427 100083 23430
rect 128997 23427 129063 23430
rect 157977 23427 158043 23430
rect 186957 23427 187023 23430
rect 215937 23427 216003 23430
rect 246297 23427 246363 23430
rect 275277 23427 275343 23430
rect 304257 23427 304323 23430
rect 333237 23427 333303 23430
rect 362217 23427 362283 23430
rect 391197 23427 391263 23430
rect 420177 23427 420243 23430
rect 449157 23427 449223 23430
rect 478137 23427 478203 23430
rect 536097 23427 536163 23430
rect 12433 22946 12499 22949
rect 12433 22944 16100 22946
rect 12433 22888 12438 22944
rect 12494 22888 16100 22944
rect 12433 22886 16100 22888
rect 79918 22886 81266 22946
rect 12433 22883 12499 22886
rect 79918 22780 79978 22886
rect 81206 22780 81266 22886
rect 456934 22886 458282 22946
rect 108836 22750 110308 22810
rect 137908 22750 139380 22810
rect 166796 22750 168268 22810
rect 195868 22750 197340 22810
rect 224940 22750 226412 22810
rect 253828 22750 255300 22810
rect 282900 22750 284372 22810
rect 311788 22750 313260 22810
rect 340860 22750 342332 22810
rect 369932 22750 371404 22810
rect 398820 22750 400292 22810
rect 427892 22750 429364 22810
rect 456934 22780 456994 22886
rect 458222 22780 458282 22886
rect 485852 22750 487324 22810
rect 514924 22750 516396 22810
rect 543812 22750 545284 22810
rect 63493 21450 63559 21453
rect 61916 21448 63559 21450
rect 61916 21392 63498 21448
rect 63554 21392 63559 21448
rect 61916 21390 63559 21392
rect 63493 21387 63559 21390
rect 79918 21390 81266 21450
rect 79918 21284 79978 21390
rect 81206 21284 81266 21390
rect 456934 21390 458282 21450
rect 108836 21254 110308 21314
rect 137908 21254 139380 21314
rect 166796 21254 168268 21314
rect 195868 21254 197340 21314
rect 224940 21254 226412 21314
rect 253828 21254 255300 21314
rect 282900 21254 284372 21314
rect 311788 21254 313260 21314
rect 340860 21254 342332 21314
rect 369932 21254 371404 21314
rect 398820 21254 400292 21314
rect 427892 21254 429364 21314
rect 456934 21284 456994 21390
rect 458222 21284 458282 21390
rect 485852 21254 487324 21314
rect 514924 21254 516396 21314
rect 543812 21254 545284 21314
rect 12433 20906 12499 20909
rect 12433 20904 16100 20906
rect 12433 20848 12438 20904
rect 12494 20848 16100 20904
rect 12433 20846 16100 20848
rect 12433 20843 12499 20846
rect 61285 20634 61351 20637
rect 61285 20632 61394 20634
rect 61285 20576 61290 20632
rect 61346 20576 61394 20632
rect 61285 20571 61394 20576
rect 61334 20196 61394 20571
rect 70393 20498 70459 20501
rect 100017 20498 100083 20501
rect 128997 20498 129063 20501
rect 157977 20498 158043 20501
rect 186957 20498 187023 20501
rect 215937 20498 216003 20501
rect 246297 20498 246363 20501
rect 275277 20498 275343 20501
rect 304257 20498 304323 20501
rect 333237 20498 333303 20501
rect 362217 20498 362283 20501
rect 391197 20498 391263 20501
rect 420177 20498 420243 20501
rect 449157 20498 449223 20501
rect 478137 20498 478203 20501
rect 536097 20498 536163 20501
rect 70393 20496 74060 20498
rect 70393 20440 70398 20496
rect 70454 20440 74060 20496
rect 70393 20438 74060 20440
rect 100017 20496 103132 20498
rect 100017 20440 100022 20496
rect 100078 20440 103132 20496
rect 100017 20438 103132 20440
rect 128997 20496 132204 20498
rect 128997 20440 129002 20496
rect 129058 20440 132204 20496
rect 128997 20438 132204 20440
rect 157977 20496 161092 20498
rect 157977 20440 157982 20496
rect 158038 20440 161092 20496
rect 157977 20438 161092 20440
rect 186957 20496 190164 20498
rect 186957 20440 186962 20496
rect 187018 20440 190164 20496
rect 186957 20438 190164 20440
rect 215937 20496 219052 20498
rect 215937 20440 215942 20496
rect 215998 20440 219052 20496
rect 215937 20438 219052 20440
rect 246297 20496 248124 20498
rect 246297 20440 246302 20496
rect 246358 20440 248124 20496
rect 246297 20438 248124 20440
rect 275277 20496 277196 20498
rect 275277 20440 275282 20496
rect 275338 20440 277196 20496
rect 275277 20438 277196 20440
rect 304257 20496 306084 20498
rect 304257 20440 304262 20496
rect 304318 20440 306084 20496
rect 304257 20438 306084 20440
rect 333237 20496 335156 20498
rect 333237 20440 333242 20496
rect 333298 20440 335156 20496
rect 333237 20438 335156 20440
rect 362217 20496 364044 20498
rect 362217 20440 362222 20496
rect 362278 20440 364044 20496
rect 362217 20438 364044 20440
rect 391197 20496 393116 20498
rect 391197 20440 391202 20496
rect 391258 20440 393116 20496
rect 391197 20438 393116 20440
rect 420177 20496 422188 20498
rect 420177 20440 420182 20496
rect 420238 20440 422188 20496
rect 420177 20438 422188 20440
rect 449157 20496 451076 20498
rect 449157 20440 449162 20496
rect 449218 20440 451076 20496
rect 449157 20438 451076 20440
rect 478137 20496 480148 20498
rect 478137 20440 478142 20496
rect 478198 20440 480148 20496
rect 536097 20496 538108 20498
rect 478137 20438 480148 20440
rect 70393 20435 70459 20438
rect 100017 20435 100083 20438
rect 128997 20435 129063 20438
rect 157977 20435 158043 20438
rect 186957 20435 187023 20438
rect 215937 20435 216003 20438
rect 246297 20435 246363 20438
rect 275277 20435 275343 20438
rect 304257 20435 304323 20438
rect 333237 20435 333303 20438
rect 362217 20435 362283 20438
rect 391197 20435 391263 20438
rect 420177 20435 420243 20438
rect 449157 20435 449223 20438
rect 478137 20435 478203 20438
rect 507117 19954 507183 19957
rect 509006 19954 509066 20468
rect 536097 20440 536102 20496
rect 536158 20440 538108 20496
rect 536097 20438 538108 20440
rect 536097 20435 536163 20438
rect 79918 19894 81266 19954
rect 79918 19788 79978 19894
rect 81206 19788 81266 19894
rect 456934 19894 458282 19954
rect 108836 19758 110308 19818
rect 137908 19758 139380 19818
rect 166796 19758 168268 19818
rect 195868 19758 197340 19818
rect 224940 19758 226412 19818
rect 253828 19758 255300 19818
rect 282900 19758 284372 19818
rect 311788 19758 313260 19818
rect 340860 19758 342332 19818
rect 369932 19758 371404 19818
rect 398820 19758 400292 19818
rect 427892 19758 429364 19818
rect 456934 19788 456994 19894
rect 458222 19788 458282 19894
rect 507117 19952 509066 19954
rect 507117 19896 507122 19952
rect 507178 19896 509066 19952
rect 507117 19894 509066 19896
rect 507117 19891 507183 19894
rect 485852 19758 487324 19818
rect 514924 19758 516396 19818
rect 543812 19758 545284 19818
rect 583520 19668 584960 19908
rect 11789 19546 11855 19549
rect 11789 19544 16100 19546
rect -960 19410 480 19500
rect 11789 19488 11794 19544
rect 11850 19488 16100 19544
rect 11789 19486 16100 19488
rect 11789 19483 11855 19486
rect 3693 19410 3759 19413
rect -960 19408 3759 19410
rect -960 19352 3698 19408
rect 3754 19352 3759 19408
rect -960 19350 3759 19352
rect -960 19260 480 19350
rect 3693 19347 3759 19350
rect 79918 18398 81266 18458
rect 79918 18292 79978 18398
rect 81206 18292 81266 18398
rect 456934 18398 458282 18458
rect 108836 18262 110308 18322
rect 137908 18262 139380 18322
rect 166796 18262 168268 18322
rect 195868 18262 197340 18322
rect 224940 18262 226412 18322
rect 253828 18262 255300 18322
rect 282900 18262 284372 18322
rect 311788 18262 313260 18322
rect 340860 18262 342332 18322
rect 369932 18262 371404 18322
rect 398820 18262 400292 18322
rect 427892 18262 429364 18322
rect 456934 18292 456994 18398
rect 458222 18292 458282 18398
rect 485852 18262 487324 18322
rect 514924 18262 516396 18322
rect 543812 18262 545284 18322
rect 64413 18186 64479 18189
rect 61916 18184 64479 18186
rect 61916 18128 64418 18184
rect 64474 18128 64479 18184
rect 61916 18126 64479 18128
rect 64413 18123 64479 18126
rect 12433 17506 12499 17509
rect 70393 17506 70459 17509
rect 99833 17506 99899 17509
rect 128813 17506 128879 17509
rect 157517 17506 157583 17509
rect 186773 17506 186839 17509
rect 215753 17506 215819 17509
rect 245653 17506 245719 17509
rect 274633 17506 274699 17509
rect 303613 17506 303679 17509
rect 332593 17506 332659 17509
rect 361573 17506 361639 17509
rect 390553 17506 390619 17509
rect 419533 17506 419599 17509
rect 448513 17506 448579 17509
rect 477493 17506 477559 17509
rect 535453 17506 535519 17509
rect 12433 17504 16100 17506
rect 12433 17448 12438 17504
rect 12494 17448 16100 17504
rect 12433 17446 16100 17448
rect 70393 17504 74060 17506
rect 70393 17448 70398 17504
rect 70454 17448 74060 17504
rect 70393 17446 74060 17448
rect 99833 17504 103132 17506
rect 99833 17448 99838 17504
rect 99894 17448 103132 17504
rect 99833 17446 103132 17448
rect 128813 17504 132204 17506
rect 128813 17448 128818 17504
rect 128874 17448 132204 17504
rect 128813 17446 132204 17448
rect 157517 17504 161092 17506
rect 157517 17448 157522 17504
rect 157578 17448 161092 17504
rect 157517 17446 161092 17448
rect 186773 17504 190164 17506
rect 186773 17448 186778 17504
rect 186834 17448 190164 17504
rect 186773 17446 190164 17448
rect 215753 17504 219052 17506
rect 215753 17448 215758 17504
rect 215814 17448 219052 17504
rect 215753 17446 219052 17448
rect 245653 17504 248124 17506
rect 245653 17448 245658 17504
rect 245714 17448 248124 17504
rect 245653 17446 248124 17448
rect 274633 17504 277196 17506
rect 274633 17448 274638 17504
rect 274694 17448 277196 17504
rect 274633 17446 277196 17448
rect 303613 17504 306084 17506
rect 303613 17448 303618 17504
rect 303674 17448 306084 17504
rect 303613 17446 306084 17448
rect 332593 17504 335156 17506
rect 332593 17448 332598 17504
rect 332654 17448 335156 17504
rect 332593 17446 335156 17448
rect 361573 17504 364044 17506
rect 361573 17448 361578 17504
rect 361634 17448 364044 17504
rect 361573 17446 364044 17448
rect 390553 17504 393116 17506
rect 390553 17448 390558 17504
rect 390614 17448 393116 17504
rect 390553 17446 393116 17448
rect 419533 17504 422188 17506
rect 419533 17448 419538 17504
rect 419594 17448 422188 17504
rect 419533 17446 422188 17448
rect 448513 17504 451076 17506
rect 448513 17448 448518 17504
rect 448574 17448 451076 17504
rect 448513 17446 451076 17448
rect 477493 17504 480148 17506
rect 477493 17448 477498 17504
rect 477554 17448 480148 17504
rect 535453 17504 538108 17506
rect 477493 17446 480148 17448
rect 12433 17443 12499 17446
rect 70393 17443 70459 17446
rect 99833 17443 99899 17446
rect 128813 17443 128879 17446
rect 157517 17443 157583 17446
rect 186773 17443 186839 17446
rect 215753 17443 215819 17446
rect 245653 17443 245719 17446
rect 274633 17443 274699 17446
rect 303613 17443 303679 17446
rect 332593 17443 332659 17446
rect 361573 17443 361639 17446
rect 390553 17443 390619 17446
rect 419533 17443 419599 17446
rect 448513 17443 448579 17446
rect 477493 17443 477559 17446
rect 506473 17098 506539 17101
rect 509006 17098 509066 17476
rect 535453 17448 535458 17504
rect 535514 17448 538108 17504
rect 535453 17446 538108 17448
rect 535453 17443 535519 17446
rect 506473 17096 509066 17098
rect 506473 17040 506478 17096
rect 506534 17040 509066 17096
rect 506473 17038 509066 17040
rect 506473 17035 506539 17038
rect 79918 16902 81266 16962
rect 64597 16826 64663 16829
rect 61916 16824 64663 16826
rect 61916 16768 64602 16824
rect 64658 16768 64663 16824
rect 79918 16796 79978 16902
rect 81206 16796 81266 16902
rect 456934 16902 458282 16962
rect 61916 16766 64663 16768
rect 108836 16766 110308 16826
rect 137908 16766 139380 16826
rect 166796 16766 168268 16826
rect 195868 16766 197340 16826
rect 224940 16766 226412 16826
rect 253828 16766 255300 16826
rect 282900 16766 284372 16826
rect 311788 16766 313260 16826
rect 340860 16766 342332 16826
rect 369932 16766 371404 16826
rect 398820 16766 400292 16826
rect 427892 16766 429364 16826
rect 456934 16796 456994 16902
rect 458222 16796 458282 16902
rect 485852 16766 487324 16826
rect 514924 16766 516396 16826
rect 543812 16766 545284 16826
rect 64597 16763 64663 16766
rect 45502 16492 45508 16556
rect 45572 16554 45578 16556
rect 46013 16554 46079 16557
rect 45572 16552 46079 16554
rect 45572 16496 46018 16552
rect 46074 16496 46079 16552
rect 45572 16494 46079 16496
rect 45572 16492 45578 16494
rect 46013 16491 46079 16494
rect 54334 16492 54340 16556
rect 54404 16554 54410 16556
rect 57605 16554 57671 16557
rect 54404 16552 57671 16554
rect 54404 16496 57610 16552
rect 57666 16496 57671 16552
rect 54404 16494 57671 16496
rect 54404 16492 54410 16494
rect 57605 16491 57671 16494
rect 3550 13500 3556 13564
rect 3620 13562 3626 13564
rect 35341 13562 35407 13565
rect 3620 13560 35407 13562
rect 3620 13504 35346 13560
rect 35402 13504 35407 13560
rect 3620 13502 35407 13504
rect 3620 13500 3626 13502
rect 35341 13499 35407 13502
rect 52729 13562 52795 13565
rect 558862 13562 558868 13564
rect 52729 13560 558868 13562
rect 52729 13504 52734 13560
rect 52790 13504 558868 13560
rect 52729 13502 558868 13504
rect 52729 13499 52795 13502
rect 558862 13500 558868 13502
rect 558932 13500 558938 13564
rect 41781 13426 41847 13429
rect 429326 13426 429332 13428
rect 41781 13424 429332 13426
rect 41781 13368 41786 13424
rect 41842 13368 429332 13424
rect 41781 13366 429332 13368
rect 41781 13363 41847 13366
rect 429326 13364 429332 13366
rect 429396 13364 429402 13428
rect 26969 13290 27035 13293
rect 397678 13290 397684 13292
rect 26969 13288 397684 13290
rect 26969 13232 26974 13288
rect 27030 13232 397684 13288
rect 26969 13230 397684 13232
rect 26969 13227 27035 13230
rect 397678 13228 397684 13230
rect 397748 13228 397754 13292
rect 48221 13154 48287 13157
rect 169702 13154 169708 13156
rect 48221 13152 169708 13154
rect 48221 13096 48226 13152
rect 48282 13096 169708 13152
rect 48221 13094 169708 13096
rect 48221 13091 48287 13094
rect 169702 13092 169708 13094
rect 169772 13092 169778 13156
rect 19241 13018 19307 13021
rect 527398 13018 527404 13020
rect 19241 13016 527404 13018
rect 19241 12960 19246 13016
rect 19302 12960 527404 13016
rect 19241 12958 527404 12960
rect 19241 12955 19307 12958
rect 527398 12956 527404 12958
rect 527468 12956 527474 13020
rect -960 6490 480 6580
rect -960 6430 674 6490
rect 583520 6476 584960 6716
rect -960 6354 480 6430
rect 614 6354 674 6430
rect -960 6340 674 6354
rect 246 6294 674 6340
rect 246 5810 306 6294
rect 246 5750 6930 5810
rect 6870 5674 6930 5750
rect 42742 5674 42748 5676
rect 6870 5614 42748 5674
rect 42742 5612 42748 5614
rect 42812 5612 42818 5676
rect 50838 3436 50844 3500
rect 50908 3498 50914 3500
rect 132953 3498 133019 3501
rect 50908 3496 133019 3498
rect 50908 3440 132958 3496
rect 133014 3440 133019 3496
rect 50908 3438 133019 3440
rect 50908 3436 50914 3438
rect 132953 3435 133019 3438
rect 39798 3300 39804 3364
rect 39868 3362 39874 3364
rect 136449 3362 136515 3365
rect 39868 3360 136515 3362
rect 39868 3304 136454 3360
rect 136510 3304 136515 3360
rect 39868 3302 136515 3304
rect 39868 3300 39874 3302
rect 136449 3299 136515 3302
<< via3 >>
rect 169708 699756 169772 699820
rect 397684 699756 397748 699820
rect 429332 699756 429396 699820
rect 527404 699756 527468 699820
rect 558868 699756 558932 699820
rect 3372 684252 3436 684316
rect 3556 606052 3620 606116
rect 45324 500924 45388 500988
rect 54340 474812 54404 474876
rect 249012 65588 249076 65652
rect 277900 65588 277964 65652
rect 306972 65588 307036 65652
rect 335860 65588 335924 65652
rect 364932 65588 364996 65652
rect 393820 65588 393884 65652
rect 422892 65588 422956 65652
rect 249012 43284 249076 43348
rect 277900 43556 277964 43620
rect 306972 43556 307036 43620
rect 335860 43556 335924 43620
rect 364932 43556 364996 43620
rect 393820 43556 393884 43620
rect 422892 43556 422956 43620
rect 3372 37844 3436 37908
rect 39804 35260 39868 35324
rect 42748 35260 42812 35324
rect 50844 35260 50908 35324
rect 45508 16492 45572 16556
rect 54340 16492 54404 16556
rect 3556 13500 3620 13564
rect 558868 13500 558932 13564
rect 429332 13364 429396 13428
rect 397684 13228 397748 13292
rect 169708 13092 169772 13156
rect 527404 12956 527468 13020
rect 42748 5612 42812 5676
rect 50844 3436 50908 3500
rect 39804 3300 39868 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 -7066 -8106 711002
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 -6106 -7146 710042
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 -5146 -6186 709082
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 -4186 -5226 708122
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 -3226 -4266 707162
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 -2266 -3306 706202
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 698454 -2346 705242
rect 37994 705798 38614 711590
rect 37994 705562 38026 705798
rect 38262 705562 38346 705798
rect 38582 705562 38614 705798
rect 37994 705478 38614 705562
rect 37994 705242 38026 705478
rect 38262 705242 38346 705478
rect 38582 705242 38614 705478
rect -2966 698218 -2934 698454
rect -2698 698218 -2614 698454
rect -2378 698218 -2346 698454
rect -2966 698134 -2346 698218
rect -2966 697898 -2934 698134
rect -2698 697898 -2614 698134
rect -2378 697898 -2346 698134
rect -2966 671454 -2346 697898
rect -2966 671218 -2934 671454
rect -2698 671218 -2614 671454
rect -2378 671218 -2346 671454
rect -2966 671134 -2346 671218
rect -2966 670898 -2934 671134
rect -2698 670898 -2614 671134
rect -2378 670898 -2346 671134
rect -2966 644454 -2346 670898
rect -2966 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 -2346 644454
rect -2966 644134 -2346 644218
rect -2966 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 -2346 644134
rect -2966 617454 -2346 643898
rect -2966 617218 -2934 617454
rect -2698 617218 -2614 617454
rect -2378 617218 -2346 617454
rect -2966 617134 -2346 617218
rect -2966 616898 -2934 617134
rect -2698 616898 -2614 617134
rect -2378 616898 -2346 617134
rect -2966 590454 -2346 616898
rect -2966 590218 -2934 590454
rect -2698 590218 -2614 590454
rect -2378 590218 -2346 590454
rect -2966 590134 -2346 590218
rect -2966 589898 -2934 590134
rect -2698 589898 -2614 590134
rect -2378 589898 -2346 590134
rect -2966 563454 -2346 589898
rect -2966 563218 -2934 563454
rect -2698 563218 -2614 563454
rect -2378 563218 -2346 563454
rect -2966 563134 -2346 563218
rect -2966 562898 -2934 563134
rect -2698 562898 -2614 563134
rect -2378 562898 -2346 563134
rect -2966 536454 -2346 562898
rect -2966 536218 -2934 536454
rect -2698 536218 -2614 536454
rect -2378 536218 -2346 536454
rect -2966 536134 -2346 536218
rect -2966 535898 -2934 536134
rect -2698 535898 -2614 536134
rect -2378 535898 -2346 536134
rect -2966 509454 -2346 535898
rect -2966 509218 -2934 509454
rect -2698 509218 -2614 509454
rect -2378 509218 -2346 509454
rect -2966 509134 -2346 509218
rect -2966 508898 -2934 509134
rect -2698 508898 -2614 509134
rect -2378 508898 -2346 509134
rect -2966 482454 -2346 508898
rect -2966 482218 -2934 482454
rect -2698 482218 -2614 482454
rect -2378 482218 -2346 482454
rect -2966 482134 -2346 482218
rect -2966 481898 -2934 482134
rect -2698 481898 -2614 482134
rect -2378 481898 -2346 482134
rect -2966 455454 -2346 481898
rect -2966 455218 -2934 455454
rect -2698 455218 -2614 455454
rect -2378 455218 -2346 455454
rect -2966 455134 -2346 455218
rect -2966 454898 -2934 455134
rect -2698 454898 -2614 455134
rect -2378 454898 -2346 455134
rect -2966 428454 -2346 454898
rect -2966 428218 -2934 428454
rect -2698 428218 -2614 428454
rect -2378 428218 -2346 428454
rect -2966 428134 -2346 428218
rect -2966 427898 -2934 428134
rect -2698 427898 -2614 428134
rect -2378 427898 -2346 428134
rect -2966 401454 -2346 427898
rect -2966 401218 -2934 401454
rect -2698 401218 -2614 401454
rect -2378 401218 -2346 401454
rect -2966 401134 -2346 401218
rect -2966 400898 -2934 401134
rect -2698 400898 -2614 401134
rect -2378 400898 -2346 401134
rect -2966 374454 -2346 400898
rect -2966 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 -2346 374454
rect -2966 374134 -2346 374218
rect -2966 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 -2346 374134
rect -2966 347454 -2346 373898
rect -2966 347218 -2934 347454
rect -2698 347218 -2614 347454
rect -2378 347218 -2346 347454
rect -2966 347134 -2346 347218
rect -2966 346898 -2934 347134
rect -2698 346898 -2614 347134
rect -2378 346898 -2346 347134
rect -2966 320454 -2346 346898
rect -2966 320218 -2934 320454
rect -2698 320218 -2614 320454
rect -2378 320218 -2346 320454
rect -2966 320134 -2346 320218
rect -2966 319898 -2934 320134
rect -2698 319898 -2614 320134
rect -2378 319898 -2346 320134
rect -2966 293454 -2346 319898
rect -2966 293218 -2934 293454
rect -2698 293218 -2614 293454
rect -2378 293218 -2346 293454
rect -2966 293134 -2346 293218
rect -2966 292898 -2934 293134
rect -2698 292898 -2614 293134
rect -2378 292898 -2346 293134
rect -2966 266454 -2346 292898
rect -2966 266218 -2934 266454
rect -2698 266218 -2614 266454
rect -2378 266218 -2346 266454
rect -2966 266134 -2346 266218
rect -2966 265898 -2934 266134
rect -2698 265898 -2614 266134
rect -2378 265898 -2346 266134
rect -2966 239454 -2346 265898
rect -2966 239218 -2934 239454
rect -2698 239218 -2614 239454
rect -2378 239218 -2346 239454
rect -2966 239134 -2346 239218
rect -2966 238898 -2934 239134
rect -2698 238898 -2614 239134
rect -2378 238898 -2346 239134
rect -2966 212454 -2346 238898
rect -2966 212218 -2934 212454
rect -2698 212218 -2614 212454
rect -2378 212218 -2346 212454
rect -2966 212134 -2346 212218
rect -2966 211898 -2934 212134
rect -2698 211898 -2614 212134
rect -2378 211898 -2346 212134
rect -2966 185454 -2346 211898
rect -2966 185218 -2934 185454
rect -2698 185218 -2614 185454
rect -2378 185218 -2346 185454
rect -2966 185134 -2346 185218
rect -2966 184898 -2934 185134
rect -2698 184898 -2614 185134
rect -2378 184898 -2346 185134
rect -2966 158454 -2346 184898
rect -2966 158218 -2934 158454
rect -2698 158218 -2614 158454
rect -2378 158218 -2346 158454
rect -2966 158134 -2346 158218
rect -2966 157898 -2934 158134
rect -2698 157898 -2614 158134
rect -2378 157898 -2346 158134
rect -2966 131454 -2346 157898
rect -2966 131218 -2934 131454
rect -2698 131218 -2614 131454
rect -2378 131218 -2346 131454
rect -2966 131134 -2346 131218
rect -2966 130898 -2934 131134
rect -2698 130898 -2614 131134
rect -2378 130898 -2346 131134
rect -2966 104454 -2346 130898
rect -2966 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 -2346 104454
rect -2966 104134 -2346 104218
rect -2966 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 -2346 104134
rect -2966 77454 -2346 103898
rect -2966 77218 -2934 77454
rect -2698 77218 -2614 77454
rect -2378 77218 -2346 77454
rect -2966 77134 -2346 77218
rect -2966 76898 -2934 77134
rect -2698 76898 -2614 77134
rect -2378 76898 -2346 77134
rect -2966 50454 -2346 76898
rect -2966 50218 -2934 50454
rect -2698 50218 -2614 50454
rect -2378 50218 -2346 50454
rect -2966 50134 -2346 50218
rect -2966 49898 -2934 50134
rect -2698 49898 -2614 50134
rect -2378 49898 -2346 50134
rect -2966 23454 -2346 49898
rect -2966 23218 -2934 23454
rect -2698 23218 -2614 23454
rect -2378 23218 -2346 23454
rect -2966 23134 -2346 23218
rect -2966 22898 -2934 23134
rect -2698 22898 -2614 23134
rect -2378 22898 -2346 23134
rect -2966 -1306 -2346 22898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 701829 -1386 704282
rect -2006 701593 -1974 701829
rect -1738 701593 -1654 701829
rect -1418 701593 -1386 701829
rect -2006 701509 -1386 701593
rect -2006 701273 -1974 701509
rect -1738 701273 -1654 701509
rect -1418 701273 -1386 701509
rect -2006 674829 -1386 701273
rect 37994 698454 38614 705242
rect 37994 698218 38026 698454
rect 38262 698218 38346 698454
rect 38582 698218 38614 698454
rect 37994 698134 38614 698218
rect 37994 697898 38026 698134
rect 38262 697898 38346 698134
rect 38582 697898 38614 698134
rect 3371 684316 3437 684317
rect 3371 684252 3372 684316
rect 3436 684252 3437 684316
rect 3371 684251 3437 684252
rect -2006 674593 -1974 674829
rect -1738 674593 -1654 674829
rect -1418 674593 -1386 674829
rect -2006 674509 -1386 674593
rect -2006 674273 -1974 674509
rect -1738 674273 -1654 674509
rect -1418 674273 -1386 674509
rect -2006 647829 -1386 674273
rect -2006 647593 -1974 647829
rect -1738 647593 -1654 647829
rect -1418 647593 -1386 647829
rect -2006 647509 -1386 647593
rect -2006 647273 -1974 647509
rect -1738 647273 -1654 647509
rect -1418 647273 -1386 647509
rect -2006 620829 -1386 647273
rect -2006 620593 -1974 620829
rect -1738 620593 -1654 620829
rect -1418 620593 -1386 620829
rect -2006 620509 -1386 620593
rect -2006 620273 -1974 620509
rect -1738 620273 -1654 620509
rect -1418 620273 -1386 620509
rect -2006 593829 -1386 620273
rect -2006 593593 -1974 593829
rect -1738 593593 -1654 593829
rect -1418 593593 -1386 593829
rect -2006 593509 -1386 593593
rect -2006 593273 -1974 593509
rect -1738 593273 -1654 593509
rect -1418 593273 -1386 593509
rect -2006 566829 -1386 593273
rect -2006 566593 -1974 566829
rect -1738 566593 -1654 566829
rect -1418 566593 -1386 566829
rect -2006 566509 -1386 566593
rect -2006 566273 -1974 566509
rect -1738 566273 -1654 566509
rect -1418 566273 -1386 566509
rect -2006 539829 -1386 566273
rect -2006 539593 -1974 539829
rect -1738 539593 -1654 539829
rect -1418 539593 -1386 539829
rect -2006 539509 -1386 539593
rect -2006 539273 -1974 539509
rect -1738 539273 -1654 539509
rect -1418 539273 -1386 539509
rect -2006 512829 -1386 539273
rect -2006 512593 -1974 512829
rect -1738 512593 -1654 512829
rect -1418 512593 -1386 512829
rect -2006 512509 -1386 512593
rect -2006 512273 -1974 512509
rect -1738 512273 -1654 512509
rect -1418 512273 -1386 512509
rect -2006 485829 -1386 512273
rect -2006 485593 -1974 485829
rect -1738 485593 -1654 485829
rect -1418 485593 -1386 485829
rect -2006 485509 -1386 485593
rect -2006 485273 -1974 485509
rect -1738 485273 -1654 485509
rect -1418 485273 -1386 485509
rect -2006 458829 -1386 485273
rect -2006 458593 -1974 458829
rect -1738 458593 -1654 458829
rect -1418 458593 -1386 458829
rect -2006 458509 -1386 458593
rect -2006 458273 -1974 458509
rect -1738 458273 -1654 458509
rect -1418 458273 -1386 458509
rect -2006 431829 -1386 458273
rect -2006 431593 -1974 431829
rect -1738 431593 -1654 431829
rect -1418 431593 -1386 431829
rect -2006 431509 -1386 431593
rect -2006 431273 -1974 431509
rect -1738 431273 -1654 431509
rect -1418 431273 -1386 431509
rect -2006 404829 -1386 431273
rect -2006 404593 -1974 404829
rect -1738 404593 -1654 404829
rect -1418 404593 -1386 404829
rect -2006 404509 -1386 404593
rect -2006 404273 -1974 404509
rect -1738 404273 -1654 404509
rect -1418 404273 -1386 404509
rect -2006 377829 -1386 404273
rect -2006 377593 -1974 377829
rect -1738 377593 -1654 377829
rect -1418 377593 -1386 377829
rect -2006 377509 -1386 377593
rect -2006 377273 -1974 377509
rect -1738 377273 -1654 377509
rect -1418 377273 -1386 377509
rect -2006 350829 -1386 377273
rect -2006 350593 -1974 350829
rect -1738 350593 -1654 350829
rect -1418 350593 -1386 350829
rect -2006 350509 -1386 350593
rect -2006 350273 -1974 350509
rect -1738 350273 -1654 350509
rect -1418 350273 -1386 350509
rect -2006 323829 -1386 350273
rect -2006 323593 -1974 323829
rect -1738 323593 -1654 323829
rect -1418 323593 -1386 323829
rect -2006 323509 -1386 323593
rect -2006 323273 -1974 323509
rect -1738 323273 -1654 323509
rect -1418 323273 -1386 323509
rect -2006 296829 -1386 323273
rect -2006 296593 -1974 296829
rect -1738 296593 -1654 296829
rect -1418 296593 -1386 296829
rect -2006 296509 -1386 296593
rect -2006 296273 -1974 296509
rect -1738 296273 -1654 296509
rect -1418 296273 -1386 296509
rect -2006 269829 -1386 296273
rect -2006 269593 -1974 269829
rect -1738 269593 -1654 269829
rect -1418 269593 -1386 269829
rect -2006 269509 -1386 269593
rect -2006 269273 -1974 269509
rect -1738 269273 -1654 269509
rect -1418 269273 -1386 269509
rect -2006 242829 -1386 269273
rect -2006 242593 -1974 242829
rect -1738 242593 -1654 242829
rect -1418 242593 -1386 242829
rect -2006 242509 -1386 242593
rect -2006 242273 -1974 242509
rect -1738 242273 -1654 242509
rect -1418 242273 -1386 242509
rect -2006 215829 -1386 242273
rect -2006 215593 -1974 215829
rect -1738 215593 -1654 215829
rect -1418 215593 -1386 215829
rect -2006 215509 -1386 215593
rect -2006 215273 -1974 215509
rect -1738 215273 -1654 215509
rect -1418 215273 -1386 215509
rect -2006 188829 -1386 215273
rect -2006 188593 -1974 188829
rect -1738 188593 -1654 188829
rect -1418 188593 -1386 188829
rect -2006 188509 -1386 188593
rect -2006 188273 -1974 188509
rect -1738 188273 -1654 188509
rect -1418 188273 -1386 188509
rect -2006 161829 -1386 188273
rect -2006 161593 -1974 161829
rect -1738 161593 -1654 161829
rect -1418 161593 -1386 161829
rect -2006 161509 -1386 161593
rect -2006 161273 -1974 161509
rect -1738 161273 -1654 161509
rect -1418 161273 -1386 161509
rect -2006 134829 -1386 161273
rect -2006 134593 -1974 134829
rect -1738 134593 -1654 134829
rect -1418 134593 -1386 134829
rect -2006 134509 -1386 134593
rect -2006 134273 -1974 134509
rect -1738 134273 -1654 134509
rect -1418 134273 -1386 134509
rect -2006 107829 -1386 134273
rect -2006 107593 -1974 107829
rect -1738 107593 -1654 107829
rect -1418 107593 -1386 107829
rect -2006 107509 -1386 107593
rect -2006 107273 -1974 107509
rect -1738 107273 -1654 107509
rect -1418 107273 -1386 107509
rect -2006 80829 -1386 107273
rect -2006 80593 -1974 80829
rect -1738 80593 -1654 80829
rect -1418 80593 -1386 80829
rect -2006 80509 -1386 80593
rect -2006 80273 -1974 80509
rect -1738 80273 -1654 80509
rect -1418 80273 -1386 80509
rect -2006 53829 -1386 80273
rect -2006 53593 -1974 53829
rect -1738 53593 -1654 53829
rect -1418 53593 -1386 53829
rect -2006 53509 -1386 53593
rect -2006 53273 -1974 53509
rect -1738 53273 -1654 53509
rect -1418 53273 -1386 53509
rect -2006 26829 -1386 53273
rect 3374 37909 3434 684251
rect 37994 671454 38614 697898
rect 37994 671218 38026 671454
rect 38262 671218 38346 671454
rect 38582 671218 38614 671454
rect 37994 671134 38614 671218
rect 37994 670898 38026 671134
rect 38262 670898 38346 671134
rect 38582 670898 38614 671134
rect 37994 644454 38614 670898
rect 37994 644218 38026 644454
rect 38262 644218 38346 644454
rect 38582 644218 38614 644454
rect 37994 644134 38614 644218
rect 37994 643898 38026 644134
rect 38262 643898 38346 644134
rect 38582 643898 38614 644134
rect 37994 617454 38614 643898
rect 37994 617218 38026 617454
rect 38262 617218 38346 617454
rect 38582 617218 38614 617454
rect 37994 617134 38614 617218
rect 37994 616898 38026 617134
rect 38262 616898 38346 617134
rect 38582 616898 38614 617134
rect 3555 606116 3621 606117
rect 3555 606052 3556 606116
rect 3620 606052 3621 606116
rect 3555 606051 3621 606052
rect 3371 37908 3437 37909
rect 3371 37844 3372 37908
rect 3436 37844 3437 37908
rect 3371 37843 3437 37844
rect -2006 26593 -1974 26829
rect -1738 26593 -1654 26829
rect -1418 26593 -1386 26829
rect -2006 26509 -1386 26593
rect -2006 26273 -1974 26509
rect -1738 26273 -1654 26509
rect -1418 26273 -1386 26509
rect -2006 -346 -1386 26273
rect 3558 13565 3618 606051
rect 37994 590454 38614 616898
rect 37994 590218 38026 590454
rect 38262 590218 38346 590454
rect 38582 590218 38614 590454
rect 37994 590134 38614 590218
rect 37994 589898 38026 590134
rect 38262 589898 38346 590134
rect 38582 589898 38614 590134
rect 37994 563454 38614 589898
rect 37994 563218 38026 563454
rect 38262 563218 38346 563454
rect 38582 563218 38614 563454
rect 37994 563134 38614 563218
rect 37994 562898 38026 563134
rect 38262 562898 38346 563134
rect 38582 562898 38614 563134
rect 37994 536454 38614 562898
rect 37994 536218 38026 536454
rect 38262 536218 38346 536454
rect 38582 536218 38614 536454
rect 37994 536134 38614 536218
rect 37994 535898 38026 536134
rect 38262 535898 38346 536134
rect 38582 535898 38614 536134
rect 37994 509454 38614 535898
rect 37994 509218 38026 509454
rect 38262 509218 38346 509454
rect 38582 509218 38614 509454
rect 37994 509134 38614 509218
rect 37994 508898 38026 509134
rect 38262 508898 38346 509134
rect 38582 508898 38614 509134
rect 37994 482454 38614 508898
rect 37994 482218 38026 482454
rect 38262 482218 38346 482454
rect 38582 482218 38614 482454
rect 37994 482134 38614 482218
rect 37994 481898 38026 482134
rect 38262 481898 38346 482134
rect 38582 481898 38614 482134
rect 37994 455454 38614 481898
rect 37994 455218 38026 455454
rect 38262 455218 38346 455454
rect 38582 455218 38614 455454
rect 37994 455134 38614 455218
rect 37994 454898 38026 455134
rect 38262 454898 38346 455134
rect 38582 454898 38614 455134
rect 37994 428454 38614 454898
rect 37994 428218 38026 428454
rect 38262 428218 38346 428454
rect 38582 428218 38614 428454
rect 37994 428134 38614 428218
rect 37994 427898 38026 428134
rect 38262 427898 38346 428134
rect 38582 427898 38614 428134
rect 37994 401454 38614 427898
rect 37994 401218 38026 401454
rect 38262 401218 38346 401454
rect 38582 401218 38614 401454
rect 37994 401134 38614 401218
rect 37994 400898 38026 401134
rect 38262 400898 38346 401134
rect 38582 400898 38614 401134
rect 37994 374454 38614 400898
rect 37994 374218 38026 374454
rect 38262 374218 38346 374454
rect 38582 374218 38614 374454
rect 37994 374134 38614 374218
rect 37994 373898 38026 374134
rect 38262 373898 38346 374134
rect 38582 373898 38614 374134
rect 37994 347454 38614 373898
rect 37994 347218 38026 347454
rect 38262 347218 38346 347454
rect 38582 347218 38614 347454
rect 37994 347134 38614 347218
rect 37994 346898 38026 347134
rect 38262 346898 38346 347134
rect 38582 346898 38614 347134
rect 37994 320454 38614 346898
rect 37994 320218 38026 320454
rect 38262 320218 38346 320454
rect 38582 320218 38614 320454
rect 37994 320134 38614 320218
rect 37994 319898 38026 320134
rect 38262 319898 38346 320134
rect 38582 319898 38614 320134
rect 37994 293454 38614 319898
rect 37994 293218 38026 293454
rect 38262 293218 38346 293454
rect 38582 293218 38614 293454
rect 37994 293134 38614 293218
rect 37994 292898 38026 293134
rect 38262 292898 38346 293134
rect 38582 292898 38614 293134
rect 37994 266454 38614 292898
rect 37994 266218 38026 266454
rect 38262 266218 38346 266454
rect 38582 266218 38614 266454
rect 37994 266134 38614 266218
rect 37994 265898 38026 266134
rect 38262 265898 38346 266134
rect 38582 265898 38614 266134
rect 37994 239454 38614 265898
rect 37994 239218 38026 239454
rect 38262 239218 38346 239454
rect 38582 239218 38614 239454
rect 37994 239134 38614 239218
rect 37994 238898 38026 239134
rect 38262 238898 38346 239134
rect 38582 238898 38614 239134
rect 37994 212454 38614 238898
rect 37994 212218 38026 212454
rect 38262 212218 38346 212454
rect 38582 212218 38614 212454
rect 37994 212134 38614 212218
rect 37994 211898 38026 212134
rect 38262 211898 38346 212134
rect 38582 211898 38614 212134
rect 37994 185454 38614 211898
rect 37994 185218 38026 185454
rect 38262 185218 38346 185454
rect 38582 185218 38614 185454
rect 37994 185134 38614 185218
rect 37994 184898 38026 185134
rect 38262 184898 38346 185134
rect 38582 184898 38614 185134
rect 37994 158454 38614 184898
rect 37994 158218 38026 158454
rect 38262 158218 38346 158454
rect 38582 158218 38614 158454
rect 37994 158134 38614 158218
rect 37994 157898 38026 158134
rect 38262 157898 38346 158134
rect 38582 157898 38614 158134
rect 37994 131454 38614 157898
rect 37994 131218 38026 131454
rect 38262 131218 38346 131454
rect 38582 131218 38614 131454
rect 37994 131134 38614 131218
rect 37994 130898 38026 131134
rect 38262 130898 38346 131134
rect 38582 130898 38614 131134
rect 37994 104454 38614 130898
rect 37994 104218 38026 104454
rect 38262 104218 38346 104454
rect 38582 104218 38614 104454
rect 37994 104134 38614 104218
rect 37994 103898 38026 104134
rect 38262 103898 38346 104134
rect 38582 103898 38614 104134
rect 37994 77454 38614 103898
rect 37994 77218 38026 77454
rect 38262 77218 38346 77454
rect 38582 77218 38614 77454
rect 37994 77134 38614 77218
rect 37994 76898 38026 77134
rect 38262 76898 38346 77134
rect 38582 76898 38614 77134
rect 37994 50454 38614 76898
rect 37994 50218 38026 50454
rect 38262 50218 38346 50454
rect 38582 50218 38614 50454
rect 37994 50134 38614 50218
rect 37994 49898 38026 50134
rect 38262 49898 38346 50134
rect 38582 49898 38614 50134
rect 37994 38000 38614 49898
rect 41494 704838 42114 711590
rect 41494 704602 41526 704838
rect 41762 704602 41846 704838
rect 42082 704602 42114 704838
rect 41494 704518 42114 704602
rect 41494 704282 41526 704518
rect 41762 704282 41846 704518
rect 42082 704282 42114 704518
rect 41494 701829 42114 704282
rect 41494 701593 41526 701829
rect 41762 701593 41846 701829
rect 42082 701593 42114 701829
rect 41494 701509 42114 701593
rect 41494 701273 41526 701509
rect 41762 701273 41846 701509
rect 42082 701273 42114 701509
rect 41494 674829 42114 701273
rect 41494 674593 41526 674829
rect 41762 674593 41846 674829
rect 42082 674593 42114 674829
rect 41494 674509 42114 674593
rect 41494 674273 41526 674509
rect 41762 674273 41846 674509
rect 42082 674273 42114 674509
rect 41494 647829 42114 674273
rect 41494 647593 41526 647829
rect 41762 647593 41846 647829
rect 42082 647593 42114 647829
rect 41494 647509 42114 647593
rect 41494 647273 41526 647509
rect 41762 647273 41846 647509
rect 42082 647273 42114 647509
rect 41494 620829 42114 647273
rect 41494 620593 41526 620829
rect 41762 620593 41846 620829
rect 42082 620593 42114 620829
rect 41494 620509 42114 620593
rect 41494 620273 41526 620509
rect 41762 620273 41846 620509
rect 42082 620273 42114 620509
rect 41494 593829 42114 620273
rect 41494 593593 41526 593829
rect 41762 593593 41846 593829
rect 42082 593593 42114 593829
rect 41494 593509 42114 593593
rect 41494 593273 41526 593509
rect 41762 593273 41846 593509
rect 42082 593273 42114 593509
rect 41494 566829 42114 593273
rect 41494 566593 41526 566829
rect 41762 566593 41846 566829
rect 42082 566593 42114 566829
rect 41494 566509 42114 566593
rect 41494 566273 41526 566509
rect 41762 566273 41846 566509
rect 42082 566273 42114 566509
rect 41494 539829 42114 566273
rect 41494 539593 41526 539829
rect 41762 539593 41846 539829
rect 42082 539593 42114 539829
rect 41494 539509 42114 539593
rect 41494 539273 41526 539509
rect 41762 539273 41846 539509
rect 42082 539273 42114 539509
rect 41494 512829 42114 539273
rect 41494 512593 41526 512829
rect 41762 512593 41846 512829
rect 42082 512593 42114 512829
rect 41494 512509 42114 512593
rect 41494 512273 41526 512509
rect 41762 512273 41846 512509
rect 42082 512273 42114 512509
rect 41494 485829 42114 512273
rect 65994 705798 66614 711590
rect 65994 705562 66026 705798
rect 66262 705562 66346 705798
rect 66582 705562 66614 705798
rect 65994 705478 66614 705562
rect 65994 705242 66026 705478
rect 66262 705242 66346 705478
rect 66582 705242 66614 705478
rect 65994 698454 66614 705242
rect 65994 698218 66026 698454
rect 66262 698218 66346 698454
rect 66582 698218 66614 698454
rect 65994 698134 66614 698218
rect 65994 697898 66026 698134
rect 66262 697898 66346 698134
rect 66582 697898 66614 698134
rect 65994 671454 66614 697898
rect 65994 671218 66026 671454
rect 66262 671218 66346 671454
rect 66582 671218 66614 671454
rect 65994 671134 66614 671218
rect 65994 670898 66026 671134
rect 66262 670898 66346 671134
rect 66582 670898 66614 671134
rect 65994 644454 66614 670898
rect 65994 644218 66026 644454
rect 66262 644218 66346 644454
rect 66582 644218 66614 644454
rect 65994 644134 66614 644218
rect 65994 643898 66026 644134
rect 66262 643898 66346 644134
rect 66582 643898 66614 644134
rect 65994 617454 66614 643898
rect 65994 617218 66026 617454
rect 66262 617218 66346 617454
rect 66582 617218 66614 617454
rect 65994 617134 66614 617218
rect 65994 616898 66026 617134
rect 66262 616898 66346 617134
rect 66582 616898 66614 617134
rect 65994 590454 66614 616898
rect 65994 590218 66026 590454
rect 66262 590218 66346 590454
rect 66582 590218 66614 590454
rect 65994 590134 66614 590218
rect 65994 589898 66026 590134
rect 66262 589898 66346 590134
rect 66582 589898 66614 590134
rect 65994 563454 66614 589898
rect 65994 563218 66026 563454
rect 66262 563218 66346 563454
rect 66582 563218 66614 563454
rect 65994 563134 66614 563218
rect 65994 562898 66026 563134
rect 66262 562898 66346 563134
rect 66582 562898 66614 563134
rect 65994 536454 66614 562898
rect 65994 536218 66026 536454
rect 66262 536218 66346 536454
rect 66582 536218 66614 536454
rect 65994 536134 66614 536218
rect 65994 535898 66026 536134
rect 66262 535898 66346 536134
rect 66582 535898 66614 536134
rect 65994 509454 66614 535898
rect 65994 509218 66026 509454
rect 66262 509218 66346 509454
rect 66582 509218 66614 509454
rect 65994 509134 66614 509218
rect 65994 508898 66026 509134
rect 66262 508898 66346 509134
rect 66582 508898 66614 509134
rect 45323 500988 45389 500989
rect 45323 500924 45324 500988
rect 45388 500924 45389 500988
rect 45323 500923 45389 500924
rect 41494 485593 41526 485829
rect 41762 485593 41846 485829
rect 42082 485593 42114 485829
rect 41494 485509 42114 485593
rect 41494 485273 41526 485509
rect 41762 485273 41846 485509
rect 42082 485273 42114 485509
rect 41494 458829 42114 485273
rect 41494 458593 41526 458829
rect 41762 458593 41846 458829
rect 42082 458593 42114 458829
rect 41494 458509 42114 458593
rect 41494 458273 41526 458509
rect 41762 458273 41846 458509
rect 42082 458273 42114 458509
rect 41494 431829 42114 458273
rect 41494 431593 41526 431829
rect 41762 431593 41846 431829
rect 42082 431593 42114 431829
rect 41494 431509 42114 431593
rect 41494 431273 41526 431509
rect 41762 431273 41846 431509
rect 42082 431273 42114 431509
rect 41494 404829 42114 431273
rect 41494 404593 41526 404829
rect 41762 404593 41846 404829
rect 42082 404593 42114 404829
rect 41494 404509 42114 404593
rect 41494 404273 41526 404509
rect 41762 404273 41846 404509
rect 42082 404273 42114 404509
rect 41494 377829 42114 404273
rect 41494 377593 41526 377829
rect 41762 377593 41846 377829
rect 42082 377593 42114 377829
rect 41494 377509 42114 377593
rect 41494 377273 41526 377509
rect 41762 377273 41846 377509
rect 42082 377273 42114 377509
rect 41494 350829 42114 377273
rect 41494 350593 41526 350829
rect 41762 350593 41846 350829
rect 42082 350593 42114 350829
rect 41494 350509 42114 350593
rect 41494 350273 41526 350509
rect 41762 350273 41846 350509
rect 42082 350273 42114 350509
rect 41494 323829 42114 350273
rect 41494 323593 41526 323829
rect 41762 323593 41846 323829
rect 42082 323593 42114 323829
rect 41494 323509 42114 323593
rect 41494 323273 41526 323509
rect 41762 323273 41846 323509
rect 42082 323273 42114 323509
rect 41494 296829 42114 323273
rect 41494 296593 41526 296829
rect 41762 296593 41846 296829
rect 42082 296593 42114 296829
rect 41494 296509 42114 296593
rect 41494 296273 41526 296509
rect 41762 296273 41846 296509
rect 42082 296273 42114 296509
rect 41494 269829 42114 296273
rect 41494 269593 41526 269829
rect 41762 269593 41846 269829
rect 42082 269593 42114 269829
rect 41494 269509 42114 269593
rect 41494 269273 41526 269509
rect 41762 269273 41846 269509
rect 42082 269273 42114 269509
rect 41494 242829 42114 269273
rect 41494 242593 41526 242829
rect 41762 242593 41846 242829
rect 42082 242593 42114 242829
rect 41494 242509 42114 242593
rect 41494 242273 41526 242509
rect 41762 242273 41846 242509
rect 42082 242273 42114 242509
rect 41494 215829 42114 242273
rect 41494 215593 41526 215829
rect 41762 215593 41846 215829
rect 42082 215593 42114 215829
rect 41494 215509 42114 215593
rect 41494 215273 41526 215509
rect 41762 215273 41846 215509
rect 42082 215273 42114 215509
rect 41494 188829 42114 215273
rect 41494 188593 41526 188829
rect 41762 188593 41846 188829
rect 42082 188593 42114 188829
rect 41494 188509 42114 188593
rect 41494 188273 41526 188509
rect 41762 188273 41846 188509
rect 42082 188273 42114 188509
rect 41494 161829 42114 188273
rect 41494 161593 41526 161829
rect 41762 161593 41846 161829
rect 42082 161593 42114 161829
rect 41494 161509 42114 161593
rect 41494 161273 41526 161509
rect 41762 161273 41846 161509
rect 42082 161273 42114 161509
rect 41494 134829 42114 161273
rect 41494 134593 41526 134829
rect 41762 134593 41846 134829
rect 42082 134593 42114 134829
rect 41494 134509 42114 134593
rect 41494 134273 41526 134509
rect 41762 134273 41846 134509
rect 42082 134273 42114 134509
rect 41494 107829 42114 134273
rect 41494 107593 41526 107829
rect 41762 107593 41846 107829
rect 42082 107593 42114 107829
rect 41494 107509 42114 107593
rect 41494 107273 41526 107509
rect 41762 107273 41846 107509
rect 42082 107273 42114 107509
rect 41494 80829 42114 107273
rect 41494 80593 41526 80829
rect 41762 80593 41846 80829
rect 42082 80593 42114 80829
rect 41494 80509 42114 80593
rect 41494 80273 41526 80509
rect 41762 80273 41846 80509
rect 42082 80273 42114 80509
rect 41494 53829 42114 80273
rect 41494 53593 41526 53829
rect 41762 53593 41846 53829
rect 42082 53593 42114 53829
rect 41494 53509 42114 53593
rect 41494 53273 41526 53509
rect 41762 53273 41846 53509
rect 42082 53273 42114 53509
rect 41494 38000 42114 53273
rect 39803 35324 39869 35325
rect 39803 35260 39804 35324
rect 39868 35260 39869 35324
rect 39803 35259 39869 35260
rect 42747 35324 42813 35325
rect 42747 35260 42748 35324
rect 42812 35260 42813 35324
rect 42747 35259 42813 35260
rect 22418 26829 22738 26861
rect 22418 26593 22460 26829
rect 22696 26593 22738 26829
rect 22418 26509 22738 26593
rect 22418 26273 22460 26509
rect 22696 26273 22738 26509
rect 22418 26241 22738 26273
rect 33366 26829 33686 26861
rect 33366 26593 33408 26829
rect 33644 26593 33686 26829
rect 33366 26509 33686 26593
rect 33366 26273 33408 26509
rect 33644 26273 33686 26509
rect 33366 26241 33686 26273
rect 27892 23454 28212 23486
rect 27892 23218 27934 23454
rect 28170 23218 28212 23454
rect 27892 23134 28212 23218
rect 27892 22898 27934 23134
rect 28170 22898 28212 23134
rect 27892 22866 28212 22898
rect 38840 23454 39160 23486
rect 38840 23218 38882 23454
rect 39118 23218 39160 23454
rect 38840 23134 39160 23218
rect 38840 22898 38882 23134
rect 39118 22898 39160 23134
rect 38840 22866 39160 22898
rect 3555 13564 3621 13565
rect 3555 13500 3556 13564
rect 3620 13500 3621 13564
rect 3555 13499 3621 13500
rect 39806 3365 39866 35259
rect 42750 5677 42810 35259
rect 44314 26829 44634 26861
rect 44314 26593 44356 26829
rect 44592 26593 44634 26829
rect 44314 26509 44634 26593
rect 44314 26273 44356 26509
rect 44592 26273 44634 26509
rect 44314 26241 44634 26273
rect 45326 16590 45386 500923
rect 65994 482454 66614 508898
rect 65994 482218 66026 482454
rect 66262 482218 66346 482454
rect 66582 482218 66614 482454
rect 65994 482134 66614 482218
rect 65994 481898 66026 482134
rect 66262 481898 66346 482134
rect 66582 481898 66614 482134
rect 54339 474876 54405 474877
rect 54339 474812 54340 474876
rect 54404 474812 54405 474876
rect 54339 474811 54405 474812
rect 50843 35324 50909 35325
rect 50843 35260 50844 35324
rect 50908 35260 50909 35324
rect 50843 35259 50909 35260
rect 49788 23454 50108 23486
rect 49788 23218 49830 23454
rect 50066 23218 50108 23454
rect 49788 23134 50108 23218
rect 49788 22898 49830 23134
rect 50066 22898 50108 23134
rect 49788 22866 50108 22898
rect 45326 16557 45570 16590
rect 45326 16556 45573 16557
rect 45326 16530 45508 16556
rect 45507 16492 45508 16530
rect 45572 16492 45573 16556
rect 45507 16491 45573 16492
rect 42747 5676 42813 5677
rect 42747 5612 42748 5676
rect 42812 5612 42813 5676
rect 42747 5611 42813 5612
rect 50846 3501 50906 35259
rect 54342 16557 54402 474811
rect 65994 455454 66614 481898
rect 65994 455218 66026 455454
rect 66262 455218 66346 455454
rect 66582 455218 66614 455454
rect 65994 455134 66614 455218
rect 65994 454898 66026 455134
rect 66262 454898 66346 455134
rect 66582 454898 66614 455134
rect 65994 428454 66614 454898
rect 65994 428218 66026 428454
rect 66262 428218 66346 428454
rect 66582 428218 66614 428454
rect 65994 428134 66614 428218
rect 65994 427898 66026 428134
rect 66262 427898 66346 428134
rect 66582 427898 66614 428134
rect 65994 401454 66614 427898
rect 65994 401218 66026 401454
rect 66262 401218 66346 401454
rect 66582 401218 66614 401454
rect 65994 401134 66614 401218
rect 65994 400898 66026 401134
rect 66262 400898 66346 401134
rect 66582 400898 66614 401134
rect 65994 374454 66614 400898
rect 65994 374218 66026 374454
rect 66262 374218 66346 374454
rect 66582 374218 66614 374454
rect 65994 374134 66614 374218
rect 65994 373898 66026 374134
rect 66262 373898 66346 374134
rect 66582 373898 66614 374134
rect 65994 347454 66614 373898
rect 65994 347218 66026 347454
rect 66262 347218 66346 347454
rect 66582 347218 66614 347454
rect 65994 347134 66614 347218
rect 65994 346898 66026 347134
rect 66262 346898 66346 347134
rect 66582 346898 66614 347134
rect 65994 320454 66614 346898
rect 65994 320218 66026 320454
rect 66262 320218 66346 320454
rect 66582 320218 66614 320454
rect 65994 320134 66614 320218
rect 65994 319898 66026 320134
rect 66262 319898 66346 320134
rect 66582 319898 66614 320134
rect 65994 293454 66614 319898
rect 65994 293218 66026 293454
rect 66262 293218 66346 293454
rect 66582 293218 66614 293454
rect 65994 293134 66614 293218
rect 65994 292898 66026 293134
rect 66262 292898 66346 293134
rect 66582 292898 66614 293134
rect 65994 266454 66614 292898
rect 65994 266218 66026 266454
rect 66262 266218 66346 266454
rect 66582 266218 66614 266454
rect 65994 266134 66614 266218
rect 65994 265898 66026 266134
rect 66262 265898 66346 266134
rect 66582 265898 66614 266134
rect 65994 239454 66614 265898
rect 65994 239218 66026 239454
rect 66262 239218 66346 239454
rect 66582 239218 66614 239454
rect 65994 239134 66614 239218
rect 65994 238898 66026 239134
rect 66262 238898 66346 239134
rect 66582 238898 66614 239134
rect 65994 212454 66614 238898
rect 65994 212218 66026 212454
rect 66262 212218 66346 212454
rect 66582 212218 66614 212454
rect 65994 212134 66614 212218
rect 65994 211898 66026 212134
rect 66262 211898 66346 212134
rect 66582 211898 66614 212134
rect 65994 185454 66614 211898
rect 65994 185218 66026 185454
rect 66262 185218 66346 185454
rect 66582 185218 66614 185454
rect 65994 185134 66614 185218
rect 65994 184898 66026 185134
rect 66262 184898 66346 185134
rect 66582 184898 66614 185134
rect 65994 158454 66614 184898
rect 65994 158218 66026 158454
rect 66262 158218 66346 158454
rect 66582 158218 66614 158454
rect 65994 158134 66614 158218
rect 65994 157898 66026 158134
rect 66262 157898 66346 158134
rect 66582 157898 66614 158134
rect 65994 131454 66614 157898
rect 65994 131218 66026 131454
rect 66262 131218 66346 131454
rect 66582 131218 66614 131454
rect 65994 131134 66614 131218
rect 65994 130898 66026 131134
rect 66262 130898 66346 131134
rect 66582 130898 66614 131134
rect 65994 104454 66614 130898
rect 65994 104218 66026 104454
rect 66262 104218 66346 104454
rect 66582 104218 66614 104454
rect 65994 104134 66614 104218
rect 65994 103898 66026 104134
rect 66262 103898 66346 104134
rect 66582 103898 66614 104134
rect 65994 77454 66614 103898
rect 65994 77218 66026 77454
rect 66262 77218 66346 77454
rect 66582 77218 66614 77454
rect 65994 77134 66614 77218
rect 65994 76898 66026 77134
rect 66262 76898 66346 77134
rect 66582 76898 66614 77134
rect 65994 50454 66614 76898
rect 65994 50218 66026 50454
rect 66262 50218 66346 50454
rect 66582 50218 66614 50454
rect 65994 50134 66614 50218
rect 65994 49898 66026 50134
rect 66262 49898 66346 50134
rect 66582 49898 66614 50134
rect 55262 26829 55582 26861
rect 55262 26593 55304 26829
rect 55540 26593 55582 26829
rect 55262 26509 55582 26593
rect 55262 26273 55304 26509
rect 55540 26273 55582 26509
rect 55262 26241 55582 26273
rect 60736 23454 61056 23486
rect 60736 23218 60778 23454
rect 61014 23218 61056 23454
rect 60736 23134 61056 23218
rect 60736 22898 60778 23134
rect 61014 22898 61056 23134
rect 60736 22866 61056 22898
rect 65994 23454 66614 49898
rect 65994 23218 66026 23454
rect 66262 23218 66346 23454
rect 66582 23218 66614 23454
rect 65994 23134 66614 23218
rect 65994 22898 66026 23134
rect 66262 22898 66346 23134
rect 66582 22898 66614 23134
rect 54339 16556 54405 16557
rect 54339 16492 54340 16556
rect 54404 16492 54405 16556
rect 54339 16491 54405 16492
rect 50843 3500 50909 3501
rect 50843 3436 50844 3500
rect 50908 3436 50909 3500
rect 50843 3435 50909 3436
rect 39803 3364 39869 3365
rect 39803 3300 39804 3364
rect 39868 3300 39869 3364
rect 39803 3299 39869 3300
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 65994 -1306 66614 22898
rect 65994 -1542 66026 -1306
rect 66262 -1542 66346 -1306
rect 66582 -1542 66614 -1306
rect 65994 -1626 66614 -1542
rect 65994 -1862 66026 -1626
rect 66262 -1862 66346 -1626
rect 66582 -1862 66614 -1626
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 65994 -7654 66614 -1862
rect 69494 704838 70114 711590
rect 69494 704602 69526 704838
rect 69762 704602 69846 704838
rect 70082 704602 70114 704838
rect 69494 704518 70114 704602
rect 69494 704282 69526 704518
rect 69762 704282 69846 704518
rect 70082 704282 70114 704518
rect 69494 701829 70114 704282
rect 69494 701593 69526 701829
rect 69762 701593 69846 701829
rect 70082 701593 70114 701829
rect 69494 701509 70114 701593
rect 69494 701273 69526 701509
rect 69762 701273 69846 701509
rect 70082 701273 70114 701509
rect 69494 674829 70114 701273
rect 69494 674593 69526 674829
rect 69762 674593 69846 674829
rect 70082 674593 70114 674829
rect 69494 674509 70114 674593
rect 69494 674273 69526 674509
rect 69762 674273 69846 674509
rect 70082 674273 70114 674509
rect 69494 647829 70114 674273
rect 69494 647593 69526 647829
rect 69762 647593 69846 647829
rect 70082 647593 70114 647829
rect 69494 647509 70114 647593
rect 69494 647273 69526 647509
rect 69762 647273 69846 647509
rect 70082 647273 70114 647509
rect 69494 620829 70114 647273
rect 69494 620593 69526 620829
rect 69762 620593 69846 620829
rect 70082 620593 70114 620829
rect 69494 620509 70114 620593
rect 69494 620273 69526 620509
rect 69762 620273 69846 620509
rect 70082 620273 70114 620509
rect 69494 593829 70114 620273
rect 69494 593593 69526 593829
rect 69762 593593 69846 593829
rect 70082 593593 70114 593829
rect 69494 593509 70114 593593
rect 69494 593273 69526 593509
rect 69762 593273 69846 593509
rect 70082 593273 70114 593509
rect 69494 566829 70114 593273
rect 69494 566593 69526 566829
rect 69762 566593 69846 566829
rect 70082 566593 70114 566829
rect 69494 566509 70114 566593
rect 69494 566273 69526 566509
rect 69762 566273 69846 566509
rect 70082 566273 70114 566509
rect 69494 539829 70114 566273
rect 69494 539593 69526 539829
rect 69762 539593 69846 539829
rect 70082 539593 70114 539829
rect 69494 539509 70114 539593
rect 69494 539273 69526 539509
rect 69762 539273 69846 539509
rect 70082 539273 70114 539509
rect 69494 512829 70114 539273
rect 69494 512593 69526 512829
rect 69762 512593 69846 512829
rect 70082 512593 70114 512829
rect 69494 512509 70114 512593
rect 69494 512273 69526 512509
rect 69762 512273 69846 512509
rect 70082 512273 70114 512509
rect 69494 485829 70114 512273
rect 69494 485593 69526 485829
rect 69762 485593 69846 485829
rect 70082 485593 70114 485829
rect 69494 485509 70114 485593
rect 69494 485273 69526 485509
rect 69762 485273 69846 485509
rect 70082 485273 70114 485509
rect 69494 458829 70114 485273
rect 69494 458593 69526 458829
rect 69762 458593 69846 458829
rect 70082 458593 70114 458829
rect 69494 458509 70114 458593
rect 69494 458273 69526 458509
rect 69762 458273 69846 458509
rect 70082 458273 70114 458509
rect 69494 431829 70114 458273
rect 69494 431593 69526 431829
rect 69762 431593 69846 431829
rect 70082 431593 70114 431829
rect 69494 431509 70114 431593
rect 69494 431273 69526 431509
rect 69762 431273 69846 431509
rect 70082 431273 70114 431509
rect 69494 404829 70114 431273
rect 69494 404593 69526 404829
rect 69762 404593 69846 404829
rect 70082 404593 70114 404829
rect 69494 404509 70114 404593
rect 69494 404273 69526 404509
rect 69762 404273 69846 404509
rect 70082 404273 70114 404509
rect 69494 377829 70114 404273
rect 69494 377593 69526 377829
rect 69762 377593 69846 377829
rect 70082 377593 70114 377829
rect 69494 377509 70114 377593
rect 69494 377273 69526 377509
rect 69762 377273 69846 377509
rect 70082 377273 70114 377509
rect 69494 350829 70114 377273
rect 69494 350593 69526 350829
rect 69762 350593 69846 350829
rect 70082 350593 70114 350829
rect 69494 350509 70114 350593
rect 69494 350273 69526 350509
rect 69762 350273 69846 350509
rect 70082 350273 70114 350509
rect 69494 323829 70114 350273
rect 69494 323593 69526 323829
rect 69762 323593 69846 323829
rect 70082 323593 70114 323829
rect 69494 323509 70114 323593
rect 69494 323273 69526 323509
rect 69762 323273 69846 323509
rect 70082 323273 70114 323509
rect 69494 296829 70114 323273
rect 69494 296593 69526 296829
rect 69762 296593 69846 296829
rect 70082 296593 70114 296829
rect 69494 296509 70114 296593
rect 69494 296273 69526 296509
rect 69762 296273 69846 296509
rect 70082 296273 70114 296509
rect 69494 269829 70114 296273
rect 69494 269593 69526 269829
rect 69762 269593 69846 269829
rect 70082 269593 70114 269829
rect 69494 269509 70114 269593
rect 69494 269273 69526 269509
rect 69762 269273 69846 269509
rect 70082 269273 70114 269509
rect 69494 242829 70114 269273
rect 69494 242593 69526 242829
rect 69762 242593 69846 242829
rect 70082 242593 70114 242829
rect 69494 242509 70114 242593
rect 69494 242273 69526 242509
rect 69762 242273 69846 242509
rect 70082 242273 70114 242509
rect 69494 215829 70114 242273
rect 69494 215593 69526 215829
rect 69762 215593 69846 215829
rect 70082 215593 70114 215829
rect 69494 215509 70114 215593
rect 69494 215273 69526 215509
rect 69762 215273 69846 215509
rect 70082 215273 70114 215509
rect 69494 188829 70114 215273
rect 69494 188593 69526 188829
rect 69762 188593 69846 188829
rect 70082 188593 70114 188829
rect 69494 188509 70114 188593
rect 69494 188273 69526 188509
rect 69762 188273 69846 188509
rect 70082 188273 70114 188509
rect 69494 161829 70114 188273
rect 69494 161593 69526 161829
rect 69762 161593 69846 161829
rect 70082 161593 70114 161829
rect 69494 161509 70114 161593
rect 69494 161273 69526 161509
rect 69762 161273 69846 161509
rect 70082 161273 70114 161509
rect 69494 134829 70114 161273
rect 69494 134593 69526 134829
rect 69762 134593 69846 134829
rect 70082 134593 70114 134829
rect 69494 134509 70114 134593
rect 69494 134273 69526 134509
rect 69762 134273 69846 134509
rect 70082 134273 70114 134509
rect 69494 107829 70114 134273
rect 69494 107593 69526 107829
rect 69762 107593 69846 107829
rect 70082 107593 70114 107829
rect 69494 107509 70114 107593
rect 69494 107273 69526 107509
rect 69762 107273 69846 107509
rect 70082 107273 70114 107509
rect 69494 80829 70114 107273
rect 69494 80593 69526 80829
rect 69762 80593 69846 80829
rect 70082 80593 70114 80829
rect 69494 80509 70114 80593
rect 69494 80273 69526 80509
rect 69762 80273 69846 80509
rect 70082 80273 70114 80509
rect 69494 53829 70114 80273
rect 69494 53593 69526 53829
rect 69762 53593 69846 53829
rect 70082 53593 70114 53829
rect 69494 53509 70114 53593
rect 69494 53273 69526 53509
rect 69762 53273 69846 53509
rect 70082 53273 70114 53509
rect 69494 26829 70114 53273
rect 93994 705798 94614 711590
rect 93994 705562 94026 705798
rect 94262 705562 94346 705798
rect 94582 705562 94614 705798
rect 93994 705478 94614 705562
rect 93994 705242 94026 705478
rect 94262 705242 94346 705478
rect 94582 705242 94614 705478
rect 93994 698454 94614 705242
rect 93994 698218 94026 698454
rect 94262 698218 94346 698454
rect 94582 698218 94614 698454
rect 93994 698134 94614 698218
rect 93994 697898 94026 698134
rect 94262 697898 94346 698134
rect 94582 697898 94614 698134
rect 93994 671454 94614 697898
rect 93994 671218 94026 671454
rect 94262 671218 94346 671454
rect 94582 671218 94614 671454
rect 93994 671134 94614 671218
rect 93994 670898 94026 671134
rect 94262 670898 94346 671134
rect 94582 670898 94614 671134
rect 93994 644454 94614 670898
rect 93994 644218 94026 644454
rect 94262 644218 94346 644454
rect 94582 644218 94614 644454
rect 93994 644134 94614 644218
rect 93994 643898 94026 644134
rect 94262 643898 94346 644134
rect 94582 643898 94614 644134
rect 93994 617454 94614 643898
rect 93994 617218 94026 617454
rect 94262 617218 94346 617454
rect 94582 617218 94614 617454
rect 93994 617134 94614 617218
rect 93994 616898 94026 617134
rect 94262 616898 94346 617134
rect 94582 616898 94614 617134
rect 93994 590454 94614 616898
rect 93994 590218 94026 590454
rect 94262 590218 94346 590454
rect 94582 590218 94614 590454
rect 93994 590134 94614 590218
rect 93994 589898 94026 590134
rect 94262 589898 94346 590134
rect 94582 589898 94614 590134
rect 93994 563454 94614 589898
rect 93994 563218 94026 563454
rect 94262 563218 94346 563454
rect 94582 563218 94614 563454
rect 93994 563134 94614 563218
rect 93994 562898 94026 563134
rect 94262 562898 94346 563134
rect 94582 562898 94614 563134
rect 93994 536454 94614 562898
rect 93994 536218 94026 536454
rect 94262 536218 94346 536454
rect 94582 536218 94614 536454
rect 93994 536134 94614 536218
rect 93994 535898 94026 536134
rect 94262 535898 94346 536134
rect 94582 535898 94614 536134
rect 93994 509454 94614 535898
rect 93994 509218 94026 509454
rect 94262 509218 94346 509454
rect 94582 509218 94614 509454
rect 93994 509134 94614 509218
rect 93994 508898 94026 509134
rect 94262 508898 94346 509134
rect 94582 508898 94614 509134
rect 93994 482454 94614 508898
rect 93994 482218 94026 482454
rect 94262 482218 94346 482454
rect 94582 482218 94614 482454
rect 93994 482134 94614 482218
rect 93994 481898 94026 482134
rect 94262 481898 94346 482134
rect 94582 481898 94614 482134
rect 93994 455454 94614 481898
rect 93994 455218 94026 455454
rect 94262 455218 94346 455454
rect 94582 455218 94614 455454
rect 93994 455134 94614 455218
rect 93994 454898 94026 455134
rect 94262 454898 94346 455134
rect 94582 454898 94614 455134
rect 93994 428454 94614 454898
rect 93994 428218 94026 428454
rect 94262 428218 94346 428454
rect 94582 428218 94614 428454
rect 93994 428134 94614 428218
rect 93994 427898 94026 428134
rect 94262 427898 94346 428134
rect 94582 427898 94614 428134
rect 93994 401454 94614 427898
rect 93994 401218 94026 401454
rect 94262 401218 94346 401454
rect 94582 401218 94614 401454
rect 93994 401134 94614 401218
rect 93994 400898 94026 401134
rect 94262 400898 94346 401134
rect 94582 400898 94614 401134
rect 93994 374454 94614 400898
rect 93994 374218 94026 374454
rect 94262 374218 94346 374454
rect 94582 374218 94614 374454
rect 93994 374134 94614 374218
rect 93994 373898 94026 374134
rect 94262 373898 94346 374134
rect 94582 373898 94614 374134
rect 93994 347454 94614 373898
rect 93994 347218 94026 347454
rect 94262 347218 94346 347454
rect 94582 347218 94614 347454
rect 93994 347134 94614 347218
rect 93994 346898 94026 347134
rect 94262 346898 94346 347134
rect 94582 346898 94614 347134
rect 93994 320454 94614 346898
rect 93994 320218 94026 320454
rect 94262 320218 94346 320454
rect 94582 320218 94614 320454
rect 93994 320134 94614 320218
rect 93994 319898 94026 320134
rect 94262 319898 94346 320134
rect 94582 319898 94614 320134
rect 93994 293454 94614 319898
rect 93994 293218 94026 293454
rect 94262 293218 94346 293454
rect 94582 293218 94614 293454
rect 93994 293134 94614 293218
rect 93994 292898 94026 293134
rect 94262 292898 94346 293134
rect 94582 292898 94614 293134
rect 93994 266454 94614 292898
rect 93994 266218 94026 266454
rect 94262 266218 94346 266454
rect 94582 266218 94614 266454
rect 93994 266134 94614 266218
rect 93994 265898 94026 266134
rect 94262 265898 94346 266134
rect 94582 265898 94614 266134
rect 93994 239454 94614 265898
rect 93994 239218 94026 239454
rect 94262 239218 94346 239454
rect 94582 239218 94614 239454
rect 93994 239134 94614 239218
rect 93994 238898 94026 239134
rect 94262 238898 94346 239134
rect 94582 238898 94614 239134
rect 93994 212454 94614 238898
rect 93994 212218 94026 212454
rect 94262 212218 94346 212454
rect 94582 212218 94614 212454
rect 93994 212134 94614 212218
rect 93994 211898 94026 212134
rect 94262 211898 94346 212134
rect 94582 211898 94614 212134
rect 93994 185454 94614 211898
rect 93994 185218 94026 185454
rect 94262 185218 94346 185454
rect 94582 185218 94614 185454
rect 93994 185134 94614 185218
rect 93994 184898 94026 185134
rect 94262 184898 94346 185134
rect 94582 184898 94614 185134
rect 93994 158454 94614 184898
rect 93994 158218 94026 158454
rect 94262 158218 94346 158454
rect 94582 158218 94614 158454
rect 93994 158134 94614 158218
rect 93994 157898 94026 158134
rect 94262 157898 94346 158134
rect 94582 157898 94614 158134
rect 93994 131454 94614 157898
rect 93994 131218 94026 131454
rect 94262 131218 94346 131454
rect 94582 131218 94614 131454
rect 93994 131134 94614 131218
rect 93994 130898 94026 131134
rect 94262 130898 94346 131134
rect 94582 130898 94614 131134
rect 93994 104454 94614 130898
rect 93994 104218 94026 104454
rect 94262 104218 94346 104454
rect 94582 104218 94614 104454
rect 93994 104134 94614 104218
rect 93994 103898 94026 104134
rect 94262 103898 94346 104134
rect 94582 103898 94614 104134
rect 93994 77454 94614 103898
rect 93994 77218 94026 77454
rect 94262 77218 94346 77454
rect 94582 77218 94614 77454
rect 93994 77134 94614 77218
rect 93994 76898 94026 77134
rect 94262 76898 94346 77134
rect 94582 76898 94614 77134
rect 93994 50454 94614 76898
rect 93994 50218 94026 50454
rect 94262 50218 94346 50454
rect 94582 50218 94614 50454
rect 93994 50134 94614 50218
rect 93994 49898 94026 50134
rect 94262 49898 94346 50134
rect 94582 49898 94614 50134
rect 93994 42000 94614 49898
rect 97494 704838 98114 711590
rect 97494 704602 97526 704838
rect 97762 704602 97846 704838
rect 98082 704602 98114 704838
rect 97494 704518 98114 704602
rect 97494 704282 97526 704518
rect 97762 704282 97846 704518
rect 98082 704282 98114 704518
rect 97494 701829 98114 704282
rect 97494 701593 97526 701829
rect 97762 701593 97846 701829
rect 98082 701593 98114 701829
rect 97494 701509 98114 701593
rect 97494 701273 97526 701509
rect 97762 701273 97846 701509
rect 98082 701273 98114 701509
rect 97494 674829 98114 701273
rect 97494 674593 97526 674829
rect 97762 674593 97846 674829
rect 98082 674593 98114 674829
rect 97494 674509 98114 674593
rect 97494 674273 97526 674509
rect 97762 674273 97846 674509
rect 98082 674273 98114 674509
rect 97494 647829 98114 674273
rect 97494 647593 97526 647829
rect 97762 647593 97846 647829
rect 98082 647593 98114 647829
rect 97494 647509 98114 647593
rect 97494 647273 97526 647509
rect 97762 647273 97846 647509
rect 98082 647273 98114 647509
rect 97494 620829 98114 647273
rect 97494 620593 97526 620829
rect 97762 620593 97846 620829
rect 98082 620593 98114 620829
rect 97494 620509 98114 620593
rect 97494 620273 97526 620509
rect 97762 620273 97846 620509
rect 98082 620273 98114 620509
rect 97494 593829 98114 620273
rect 97494 593593 97526 593829
rect 97762 593593 97846 593829
rect 98082 593593 98114 593829
rect 97494 593509 98114 593593
rect 97494 593273 97526 593509
rect 97762 593273 97846 593509
rect 98082 593273 98114 593509
rect 97494 566829 98114 593273
rect 97494 566593 97526 566829
rect 97762 566593 97846 566829
rect 98082 566593 98114 566829
rect 97494 566509 98114 566593
rect 97494 566273 97526 566509
rect 97762 566273 97846 566509
rect 98082 566273 98114 566509
rect 97494 539829 98114 566273
rect 97494 539593 97526 539829
rect 97762 539593 97846 539829
rect 98082 539593 98114 539829
rect 97494 539509 98114 539593
rect 97494 539273 97526 539509
rect 97762 539273 97846 539509
rect 98082 539273 98114 539509
rect 97494 512829 98114 539273
rect 97494 512593 97526 512829
rect 97762 512593 97846 512829
rect 98082 512593 98114 512829
rect 97494 512509 98114 512593
rect 97494 512273 97526 512509
rect 97762 512273 97846 512509
rect 98082 512273 98114 512509
rect 97494 485829 98114 512273
rect 97494 485593 97526 485829
rect 97762 485593 97846 485829
rect 98082 485593 98114 485829
rect 97494 485509 98114 485593
rect 97494 485273 97526 485509
rect 97762 485273 97846 485509
rect 98082 485273 98114 485509
rect 97494 458829 98114 485273
rect 97494 458593 97526 458829
rect 97762 458593 97846 458829
rect 98082 458593 98114 458829
rect 97494 458509 98114 458593
rect 97494 458273 97526 458509
rect 97762 458273 97846 458509
rect 98082 458273 98114 458509
rect 97494 431829 98114 458273
rect 97494 431593 97526 431829
rect 97762 431593 97846 431829
rect 98082 431593 98114 431829
rect 97494 431509 98114 431593
rect 97494 431273 97526 431509
rect 97762 431273 97846 431509
rect 98082 431273 98114 431509
rect 97494 404829 98114 431273
rect 97494 404593 97526 404829
rect 97762 404593 97846 404829
rect 98082 404593 98114 404829
rect 97494 404509 98114 404593
rect 97494 404273 97526 404509
rect 97762 404273 97846 404509
rect 98082 404273 98114 404509
rect 97494 377829 98114 404273
rect 97494 377593 97526 377829
rect 97762 377593 97846 377829
rect 98082 377593 98114 377829
rect 97494 377509 98114 377593
rect 97494 377273 97526 377509
rect 97762 377273 97846 377509
rect 98082 377273 98114 377509
rect 97494 350829 98114 377273
rect 97494 350593 97526 350829
rect 97762 350593 97846 350829
rect 98082 350593 98114 350829
rect 97494 350509 98114 350593
rect 97494 350273 97526 350509
rect 97762 350273 97846 350509
rect 98082 350273 98114 350509
rect 97494 323829 98114 350273
rect 97494 323593 97526 323829
rect 97762 323593 97846 323829
rect 98082 323593 98114 323829
rect 97494 323509 98114 323593
rect 97494 323273 97526 323509
rect 97762 323273 97846 323509
rect 98082 323273 98114 323509
rect 97494 296829 98114 323273
rect 97494 296593 97526 296829
rect 97762 296593 97846 296829
rect 98082 296593 98114 296829
rect 97494 296509 98114 296593
rect 97494 296273 97526 296509
rect 97762 296273 97846 296509
rect 98082 296273 98114 296509
rect 97494 269829 98114 296273
rect 97494 269593 97526 269829
rect 97762 269593 97846 269829
rect 98082 269593 98114 269829
rect 97494 269509 98114 269593
rect 97494 269273 97526 269509
rect 97762 269273 97846 269509
rect 98082 269273 98114 269509
rect 97494 242829 98114 269273
rect 97494 242593 97526 242829
rect 97762 242593 97846 242829
rect 98082 242593 98114 242829
rect 97494 242509 98114 242593
rect 97494 242273 97526 242509
rect 97762 242273 97846 242509
rect 98082 242273 98114 242509
rect 97494 215829 98114 242273
rect 97494 215593 97526 215829
rect 97762 215593 97846 215829
rect 98082 215593 98114 215829
rect 97494 215509 98114 215593
rect 97494 215273 97526 215509
rect 97762 215273 97846 215509
rect 98082 215273 98114 215509
rect 97494 188829 98114 215273
rect 97494 188593 97526 188829
rect 97762 188593 97846 188829
rect 98082 188593 98114 188829
rect 97494 188509 98114 188593
rect 97494 188273 97526 188509
rect 97762 188273 97846 188509
rect 98082 188273 98114 188509
rect 97494 161829 98114 188273
rect 97494 161593 97526 161829
rect 97762 161593 97846 161829
rect 98082 161593 98114 161829
rect 97494 161509 98114 161593
rect 97494 161273 97526 161509
rect 97762 161273 97846 161509
rect 98082 161273 98114 161509
rect 97494 134829 98114 161273
rect 97494 134593 97526 134829
rect 97762 134593 97846 134829
rect 98082 134593 98114 134829
rect 97494 134509 98114 134593
rect 97494 134273 97526 134509
rect 97762 134273 97846 134509
rect 98082 134273 98114 134509
rect 97494 107829 98114 134273
rect 97494 107593 97526 107829
rect 97762 107593 97846 107829
rect 98082 107593 98114 107829
rect 97494 107509 98114 107593
rect 97494 107273 97526 107509
rect 97762 107273 97846 107509
rect 98082 107273 98114 107509
rect 97494 80829 98114 107273
rect 97494 80593 97526 80829
rect 97762 80593 97846 80829
rect 98082 80593 98114 80829
rect 97494 80509 98114 80593
rect 97494 80273 97526 80509
rect 97762 80273 97846 80509
rect 98082 80273 98114 80509
rect 97494 53829 98114 80273
rect 97494 53593 97526 53829
rect 97762 53593 97846 53829
rect 98082 53593 98114 53829
rect 97494 53509 98114 53593
rect 97494 53273 97526 53509
rect 97762 53273 97846 53509
rect 98082 53273 98114 53509
rect 97494 42000 98114 53273
rect 121994 705798 122614 711590
rect 121994 705562 122026 705798
rect 122262 705562 122346 705798
rect 122582 705562 122614 705798
rect 121994 705478 122614 705562
rect 121994 705242 122026 705478
rect 122262 705242 122346 705478
rect 122582 705242 122614 705478
rect 121994 698454 122614 705242
rect 121994 698218 122026 698454
rect 122262 698218 122346 698454
rect 122582 698218 122614 698454
rect 121994 698134 122614 698218
rect 121994 697898 122026 698134
rect 122262 697898 122346 698134
rect 122582 697898 122614 698134
rect 121994 671454 122614 697898
rect 121994 671218 122026 671454
rect 122262 671218 122346 671454
rect 122582 671218 122614 671454
rect 121994 671134 122614 671218
rect 121994 670898 122026 671134
rect 122262 670898 122346 671134
rect 122582 670898 122614 671134
rect 121994 644454 122614 670898
rect 121994 644218 122026 644454
rect 122262 644218 122346 644454
rect 122582 644218 122614 644454
rect 121994 644134 122614 644218
rect 121994 643898 122026 644134
rect 122262 643898 122346 644134
rect 122582 643898 122614 644134
rect 121994 617454 122614 643898
rect 121994 617218 122026 617454
rect 122262 617218 122346 617454
rect 122582 617218 122614 617454
rect 121994 617134 122614 617218
rect 121994 616898 122026 617134
rect 122262 616898 122346 617134
rect 122582 616898 122614 617134
rect 121994 590454 122614 616898
rect 121994 590218 122026 590454
rect 122262 590218 122346 590454
rect 122582 590218 122614 590454
rect 121994 590134 122614 590218
rect 121994 589898 122026 590134
rect 122262 589898 122346 590134
rect 122582 589898 122614 590134
rect 121994 563454 122614 589898
rect 121994 563218 122026 563454
rect 122262 563218 122346 563454
rect 122582 563218 122614 563454
rect 121994 563134 122614 563218
rect 121994 562898 122026 563134
rect 122262 562898 122346 563134
rect 122582 562898 122614 563134
rect 121994 536454 122614 562898
rect 121994 536218 122026 536454
rect 122262 536218 122346 536454
rect 122582 536218 122614 536454
rect 121994 536134 122614 536218
rect 121994 535898 122026 536134
rect 122262 535898 122346 536134
rect 122582 535898 122614 536134
rect 121994 509454 122614 535898
rect 121994 509218 122026 509454
rect 122262 509218 122346 509454
rect 122582 509218 122614 509454
rect 121994 509134 122614 509218
rect 121994 508898 122026 509134
rect 122262 508898 122346 509134
rect 122582 508898 122614 509134
rect 121994 482454 122614 508898
rect 121994 482218 122026 482454
rect 122262 482218 122346 482454
rect 122582 482218 122614 482454
rect 121994 482134 122614 482218
rect 121994 481898 122026 482134
rect 122262 481898 122346 482134
rect 122582 481898 122614 482134
rect 121994 455454 122614 481898
rect 121994 455218 122026 455454
rect 122262 455218 122346 455454
rect 122582 455218 122614 455454
rect 121994 455134 122614 455218
rect 121994 454898 122026 455134
rect 122262 454898 122346 455134
rect 122582 454898 122614 455134
rect 121994 428454 122614 454898
rect 121994 428218 122026 428454
rect 122262 428218 122346 428454
rect 122582 428218 122614 428454
rect 121994 428134 122614 428218
rect 121994 427898 122026 428134
rect 122262 427898 122346 428134
rect 122582 427898 122614 428134
rect 121994 401454 122614 427898
rect 121994 401218 122026 401454
rect 122262 401218 122346 401454
rect 122582 401218 122614 401454
rect 121994 401134 122614 401218
rect 121994 400898 122026 401134
rect 122262 400898 122346 401134
rect 122582 400898 122614 401134
rect 121994 374454 122614 400898
rect 121994 374218 122026 374454
rect 122262 374218 122346 374454
rect 122582 374218 122614 374454
rect 121994 374134 122614 374218
rect 121994 373898 122026 374134
rect 122262 373898 122346 374134
rect 122582 373898 122614 374134
rect 121994 347454 122614 373898
rect 121994 347218 122026 347454
rect 122262 347218 122346 347454
rect 122582 347218 122614 347454
rect 121994 347134 122614 347218
rect 121994 346898 122026 347134
rect 122262 346898 122346 347134
rect 122582 346898 122614 347134
rect 121994 320454 122614 346898
rect 121994 320218 122026 320454
rect 122262 320218 122346 320454
rect 122582 320218 122614 320454
rect 121994 320134 122614 320218
rect 121994 319898 122026 320134
rect 122262 319898 122346 320134
rect 122582 319898 122614 320134
rect 121994 293454 122614 319898
rect 121994 293218 122026 293454
rect 122262 293218 122346 293454
rect 122582 293218 122614 293454
rect 121994 293134 122614 293218
rect 121994 292898 122026 293134
rect 122262 292898 122346 293134
rect 122582 292898 122614 293134
rect 121994 266454 122614 292898
rect 121994 266218 122026 266454
rect 122262 266218 122346 266454
rect 122582 266218 122614 266454
rect 121994 266134 122614 266218
rect 121994 265898 122026 266134
rect 122262 265898 122346 266134
rect 122582 265898 122614 266134
rect 121994 239454 122614 265898
rect 121994 239218 122026 239454
rect 122262 239218 122346 239454
rect 122582 239218 122614 239454
rect 121994 239134 122614 239218
rect 121994 238898 122026 239134
rect 122262 238898 122346 239134
rect 122582 238898 122614 239134
rect 121994 212454 122614 238898
rect 121994 212218 122026 212454
rect 122262 212218 122346 212454
rect 122582 212218 122614 212454
rect 121994 212134 122614 212218
rect 121994 211898 122026 212134
rect 122262 211898 122346 212134
rect 122582 211898 122614 212134
rect 121994 185454 122614 211898
rect 121994 185218 122026 185454
rect 122262 185218 122346 185454
rect 122582 185218 122614 185454
rect 121994 185134 122614 185218
rect 121994 184898 122026 185134
rect 122262 184898 122346 185134
rect 122582 184898 122614 185134
rect 121994 158454 122614 184898
rect 121994 158218 122026 158454
rect 122262 158218 122346 158454
rect 122582 158218 122614 158454
rect 121994 158134 122614 158218
rect 121994 157898 122026 158134
rect 122262 157898 122346 158134
rect 122582 157898 122614 158134
rect 121994 131454 122614 157898
rect 121994 131218 122026 131454
rect 122262 131218 122346 131454
rect 122582 131218 122614 131454
rect 121994 131134 122614 131218
rect 121994 130898 122026 131134
rect 122262 130898 122346 131134
rect 122582 130898 122614 131134
rect 121994 104454 122614 130898
rect 121994 104218 122026 104454
rect 122262 104218 122346 104454
rect 122582 104218 122614 104454
rect 121994 104134 122614 104218
rect 121994 103898 122026 104134
rect 122262 103898 122346 104134
rect 122582 103898 122614 104134
rect 121994 77454 122614 103898
rect 121994 77218 122026 77454
rect 122262 77218 122346 77454
rect 122582 77218 122614 77454
rect 121994 77134 122614 77218
rect 121994 76898 122026 77134
rect 122262 76898 122346 77134
rect 122582 76898 122614 77134
rect 121994 50454 122614 76898
rect 121994 50218 122026 50454
rect 122262 50218 122346 50454
rect 122582 50218 122614 50454
rect 121994 50134 122614 50218
rect 121994 49898 122026 50134
rect 122262 49898 122346 50134
rect 122582 49898 122614 50134
rect 121994 42000 122614 49898
rect 125494 704838 126114 711590
rect 125494 704602 125526 704838
rect 125762 704602 125846 704838
rect 126082 704602 126114 704838
rect 125494 704518 126114 704602
rect 125494 704282 125526 704518
rect 125762 704282 125846 704518
rect 126082 704282 126114 704518
rect 125494 701829 126114 704282
rect 125494 701593 125526 701829
rect 125762 701593 125846 701829
rect 126082 701593 126114 701829
rect 125494 701509 126114 701593
rect 125494 701273 125526 701509
rect 125762 701273 125846 701509
rect 126082 701273 126114 701509
rect 125494 674829 126114 701273
rect 125494 674593 125526 674829
rect 125762 674593 125846 674829
rect 126082 674593 126114 674829
rect 125494 674509 126114 674593
rect 125494 674273 125526 674509
rect 125762 674273 125846 674509
rect 126082 674273 126114 674509
rect 125494 647829 126114 674273
rect 125494 647593 125526 647829
rect 125762 647593 125846 647829
rect 126082 647593 126114 647829
rect 125494 647509 126114 647593
rect 125494 647273 125526 647509
rect 125762 647273 125846 647509
rect 126082 647273 126114 647509
rect 125494 620829 126114 647273
rect 125494 620593 125526 620829
rect 125762 620593 125846 620829
rect 126082 620593 126114 620829
rect 125494 620509 126114 620593
rect 125494 620273 125526 620509
rect 125762 620273 125846 620509
rect 126082 620273 126114 620509
rect 125494 593829 126114 620273
rect 125494 593593 125526 593829
rect 125762 593593 125846 593829
rect 126082 593593 126114 593829
rect 125494 593509 126114 593593
rect 125494 593273 125526 593509
rect 125762 593273 125846 593509
rect 126082 593273 126114 593509
rect 125494 566829 126114 593273
rect 125494 566593 125526 566829
rect 125762 566593 125846 566829
rect 126082 566593 126114 566829
rect 125494 566509 126114 566593
rect 125494 566273 125526 566509
rect 125762 566273 125846 566509
rect 126082 566273 126114 566509
rect 125494 539829 126114 566273
rect 125494 539593 125526 539829
rect 125762 539593 125846 539829
rect 126082 539593 126114 539829
rect 125494 539509 126114 539593
rect 125494 539273 125526 539509
rect 125762 539273 125846 539509
rect 126082 539273 126114 539509
rect 125494 512829 126114 539273
rect 125494 512593 125526 512829
rect 125762 512593 125846 512829
rect 126082 512593 126114 512829
rect 125494 512509 126114 512593
rect 125494 512273 125526 512509
rect 125762 512273 125846 512509
rect 126082 512273 126114 512509
rect 125494 485829 126114 512273
rect 125494 485593 125526 485829
rect 125762 485593 125846 485829
rect 126082 485593 126114 485829
rect 125494 485509 126114 485593
rect 125494 485273 125526 485509
rect 125762 485273 125846 485509
rect 126082 485273 126114 485509
rect 125494 458829 126114 485273
rect 125494 458593 125526 458829
rect 125762 458593 125846 458829
rect 126082 458593 126114 458829
rect 125494 458509 126114 458593
rect 125494 458273 125526 458509
rect 125762 458273 125846 458509
rect 126082 458273 126114 458509
rect 125494 431829 126114 458273
rect 125494 431593 125526 431829
rect 125762 431593 125846 431829
rect 126082 431593 126114 431829
rect 125494 431509 126114 431593
rect 125494 431273 125526 431509
rect 125762 431273 125846 431509
rect 126082 431273 126114 431509
rect 125494 404829 126114 431273
rect 125494 404593 125526 404829
rect 125762 404593 125846 404829
rect 126082 404593 126114 404829
rect 125494 404509 126114 404593
rect 125494 404273 125526 404509
rect 125762 404273 125846 404509
rect 126082 404273 126114 404509
rect 125494 377829 126114 404273
rect 125494 377593 125526 377829
rect 125762 377593 125846 377829
rect 126082 377593 126114 377829
rect 125494 377509 126114 377593
rect 125494 377273 125526 377509
rect 125762 377273 125846 377509
rect 126082 377273 126114 377509
rect 125494 350829 126114 377273
rect 125494 350593 125526 350829
rect 125762 350593 125846 350829
rect 126082 350593 126114 350829
rect 125494 350509 126114 350593
rect 125494 350273 125526 350509
rect 125762 350273 125846 350509
rect 126082 350273 126114 350509
rect 125494 323829 126114 350273
rect 125494 323593 125526 323829
rect 125762 323593 125846 323829
rect 126082 323593 126114 323829
rect 125494 323509 126114 323593
rect 125494 323273 125526 323509
rect 125762 323273 125846 323509
rect 126082 323273 126114 323509
rect 125494 296829 126114 323273
rect 125494 296593 125526 296829
rect 125762 296593 125846 296829
rect 126082 296593 126114 296829
rect 125494 296509 126114 296593
rect 125494 296273 125526 296509
rect 125762 296273 125846 296509
rect 126082 296273 126114 296509
rect 125494 269829 126114 296273
rect 125494 269593 125526 269829
rect 125762 269593 125846 269829
rect 126082 269593 126114 269829
rect 125494 269509 126114 269593
rect 125494 269273 125526 269509
rect 125762 269273 125846 269509
rect 126082 269273 126114 269509
rect 125494 242829 126114 269273
rect 125494 242593 125526 242829
rect 125762 242593 125846 242829
rect 126082 242593 126114 242829
rect 125494 242509 126114 242593
rect 125494 242273 125526 242509
rect 125762 242273 125846 242509
rect 126082 242273 126114 242509
rect 125494 215829 126114 242273
rect 125494 215593 125526 215829
rect 125762 215593 125846 215829
rect 126082 215593 126114 215829
rect 125494 215509 126114 215593
rect 125494 215273 125526 215509
rect 125762 215273 125846 215509
rect 126082 215273 126114 215509
rect 125494 188829 126114 215273
rect 125494 188593 125526 188829
rect 125762 188593 125846 188829
rect 126082 188593 126114 188829
rect 125494 188509 126114 188593
rect 125494 188273 125526 188509
rect 125762 188273 125846 188509
rect 126082 188273 126114 188509
rect 125494 161829 126114 188273
rect 125494 161593 125526 161829
rect 125762 161593 125846 161829
rect 126082 161593 126114 161829
rect 125494 161509 126114 161593
rect 125494 161273 125526 161509
rect 125762 161273 125846 161509
rect 126082 161273 126114 161509
rect 125494 134829 126114 161273
rect 125494 134593 125526 134829
rect 125762 134593 125846 134829
rect 126082 134593 126114 134829
rect 125494 134509 126114 134593
rect 125494 134273 125526 134509
rect 125762 134273 125846 134509
rect 126082 134273 126114 134509
rect 125494 107829 126114 134273
rect 125494 107593 125526 107829
rect 125762 107593 125846 107829
rect 126082 107593 126114 107829
rect 125494 107509 126114 107593
rect 125494 107273 125526 107509
rect 125762 107273 125846 107509
rect 126082 107273 126114 107509
rect 125494 80829 126114 107273
rect 125494 80593 125526 80829
rect 125762 80593 125846 80829
rect 126082 80593 126114 80829
rect 125494 80509 126114 80593
rect 125494 80273 125526 80509
rect 125762 80273 125846 80509
rect 126082 80273 126114 80509
rect 125494 53829 126114 80273
rect 125494 53593 125526 53829
rect 125762 53593 125846 53829
rect 126082 53593 126114 53829
rect 125494 53509 126114 53593
rect 125494 53273 125526 53509
rect 125762 53273 125846 53509
rect 126082 53273 126114 53509
rect 125494 42000 126114 53273
rect 149994 705798 150614 711590
rect 149994 705562 150026 705798
rect 150262 705562 150346 705798
rect 150582 705562 150614 705798
rect 149994 705478 150614 705562
rect 149994 705242 150026 705478
rect 150262 705242 150346 705478
rect 150582 705242 150614 705478
rect 149994 698454 150614 705242
rect 149994 698218 150026 698454
rect 150262 698218 150346 698454
rect 150582 698218 150614 698454
rect 149994 698134 150614 698218
rect 149994 697898 150026 698134
rect 150262 697898 150346 698134
rect 150582 697898 150614 698134
rect 149994 671454 150614 697898
rect 149994 671218 150026 671454
rect 150262 671218 150346 671454
rect 150582 671218 150614 671454
rect 149994 671134 150614 671218
rect 149994 670898 150026 671134
rect 150262 670898 150346 671134
rect 150582 670898 150614 671134
rect 149994 644454 150614 670898
rect 149994 644218 150026 644454
rect 150262 644218 150346 644454
rect 150582 644218 150614 644454
rect 149994 644134 150614 644218
rect 149994 643898 150026 644134
rect 150262 643898 150346 644134
rect 150582 643898 150614 644134
rect 149994 617454 150614 643898
rect 149994 617218 150026 617454
rect 150262 617218 150346 617454
rect 150582 617218 150614 617454
rect 149994 617134 150614 617218
rect 149994 616898 150026 617134
rect 150262 616898 150346 617134
rect 150582 616898 150614 617134
rect 149994 590454 150614 616898
rect 149994 590218 150026 590454
rect 150262 590218 150346 590454
rect 150582 590218 150614 590454
rect 149994 590134 150614 590218
rect 149994 589898 150026 590134
rect 150262 589898 150346 590134
rect 150582 589898 150614 590134
rect 149994 563454 150614 589898
rect 149994 563218 150026 563454
rect 150262 563218 150346 563454
rect 150582 563218 150614 563454
rect 149994 563134 150614 563218
rect 149994 562898 150026 563134
rect 150262 562898 150346 563134
rect 150582 562898 150614 563134
rect 149994 536454 150614 562898
rect 149994 536218 150026 536454
rect 150262 536218 150346 536454
rect 150582 536218 150614 536454
rect 149994 536134 150614 536218
rect 149994 535898 150026 536134
rect 150262 535898 150346 536134
rect 150582 535898 150614 536134
rect 149994 509454 150614 535898
rect 149994 509218 150026 509454
rect 150262 509218 150346 509454
rect 150582 509218 150614 509454
rect 149994 509134 150614 509218
rect 149994 508898 150026 509134
rect 150262 508898 150346 509134
rect 150582 508898 150614 509134
rect 149994 482454 150614 508898
rect 149994 482218 150026 482454
rect 150262 482218 150346 482454
rect 150582 482218 150614 482454
rect 149994 482134 150614 482218
rect 149994 481898 150026 482134
rect 150262 481898 150346 482134
rect 150582 481898 150614 482134
rect 149994 455454 150614 481898
rect 149994 455218 150026 455454
rect 150262 455218 150346 455454
rect 150582 455218 150614 455454
rect 149994 455134 150614 455218
rect 149994 454898 150026 455134
rect 150262 454898 150346 455134
rect 150582 454898 150614 455134
rect 149994 428454 150614 454898
rect 149994 428218 150026 428454
rect 150262 428218 150346 428454
rect 150582 428218 150614 428454
rect 149994 428134 150614 428218
rect 149994 427898 150026 428134
rect 150262 427898 150346 428134
rect 150582 427898 150614 428134
rect 149994 401454 150614 427898
rect 149994 401218 150026 401454
rect 150262 401218 150346 401454
rect 150582 401218 150614 401454
rect 149994 401134 150614 401218
rect 149994 400898 150026 401134
rect 150262 400898 150346 401134
rect 150582 400898 150614 401134
rect 149994 374454 150614 400898
rect 149994 374218 150026 374454
rect 150262 374218 150346 374454
rect 150582 374218 150614 374454
rect 149994 374134 150614 374218
rect 149994 373898 150026 374134
rect 150262 373898 150346 374134
rect 150582 373898 150614 374134
rect 149994 347454 150614 373898
rect 149994 347218 150026 347454
rect 150262 347218 150346 347454
rect 150582 347218 150614 347454
rect 149994 347134 150614 347218
rect 149994 346898 150026 347134
rect 150262 346898 150346 347134
rect 150582 346898 150614 347134
rect 149994 320454 150614 346898
rect 149994 320218 150026 320454
rect 150262 320218 150346 320454
rect 150582 320218 150614 320454
rect 149994 320134 150614 320218
rect 149994 319898 150026 320134
rect 150262 319898 150346 320134
rect 150582 319898 150614 320134
rect 149994 293454 150614 319898
rect 149994 293218 150026 293454
rect 150262 293218 150346 293454
rect 150582 293218 150614 293454
rect 149994 293134 150614 293218
rect 149994 292898 150026 293134
rect 150262 292898 150346 293134
rect 150582 292898 150614 293134
rect 149994 266454 150614 292898
rect 149994 266218 150026 266454
rect 150262 266218 150346 266454
rect 150582 266218 150614 266454
rect 149994 266134 150614 266218
rect 149994 265898 150026 266134
rect 150262 265898 150346 266134
rect 150582 265898 150614 266134
rect 149994 239454 150614 265898
rect 149994 239218 150026 239454
rect 150262 239218 150346 239454
rect 150582 239218 150614 239454
rect 149994 239134 150614 239218
rect 149994 238898 150026 239134
rect 150262 238898 150346 239134
rect 150582 238898 150614 239134
rect 149994 212454 150614 238898
rect 149994 212218 150026 212454
rect 150262 212218 150346 212454
rect 150582 212218 150614 212454
rect 149994 212134 150614 212218
rect 149994 211898 150026 212134
rect 150262 211898 150346 212134
rect 150582 211898 150614 212134
rect 149994 185454 150614 211898
rect 149994 185218 150026 185454
rect 150262 185218 150346 185454
rect 150582 185218 150614 185454
rect 149994 185134 150614 185218
rect 149994 184898 150026 185134
rect 150262 184898 150346 185134
rect 150582 184898 150614 185134
rect 149994 158454 150614 184898
rect 149994 158218 150026 158454
rect 150262 158218 150346 158454
rect 150582 158218 150614 158454
rect 149994 158134 150614 158218
rect 149994 157898 150026 158134
rect 150262 157898 150346 158134
rect 150582 157898 150614 158134
rect 149994 131454 150614 157898
rect 149994 131218 150026 131454
rect 150262 131218 150346 131454
rect 150582 131218 150614 131454
rect 149994 131134 150614 131218
rect 149994 130898 150026 131134
rect 150262 130898 150346 131134
rect 150582 130898 150614 131134
rect 149994 104454 150614 130898
rect 149994 104218 150026 104454
rect 150262 104218 150346 104454
rect 150582 104218 150614 104454
rect 149994 104134 150614 104218
rect 149994 103898 150026 104134
rect 150262 103898 150346 104134
rect 150582 103898 150614 104134
rect 149994 77454 150614 103898
rect 149994 77218 150026 77454
rect 150262 77218 150346 77454
rect 150582 77218 150614 77454
rect 149994 77134 150614 77218
rect 149994 76898 150026 77134
rect 150262 76898 150346 77134
rect 150582 76898 150614 77134
rect 149994 50454 150614 76898
rect 149994 50218 150026 50454
rect 150262 50218 150346 50454
rect 150582 50218 150614 50454
rect 149994 50134 150614 50218
rect 149994 49898 150026 50134
rect 150262 49898 150346 50134
rect 150582 49898 150614 50134
rect 149994 42000 150614 49898
rect 153494 704838 154114 711590
rect 153494 704602 153526 704838
rect 153762 704602 153846 704838
rect 154082 704602 154114 704838
rect 153494 704518 154114 704602
rect 153494 704282 153526 704518
rect 153762 704282 153846 704518
rect 154082 704282 154114 704518
rect 153494 701829 154114 704282
rect 153494 701593 153526 701829
rect 153762 701593 153846 701829
rect 154082 701593 154114 701829
rect 153494 701509 154114 701593
rect 153494 701273 153526 701509
rect 153762 701273 153846 701509
rect 154082 701273 154114 701509
rect 153494 674829 154114 701273
rect 177994 705798 178614 711590
rect 177994 705562 178026 705798
rect 178262 705562 178346 705798
rect 178582 705562 178614 705798
rect 177994 705478 178614 705562
rect 177994 705242 178026 705478
rect 178262 705242 178346 705478
rect 178582 705242 178614 705478
rect 169707 699820 169773 699821
rect 169707 699756 169708 699820
rect 169772 699756 169773 699820
rect 169707 699755 169773 699756
rect 153494 674593 153526 674829
rect 153762 674593 153846 674829
rect 154082 674593 154114 674829
rect 153494 674509 154114 674593
rect 153494 674273 153526 674509
rect 153762 674273 153846 674509
rect 154082 674273 154114 674509
rect 153494 647829 154114 674273
rect 153494 647593 153526 647829
rect 153762 647593 153846 647829
rect 154082 647593 154114 647829
rect 153494 647509 154114 647593
rect 153494 647273 153526 647509
rect 153762 647273 153846 647509
rect 154082 647273 154114 647509
rect 153494 620829 154114 647273
rect 153494 620593 153526 620829
rect 153762 620593 153846 620829
rect 154082 620593 154114 620829
rect 153494 620509 154114 620593
rect 153494 620273 153526 620509
rect 153762 620273 153846 620509
rect 154082 620273 154114 620509
rect 153494 593829 154114 620273
rect 153494 593593 153526 593829
rect 153762 593593 153846 593829
rect 154082 593593 154114 593829
rect 153494 593509 154114 593593
rect 153494 593273 153526 593509
rect 153762 593273 153846 593509
rect 154082 593273 154114 593509
rect 153494 566829 154114 593273
rect 153494 566593 153526 566829
rect 153762 566593 153846 566829
rect 154082 566593 154114 566829
rect 153494 566509 154114 566593
rect 153494 566273 153526 566509
rect 153762 566273 153846 566509
rect 154082 566273 154114 566509
rect 153494 539829 154114 566273
rect 153494 539593 153526 539829
rect 153762 539593 153846 539829
rect 154082 539593 154114 539829
rect 153494 539509 154114 539593
rect 153494 539273 153526 539509
rect 153762 539273 153846 539509
rect 154082 539273 154114 539509
rect 153494 512829 154114 539273
rect 153494 512593 153526 512829
rect 153762 512593 153846 512829
rect 154082 512593 154114 512829
rect 153494 512509 154114 512593
rect 153494 512273 153526 512509
rect 153762 512273 153846 512509
rect 154082 512273 154114 512509
rect 153494 485829 154114 512273
rect 153494 485593 153526 485829
rect 153762 485593 153846 485829
rect 154082 485593 154114 485829
rect 153494 485509 154114 485593
rect 153494 485273 153526 485509
rect 153762 485273 153846 485509
rect 154082 485273 154114 485509
rect 153494 458829 154114 485273
rect 153494 458593 153526 458829
rect 153762 458593 153846 458829
rect 154082 458593 154114 458829
rect 153494 458509 154114 458593
rect 153494 458273 153526 458509
rect 153762 458273 153846 458509
rect 154082 458273 154114 458509
rect 153494 431829 154114 458273
rect 153494 431593 153526 431829
rect 153762 431593 153846 431829
rect 154082 431593 154114 431829
rect 153494 431509 154114 431593
rect 153494 431273 153526 431509
rect 153762 431273 153846 431509
rect 154082 431273 154114 431509
rect 153494 404829 154114 431273
rect 153494 404593 153526 404829
rect 153762 404593 153846 404829
rect 154082 404593 154114 404829
rect 153494 404509 154114 404593
rect 153494 404273 153526 404509
rect 153762 404273 153846 404509
rect 154082 404273 154114 404509
rect 153494 377829 154114 404273
rect 153494 377593 153526 377829
rect 153762 377593 153846 377829
rect 154082 377593 154114 377829
rect 153494 377509 154114 377593
rect 153494 377273 153526 377509
rect 153762 377273 153846 377509
rect 154082 377273 154114 377509
rect 153494 350829 154114 377273
rect 153494 350593 153526 350829
rect 153762 350593 153846 350829
rect 154082 350593 154114 350829
rect 153494 350509 154114 350593
rect 153494 350273 153526 350509
rect 153762 350273 153846 350509
rect 154082 350273 154114 350509
rect 153494 323829 154114 350273
rect 153494 323593 153526 323829
rect 153762 323593 153846 323829
rect 154082 323593 154114 323829
rect 153494 323509 154114 323593
rect 153494 323273 153526 323509
rect 153762 323273 153846 323509
rect 154082 323273 154114 323509
rect 153494 296829 154114 323273
rect 153494 296593 153526 296829
rect 153762 296593 153846 296829
rect 154082 296593 154114 296829
rect 153494 296509 154114 296593
rect 153494 296273 153526 296509
rect 153762 296273 153846 296509
rect 154082 296273 154114 296509
rect 153494 269829 154114 296273
rect 153494 269593 153526 269829
rect 153762 269593 153846 269829
rect 154082 269593 154114 269829
rect 153494 269509 154114 269593
rect 153494 269273 153526 269509
rect 153762 269273 153846 269509
rect 154082 269273 154114 269509
rect 153494 242829 154114 269273
rect 153494 242593 153526 242829
rect 153762 242593 153846 242829
rect 154082 242593 154114 242829
rect 153494 242509 154114 242593
rect 153494 242273 153526 242509
rect 153762 242273 153846 242509
rect 154082 242273 154114 242509
rect 153494 215829 154114 242273
rect 153494 215593 153526 215829
rect 153762 215593 153846 215829
rect 154082 215593 154114 215829
rect 153494 215509 154114 215593
rect 153494 215273 153526 215509
rect 153762 215273 153846 215509
rect 154082 215273 154114 215509
rect 153494 188829 154114 215273
rect 153494 188593 153526 188829
rect 153762 188593 153846 188829
rect 154082 188593 154114 188829
rect 153494 188509 154114 188593
rect 153494 188273 153526 188509
rect 153762 188273 153846 188509
rect 154082 188273 154114 188509
rect 153494 161829 154114 188273
rect 153494 161593 153526 161829
rect 153762 161593 153846 161829
rect 154082 161593 154114 161829
rect 153494 161509 154114 161593
rect 153494 161273 153526 161509
rect 153762 161273 153846 161509
rect 154082 161273 154114 161509
rect 153494 134829 154114 161273
rect 153494 134593 153526 134829
rect 153762 134593 153846 134829
rect 154082 134593 154114 134829
rect 153494 134509 154114 134593
rect 153494 134273 153526 134509
rect 153762 134273 153846 134509
rect 154082 134273 154114 134509
rect 153494 107829 154114 134273
rect 153494 107593 153526 107829
rect 153762 107593 153846 107829
rect 154082 107593 154114 107829
rect 153494 107509 154114 107593
rect 153494 107273 153526 107509
rect 153762 107273 153846 107509
rect 154082 107273 154114 107509
rect 153494 80829 154114 107273
rect 153494 80593 153526 80829
rect 153762 80593 153846 80829
rect 154082 80593 154114 80829
rect 153494 80509 154114 80593
rect 153494 80273 153526 80509
rect 153762 80273 153846 80509
rect 154082 80273 154114 80509
rect 153494 53829 154114 80273
rect 153494 53593 153526 53829
rect 153762 53593 153846 53829
rect 154082 53593 154114 53829
rect 153494 53509 154114 53593
rect 153494 53273 153526 53509
rect 153762 53273 153846 53509
rect 154082 53273 154114 53509
rect 153494 42000 154114 53273
rect 69494 26593 69526 26829
rect 69762 26593 69846 26829
rect 70082 26593 70114 26829
rect 69494 26509 70114 26593
rect 69494 26273 69526 26509
rect 69762 26273 69846 26509
rect 70082 26273 70114 26509
rect 69494 -346 70114 26273
rect 75418 26829 75738 26861
rect 75418 26593 75460 26829
rect 75696 26593 75738 26829
rect 75418 26509 75738 26593
rect 75418 26273 75460 26509
rect 75696 26273 75738 26509
rect 75418 26241 75738 26273
rect 76366 26829 76686 26861
rect 76366 26593 76408 26829
rect 76644 26593 76686 26829
rect 76366 26509 76686 26593
rect 76366 26273 76408 26509
rect 76644 26273 76686 26509
rect 76366 26241 76686 26273
rect 77314 26829 77634 26861
rect 77314 26593 77356 26829
rect 77592 26593 77634 26829
rect 77314 26509 77634 26593
rect 77314 26273 77356 26509
rect 77592 26273 77634 26509
rect 77314 26241 77634 26273
rect 78262 26829 78582 26861
rect 78262 26593 78304 26829
rect 78540 26593 78582 26829
rect 78262 26509 78582 26593
rect 78262 26273 78304 26509
rect 78540 26273 78582 26509
rect 78262 26241 78582 26273
rect 84118 26829 84438 26861
rect 84118 26593 84160 26829
rect 84396 26593 84438 26829
rect 84118 26509 84438 26593
rect 84118 26273 84160 26509
rect 84396 26273 84438 26509
rect 84118 26241 84438 26273
rect 88066 26829 88386 26861
rect 88066 26593 88108 26829
rect 88344 26593 88386 26829
rect 88066 26509 88386 26593
rect 88066 26273 88108 26509
rect 88344 26273 88386 26509
rect 88066 26241 88386 26273
rect 92014 26829 92334 26861
rect 92014 26593 92056 26829
rect 92292 26593 92334 26829
rect 92014 26509 92334 26593
rect 92014 26273 92056 26509
rect 92292 26273 92334 26509
rect 92014 26241 92334 26273
rect 95962 26829 96282 26861
rect 95962 26593 96004 26829
rect 96240 26593 96282 26829
rect 95962 26509 96282 26593
rect 95962 26273 96004 26509
rect 96240 26273 96282 26509
rect 95962 26241 96282 26273
rect 104418 26829 104738 26861
rect 104418 26593 104460 26829
rect 104696 26593 104738 26829
rect 104418 26509 104738 26593
rect 104418 26273 104460 26509
rect 104696 26273 104738 26509
rect 104418 26241 104738 26273
rect 105366 26829 105686 26861
rect 105366 26593 105408 26829
rect 105644 26593 105686 26829
rect 105366 26509 105686 26593
rect 105366 26273 105408 26509
rect 105644 26273 105686 26509
rect 105366 26241 105686 26273
rect 106314 26829 106634 26861
rect 106314 26593 106356 26829
rect 106592 26593 106634 26829
rect 106314 26509 106634 26593
rect 106314 26273 106356 26509
rect 106592 26273 106634 26509
rect 106314 26241 106634 26273
rect 107262 26829 107582 26861
rect 107262 26593 107304 26829
rect 107540 26593 107582 26829
rect 107262 26509 107582 26593
rect 107262 26273 107304 26509
rect 107540 26273 107582 26509
rect 107262 26241 107582 26273
rect 113118 26829 113438 26861
rect 113118 26593 113160 26829
rect 113396 26593 113438 26829
rect 113118 26509 113438 26593
rect 113118 26273 113160 26509
rect 113396 26273 113438 26509
rect 113118 26241 113438 26273
rect 117066 26829 117386 26861
rect 117066 26593 117108 26829
rect 117344 26593 117386 26829
rect 117066 26509 117386 26593
rect 117066 26273 117108 26509
rect 117344 26273 117386 26509
rect 117066 26241 117386 26273
rect 121014 26829 121334 26861
rect 121014 26593 121056 26829
rect 121292 26593 121334 26829
rect 121014 26509 121334 26593
rect 121014 26273 121056 26509
rect 121292 26273 121334 26509
rect 121014 26241 121334 26273
rect 124962 26829 125282 26861
rect 124962 26593 125004 26829
rect 125240 26593 125282 26829
rect 124962 26509 125282 26593
rect 124962 26273 125004 26509
rect 125240 26273 125282 26509
rect 124962 26241 125282 26273
rect 133418 26829 133738 26861
rect 133418 26593 133460 26829
rect 133696 26593 133738 26829
rect 133418 26509 133738 26593
rect 133418 26273 133460 26509
rect 133696 26273 133738 26509
rect 133418 26241 133738 26273
rect 134366 26829 134686 26861
rect 134366 26593 134408 26829
rect 134644 26593 134686 26829
rect 134366 26509 134686 26593
rect 134366 26273 134408 26509
rect 134644 26273 134686 26509
rect 134366 26241 134686 26273
rect 135314 26829 135634 26861
rect 135314 26593 135356 26829
rect 135592 26593 135634 26829
rect 135314 26509 135634 26593
rect 135314 26273 135356 26509
rect 135592 26273 135634 26509
rect 135314 26241 135634 26273
rect 136262 26829 136582 26861
rect 136262 26593 136304 26829
rect 136540 26593 136582 26829
rect 136262 26509 136582 26593
rect 136262 26273 136304 26509
rect 136540 26273 136582 26509
rect 136262 26241 136582 26273
rect 142118 26829 142438 26861
rect 142118 26593 142160 26829
rect 142396 26593 142438 26829
rect 142118 26509 142438 26593
rect 142118 26273 142160 26509
rect 142396 26273 142438 26509
rect 142118 26241 142438 26273
rect 146066 26829 146386 26861
rect 146066 26593 146108 26829
rect 146344 26593 146386 26829
rect 146066 26509 146386 26593
rect 146066 26273 146108 26509
rect 146344 26273 146386 26509
rect 146066 26241 146386 26273
rect 150014 26829 150334 26861
rect 150014 26593 150056 26829
rect 150292 26593 150334 26829
rect 150014 26509 150334 26593
rect 150014 26273 150056 26509
rect 150292 26273 150334 26509
rect 150014 26241 150334 26273
rect 153962 26829 154282 26861
rect 153962 26593 154004 26829
rect 154240 26593 154282 26829
rect 153962 26509 154282 26593
rect 153962 26273 154004 26509
rect 154240 26273 154282 26509
rect 153962 26241 154282 26273
rect 162418 26829 162738 26861
rect 162418 26593 162460 26829
rect 162696 26593 162738 26829
rect 162418 26509 162738 26593
rect 162418 26273 162460 26509
rect 162696 26273 162738 26509
rect 162418 26241 162738 26273
rect 163366 26829 163686 26861
rect 163366 26593 163408 26829
rect 163644 26593 163686 26829
rect 163366 26509 163686 26593
rect 163366 26273 163408 26509
rect 163644 26273 163686 26509
rect 163366 26241 163686 26273
rect 164314 26829 164634 26861
rect 164314 26593 164356 26829
rect 164592 26593 164634 26829
rect 164314 26509 164634 26593
rect 164314 26273 164356 26509
rect 164592 26273 164634 26509
rect 164314 26241 164634 26273
rect 165262 26829 165582 26861
rect 165262 26593 165304 26829
rect 165540 26593 165582 26829
rect 165262 26509 165582 26593
rect 165262 26273 165304 26509
rect 165540 26273 165582 26509
rect 165262 26241 165582 26273
rect 75892 23454 76212 23486
rect 75892 23218 75934 23454
rect 76170 23218 76212 23454
rect 75892 23134 76212 23218
rect 75892 22898 75934 23134
rect 76170 22898 76212 23134
rect 75892 22866 76212 22898
rect 76840 23454 77160 23486
rect 76840 23218 76882 23454
rect 77118 23218 77160 23454
rect 76840 23134 77160 23218
rect 76840 22898 76882 23134
rect 77118 22898 77160 23134
rect 76840 22866 77160 22898
rect 77788 23454 78108 23486
rect 77788 23218 77830 23454
rect 78066 23218 78108 23454
rect 77788 23134 78108 23218
rect 77788 22898 77830 23134
rect 78066 22898 78108 23134
rect 77788 22866 78108 22898
rect 86092 23454 86412 23486
rect 86092 23218 86134 23454
rect 86370 23218 86412 23454
rect 86092 23134 86412 23218
rect 86092 22898 86134 23134
rect 86370 22898 86412 23134
rect 86092 22866 86412 22898
rect 90040 23454 90360 23486
rect 90040 23218 90082 23454
rect 90318 23218 90360 23454
rect 90040 23134 90360 23218
rect 90040 22898 90082 23134
rect 90318 22898 90360 23134
rect 90040 22866 90360 22898
rect 93988 23454 94308 23486
rect 93988 23218 94030 23454
rect 94266 23218 94308 23454
rect 93988 23134 94308 23218
rect 93988 22898 94030 23134
rect 94266 22898 94308 23134
rect 93988 22866 94308 22898
rect 104892 23454 105212 23486
rect 104892 23218 104934 23454
rect 105170 23218 105212 23454
rect 104892 23134 105212 23218
rect 104892 22898 104934 23134
rect 105170 22898 105212 23134
rect 104892 22866 105212 22898
rect 105840 23454 106160 23486
rect 105840 23218 105882 23454
rect 106118 23218 106160 23454
rect 105840 23134 106160 23218
rect 105840 22898 105882 23134
rect 106118 22898 106160 23134
rect 105840 22866 106160 22898
rect 106788 23454 107108 23486
rect 106788 23218 106830 23454
rect 107066 23218 107108 23454
rect 106788 23134 107108 23218
rect 106788 22898 106830 23134
rect 107066 22898 107108 23134
rect 106788 22866 107108 22898
rect 115092 23454 115412 23486
rect 115092 23218 115134 23454
rect 115370 23218 115412 23454
rect 115092 23134 115412 23218
rect 115092 22898 115134 23134
rect 115370 22898 115412 23134
rect 115092 22866 115412 22898
rect 119040 23454 119360 23486
rect 119040 23218 119082 23454
rect 119318 23218 119360 23454
rect 119040 23134 119360 23218
rect 119040 22898 119082 23134
rect 119318 22898 119360 23134
rect 119040 22866 119360 22898
rect 122988 23454 123308 23486
rect 122988 23218 123030 23454
rect 123266 23218 123308 23454
rect 122988 23134 123308 23218
rect 122988 22898 123030 23134
rect 123266 22898 123308 23134
rect 122988 22866 123308 22898
rect 133892 23454 134212 23486
rect 133892 23218 133934 23454
rect 134170 23218 134212 23454
rect 133892 23134 134212 23218
rect 133892 22898 133934 23134
rect 134170 22898 134212 23134
rect 133892 22866 134212 22898
rect 134840 23454 135160 23486
rect 134840 23218 134882 23454
rect 135118 23218 135160 23454
rect 134840 23134 135160 23218
rect 134840 22898 134882 23134
rect 135118 22898 135160 23134
rect 134840 22866 135160 22898
rect 135788 23454 136108 23486
rect 135788 23218 135830 23454
rect 136066 23218 136108 23454
rect 135788 23134 136108 23218
rect 135788 22898 135830 23134
rect 136066 22898 136108 23134
rect 135788 22866 136108 22898
rect 144092 23454 144412 23486
rect 144092 23218 144134 23454
rect 144370 23218 144412 23454
rect 144092 23134 144412 23218
rect 144092 22898 144134 23134
rect 144370 22898 144412 23134
rect 144092 22866 144412 22898
rect 148040 23454 148360 23486
rect 148040 23218 148082 23454
rect 148318 23218 148360 23454
rect 148040 23134 148360 23218
rect 148040 22898 148082 23134
rect 148318 22898 148360 23134
rect 148040 22866 148360 22898
rect 151988 23454 152308 23486
rect 151988 23218 152030 23454
rect 152266 23218 152308 23454
rect 151988 23134 152308 23218
rect 151988 22898 152030 23134
rect 152266 22898 152308 23134
rect 151988 22866 152308 22898
rect 162892 23454 163212 23486
rect 162892 23218 162934 23454
rect 163170 23218 163212 23454
rect 162892 23134 163212 23218
rect 162892 22898 162934 23134
rect 163170 22898 163212 23134
rect 162892 22866 163212 22898
rect 163840 23454 164160 23486
rect 163840 23218 163882 23454
rect 164118 23218 164160 23454
rect 163840 23134 164160 23218
rect 163840 22898 163882 23134
rect 164118 22898 164160 23134
rect 163840 22866 164160 22898
rect 164788 23454 165108 23486
rect 164788 23218 164830 23454
rect 165066 23218 165108 23454
rect 164788 23134 165108 23218
rect 164788 22898 164830 23134
rect 165066 22898 165108 23134
rect 164788 22866 165108 22898
rect 169710 13157 169770 699755
rect 177994 698454 178614 705242
rect 177994 698218 178026 698454
rect 178262 698218 178346 698454
rect 178582 698218 178614 698454
rect 177994 698134 178614 698218
rect 177994 697898 178026 698134
rect 178262 697898 178346 698134
rect 178582 697898 178614 698134
rect 177994 671454 178614 697898
rect 177994 671218 178026 671454
rect 178262 671218 178346 671454
rect 178582 671218 178614 671454
rect 177994 671134 178614 671218
rect 177994 670898 178026 671134
rect 178262 670898 178346 671134
rect 178582 670898 178614 671134
rect 177994 644454 178614 670898
rect 177994 644218 178026 644454
rect 178262 644218 178346 644454
rect 178582 644218 178614 644454
rect 177994 644134 178614 644218
rect 177994 643898 178026 644134
rect 178262 643898 178346 644134
rect 178582 643898 178614 644134
rect 177994 617454 178614 643898
rect 177994 617218 178026 617454
rect 178262 617218 178346 617454
rect 178582 617218 178614 617454
rect 177994 617134 178614 617218
rect 177994 616898 178026 617134
rect 178262 616898 178346 617134
rect 178582 616898 178614 617134
rect 177994 590454 178614 616898
rect 177994 590218 178026 590454
rect 178262 590218 178346 590454
rect 178582 590218 178614 590454
rect 177994 590134 178614 590218
rect 177994 589898 178026 590134
rect 178262 589898 178346 590134
rect 178582 589898 178614 590134
rect 177994 563454 178614 589898
rect 177994 563218 178026 563454
rect 178262 563218 178346 563454
rect 178582 563218 178614 563454
rect 177994 563134 178614 563218
rect 177994 562898 178026 563134
rect 178262 562898 178346 563134
rect 178582 562898 178614 563134
rect 177994 536454 178614 562898
rect 177994 536218 178026 536454
rect 178262 536218 178346 536454
rect 178582 536218 178614 536454
rect 177994 536134 178614 536218
rect 177994 535898 178026 536134
rect 178262 535898 178346 536134
rect 178582 535898 178614 536134
rect 177994 509454 178614 535898
rect 177994 509218 178026 509454
rect 178262 509218 178346 509454
rect 178582 509218 178614 509454
rect 177994 509134 178614 509218
rect 177994 508898 178026 509134
rect 178262 508898 178346 509134
rect 178582 508898 178614 509134
rect 177994 482454 178614 508898
rect 177994 482218 178026 482454
rect 178262 482218 178346 482454
rect 178582 482218 178614 482454
rect 177994 482134 178614 482218
rect 177994 481898 178026 482134
rect 178262 481898 178346 482134
rect 178582 481898 178614 482134
rect 177994 455454 178614 481898
rect 177994 455218 178026 455454
rect 178262 455218 178346 455454
rect 178582 455218 178614 455454
rect 177994 455134 178614 455218
rect 177994 454898 178026 455134
rect 178262 454898 178346 455134
rect 178582 454898 178614 455134
rect 177994 428454 178614 454898
rect 177994 428218 178026 428454
rect 178262 428218 178346 428454
rect 178582 428218 178614 428454
rect 177994 428134 178614 428218
rect 177994 427898 178026 428134
rect 178262 427898 178346 428134
rect 178582 427898 178614 428134
rect 177994 401454 178614 427898
rect 177994 401218 178026 401454
rect 178262 401218 178346 401454
rect 178582 401218 178614 401454
rect 177994 401134 178614 401218
rect 177994 400898 178026 401134
rect 178262 400898 178346 401134
rect 178582 400898 178614 401134
rect 177994 374454 178614 400898
rect 177994 374218 178026 374454
rect 178262 374218 178346 374454
rect 178582 374218 178614 374454
rect 177994 374134 178614 374218
rect 177994 373898 178026 374134
rect 178262 373898 178346 374134
rect 178582 373898 178614 374134
rect 177994 347454 178614 373898
rect 177994 347218 178026 347454
rect 178262 347218 178346 347454
rect 178582 347218 178614 347454
rect 177994 347134 178614 347218
rect 177994 346898 178026 347134
rect 178262 346898 178346 347134
rect 178582 346898 178614 347134
rect 177994 320454 178614 346898
rect 177994 320218 178026 320454
rect 178262 320218 178346 320454
rect 178582 320218 178614 320454
rect 177994 320134 178614 320218
rect 177994 319898 178026 320134
rect 178262 319898 178346 320134
rect 178582 319898 178614 320134
rect 177994 293454 178614 319898
rect 177994 293218 178026 293454
rect 178262 293218 178346 293454
rect 178582 293218 178614 293454
rect 177994 293134 178614 293218
rect 177994 292898 178026 293134
rect 178262 292898 178346 293134
rect 178582 292898 178614 293134
rect 177994 266454 178614 292898
rect 177994 266218 178026 266454
rect 178262 266218 178346 266454
rect 178582 266218 178614 266454
rect 177994 266134 178614 266218
rect 177994 265898 178026 266134
rect 178262 265898 178346 266134
rect 178582 265898 178614 266134
rect 177994 239454 178614 265898
rect 177994 239218 178026 239454
rect 178262 239218 178346 239454
rect 178582 239218 178614 239454
rect 177994 239134 178614 239218
rect 177994 238898 178026 239134
rect 178262 238898 178346 239134
rect 178582 238898 178614 239134
rect 177994 212454 178614 238898
rect 177994 212218 178026 212454
rect 178262 212218 178346 212454
rect 178582 212218 178614 212454
rect 177994 212134 178614 212218
rect 177994 211898 178026 212134
rect 178262 211898 178346 212134
rect 178582 211898 178614 212134
rect 177994 185454 178614 211898
rect 177994 185218 178026 185454
rect 178262 185218 178346 185454
rect 178582 185218 178614 185454
rect 177994 185134 178614 185218
rect 177994 184898 178026 185134
rect 178262 184898 178346 185134
rect 178582 184898 178614 185134
rect 177994 158454 178614 184898
rect 177994 158218 178026 158454
rect 178262 158218 178346 158454
rect 178582 158218 178614 158454
rect 177994 158134 178614 158218
rect 177994 157898 178026 158134
rect 178262 157898 178346 158134
rect 178582 157898 178614 158134
rect 177994 131454 178614 157898
rect 177994 131218 178026 131454
rect 178262 131218 178346 131454
rect 178582 131218 178614 131454
rect 177994 131134 178614 131218
rect 177994 130898 178026 131134
rect 178262 130898 178346 131134
rect 178582 130898 178614 131134
rect 177994 104454 178614 130898
rect 177994 104218 178026 104454
rect 178262 104218 178346 104454
rect 178582 104218 178614 104454
rect 177994 104134 178614 104218
rect 177994 103898 178026 104134
rect 178262 103898 178346 104134
rect 178582 103898 178614 104134
rect 177994 77454 178614 103898
rect 177994 77218 178026 77454
rect 178262 77218 178346 77454
rect 178582 77218 178614 77454
rect 177994 77134 178614 77218
rect 177994 76898 178026 77134
rect 178262 76898 178346 77134
rect 178582 76898 178614 77134
rect 177994 50454 178614 76898
rect 177994 50218 178026 50454
rect 178262 50218 178346 50454
rect 178582 50218 178614 50454
rect 177994 50134 178614 50218
rect 177994 49898 178026 50134
rect 178262 49898 178346 50134
rect 178582 49898 178614 50134
rect 177994 42000 178614 49898
rect 181494 704838 182114 711590
rect 181494 704602 181526 704838
rect 181762 704602 181846 704838
rect 182082 704602 182114 704838
rect 181494 704518 182114 704602
rect 181494 704282 181526 704518
rect 181762 704282 181846 704518
rect 182082 704282 182114 704518
rect 181494 701829 182114 704282
rect 181494 701593 181526 701829
rect 181762 701593 181846 701829
rect 182082 701593 182114 701829
rect 181494 701509 182114 701593
rect 181494 701273 181526 701509
rect 181762 701273 181846 701509
rect 182082 701273 182114 701509
rect 181494 674829 182114 701273
rect 181494 674593 181526 674829
rect 181762 674593 181846 674829
rect 182082 674593 182114 674829
rect 181494 674509 182114 674593
rect 181494 674273 181526 674509
rect 181762 674273 181846 674509
rect 182082 674273 182114 674509
rect 181494 647829 182114 674273
rect 181494 647593 181526 647829
rect 181762 647593 181846 647829
rect 182082 647593 182114 647829
rect 181494 647509 182114 647593
rect 181494 647273 181526 647509
rect 181762 647273 181846 647509
rect 182082 647273 182114 647509
rect 181494 620829 182114 647273
rect 181494 620593 181526 620829
rect 181762 620593 181846 620829
rect 182082 620593 182114 620829
rect 181494 620509 182114 620593
rect 181494 620273 181526 620509
rect 181762 620273 181846 620509
rect 182082 620273 182114 620509
rect 181494 593829 182114 620273
rect 181494 593593 181526 593829
rect 181762 593593 181846 593829
rect 182082 593593 182114 593829
rect 181494 593509 182114 593593
rect 181494 593273 181526 593509
rect 181762 593273 181846 593509
rect 182082 593273 182114 593509
rect 181494 566829 182114 593273
rect 181494 566593 181526 566829
rect 181762 566593 181846 566829
rect 182082 566593 182114 566829
rect 181494 566509 182114 566593
rect 181494 566273 181526 566509
rect 181762 566273 181846 566509
rect 182082 566273 182114 566509
rect 181494 539829 182114 566273
rect 181494 539593 181526 539829
rect 181762 539593 181846 539829
rect 182082 539593 182114 539829
rect 181494 539509 182114 539593
rect 181494 539273 181526 539509
rect 181762 539273 181846 539509
rect 182082 539273 182114 539509
rect 181494 512829 182114 539273
rect 181494 512593 181526 512829
rect 181762 512593 181846 512829
rect 182082 512593 182114 512829
rect 181494 512509 182114 512593
rect 181494 512273 181526 512509
rect 181762 512273 181846 512509
rect 182082 512273 182114 512509
rect 181494 485829 182114 512273
rect 181494 485593 181526 485829
rect 181762 485593 181846 485829
rect 182082 485593 182114 485829
rect 181494 485509 182114 485593
rect 181494 485273 181526 485509
rect 181762 485273 181846 485509
rect 182082 485273 182114 485509
rect 181494 458829 182114 485273
rect 181494 458593 181526 458829
rect 181762 458593 181846 458829
rect 182082 458593 182114 458829
rect 181494 458509 182114 458593
rect 181494 458273 181526 458509
rect 181762 458273 181846 458509
rect 182082 458273 182114 458509
rect 181494 431829 182114 458273
rect 181494 431593 181526 431829
rect 181762 431593 181846 431829
rect 182082 431593 182114 431829
rect 181494 431509 182114 431593
rect 181494 431273 181526 431509
rect 181762 431273 181846 431509
rect 182082 431273 182114 431509
rect 181494 404829 182114 431273
rect 181494 404593 181526 404829
rect 181762 404593 181846 404829
rect 182082 404593 182114 404829
rect 181494 404509 182114 404593
rect 181494 404273 181526 404509
rect 181762 404273 181846 404509
rect 182082 404273 182114 404509
rect 181494 377829 182114 404273
rect 181494 377593 181526 377829
rect 181762 377593 181846 377829
rect 182082 377593 182114 377829
rect 181494 377509 182114 377593
rect 181494 377273 181526 377509
rect 181762 377273 181846 377509
rect 182082 377273 182114 377509
rect 181494 350829 182114 377273
rect 181494 350593 181526 350829
rect 181762 350593 181846 350829
rect 182082 350593 182114 350829
rect 181494 350509 182114 350593
rect 181494 350273 181526 350509
rect 181762 350273 181846 350509
rect 182082 350273 182114 350509
rect 181494 323829 182114 350273
rect 181494 323593 181526 323829
rect 181762 323593 181846 323829
rect 182082 323593 182114 323829
rect 181494 323509 182114 323593
rect 181494 323273 181526 323509
rect 181762 323273 181846 323509
rect 182082 323273 182114 323509
rect 181494 296829 182114 323273
rect 181494 296593 181526 296829
rect 181762 296593 181846 296829
rect 182082 296593 182114 296829
rect 181494 296509 182114 296593
rect 181494 296273 181526 296509
rect 181762 296273 181846 296509
rect 182082 296273 182114 296509
rect 181494 269829 182114 296273
rect 181494 269593 181526 269829
rect 181762 269593 181846 269829
rect 182082 269593 182114 269829
rect 181494 269509 182114 269593
rect 181494 269273 181526 269509
rect 181762 269273 181846 269509
rect 182082 269273 182114 269509
rect 181494 242829 182114 269273
rect 181494 242593 181526 242829
rect 181762 242593 181846 242829
rect 182082 242593 182114 242829
rect 181494 242509 182114 242593
rect 181494 242273 181526 242509
rect 181762 242273 181846 242509
rect 182082 242273 182114 242509
rect 181494 215829 182114 242273
rect 181494 215593 181526 215829
rect 181762 215593 181846 215829
rect 182082 215593 182114 215829
rect 181494 215509 182114 215593
rect 181494 215273 181526 215509
rect 181762 215273 181846 215509
rect 182082 215273 182114 215509
rect 181494 188829 182114 215273
rect 181494 188593 181526 188829
rect 181762 188593 181846 188829
rect 182082 188593 182114 188829
rect 181494 188509 182114 188593
rect 181494 188273 181526 188509
rect 181762 188273 181846 188509
rect 182082 188273 182114 188509
rect 181494 161829 182114 188273
rect 181494 161593 181526 161829
rect 181762 161593 181846 161829
rect 182082 161593 182114 161829
rect 181494 161509 182114 161593
rect 181494 161273 181526 161509
rect 181762 161273 181846 161509
rect 182082 161273 182114 161509
rect 181494 134829 182114 161273
rect 181494 134593 181526 134829
rect 181762 134593 181846 134829
rect 182082 134593 182114 134829
rect 181494 134509 182114 134593
rect 181494 134273 181526 134509
rect 181762 134273 181846 134509
rect 182082 134273 182114 134509
rect 181494 107829 182114 134273
rect 181494 107593 181526 107829
rect 181762 107593 181846 107829
rect 182082 107593 182114 107829
rect 181494 107509 182114 107593
rect 181494 107273 181526 107509
rect 181762 107273 181846 107509
rect 182082 107273 182114 107509
rect 181494 80829 182114 107273
rect 181494 80593 181526 80829
rect 181762 80593 181846 80829
rect 182082 80593 182114 80829
rect 181494 80509 182114 80593
rect 181494 80273 181526 80509
rect 181762 80273 181846 80509
rect 182082 80273 182114 80509
rect 181494 53829 182114 80273
rect 205994 705798 206614 711590
rect 205994 705562 206026 705798
rect 206262 705562 206346 705798
rect 206582 705562 206614 705798
rect 205994 705478 206614 705562
rect 205994 705242 206026 705478
rect 206262 705242 206346 705478
rect 206582 705242 206614 705478
rect 205994 698454 206614 705242
rect 205994 698218 206026 698454
rect 206262 698218 206346 698454
rect 206582 698218 206614 698454
rect 205994 698134 206614 698218
rect 205994 697898 206026 698134
rect 206262 697898 206346 698134
rect 206582 697898 206614 698134
rect 205994 671454 206614 697898
rect 205994 671218 206026 671454
rect 206262 671218 206346 671454
rect 206582 671218 206614 671454
rect 205994 671134 206614 671218
rect 205994 670898 206026 671134
rect 206262 670898 206346 671134
rect 206582 670898 206614 671134
rect 205994 644454 206614 670898
rect 205994 644218 206026 644454
rect 206262 644218 206346 644454
rect 206582 644218 206614 644454
rect 205994 644134 206614 644218
rect 205994 643898 206026 644134
rect 206262 643898 206346 644134
rect 206582 643898 206614 644134
rect 205994 617454 206614 643898
rect 205994 617218 206026 617454
rect 206262 617218 206346 617454
rect 206582 617218 206614 617454
rect 205994 617134 206614 617218
rect 205994 616898 206026 617134
rect 206262 616898 206346 617134
rect 206582 616898 206614 617134
rect 205994 590454 206614 616898
rect 205994 590218 206026 590454
rect 206262 590218 206346 590454
rect 206582 590218 206614 590454
rect 205994 590134 206614 590218
rect 205994 589898 206026 590134
rect 206262 589898 206346 590134
rect 206582 589898 206614 590134
rect 205994 563454 206614 589898
rect 205994 563218 206026 563454
rect 206262 563218 206346 563454
rect 206582 563218 206614 563454
rect 205994 563134 206614 563218
rect 205994 562898 206026 563134
rect 206262 562898 206346 563134
rect 206582 562898 206614 563134
rect 205994 536454 206614 562898
rect 205994 536218 206026 536454
rect 206262 536218 206346 536454
rect 206582 536218 206614 536454
rect 205994 536134 206614 536218
rect 205994 535898 206026 536134
rect 206262 535898 206346 536134
rect 206582 535898 206614 536134
rect 205994 509454 206614 535898
rect 205994 509218 206026 509454
rect 206262 509218 206346 509454
rect 206582 509218 206614 509454
rect 205994 509134 206614 509218
rect 205994 508898 206026 509134
rect 206262 508898 206346 509134
rect 206582 508898 206614 509134
rect 205994 482454 206614 508898
rect 205994 482218 206026 482454
rect 206262 482218 206346 482454
rect 206582 482218 206614 482454
rect 205994 482134 206614 482218
rect 205994 481898 206026 482134
rect 206262 481898 206346 482134
rect 206582 481898 206614 482134
rect 205994 455454 206614 481898
rect 205994 455218 206026 455454
rect 206262 455218 206346 455454
rect 206582 455218 206614 455454
rect 205994 455134 206614 455218
rect 205994 454898 206026 455134
rect 206262 454898 206346 455134
rect 206582 454898 206614 455134
rect 205994 428454 206614 454898
rect 205994 428218 206026 428454
rect 206262 428218 206346 428454
rect 206582 428218 206614 428454
rect 205994 428134 206614 428218
rect 205994 427898 206026 428134
rect 206262 427898 206346 428134
rect 206582 427898 206614 428134
rect 205994 401454 206614 427898
rect 205994 401218 206026 401454
rect 206262 401218 206346 401454
rect 206582 401218 206614 401454
rect 205994 401134 206614 401218
rect 205994 400898 206026 401134
rect 206262 400898 206346 401134
rect 206582 400898 206614 401134
rect 205994 374454 206614 400898
rect 205994 374218 206026 374454
rect 206262 374218 206346 374454
rect 206582 374218 206614 374454
rect 205994 374134 206614 374218
rect 205994 373898 206026 374134
rect 206262 373898 206346 374134
rect 206582 373898 206614 374134
rect 205994 347454 206614 373898
rect 205994 347218 206026 347454
rect 206262 347218 206346 347454
rect 206582 347218 206614 347454
rect 205994 347134 206614 347218
rect 205994 346898 206026 347134
rect 206262 346898 206346 347134
rect 206582 346898 206614 347134
rect 205994 320454 206614 346898
rect 205994 320218 206026 320454
rect 206262 320218 206346 320454
rect 206582 320218 206614 320454
rect 205994 320134 206614 320218
rect 205994 319898 206026 320134
rect 206262 319898 206346 320134
rect 206582 319898 206614 320134
rect 205994 293454 206614 319898
rect 205994 293218 206026 293454
rect 206262 293218 206346 293454
rect 206582 293218 206614 293454
rect 205994 293134 206614 293218
rect 205994 292898 206026 293134
rect 206262 292898 206346 293134
rect 206582 292898 206614 293134
rect 205994 266454 206614 292898
rect 205994 266218 206026 266454
rect 206262 266218 206346 266454
rect 206582 266218 206614 266454
rect 205994 266134 206614 266218
rect 205994 265898 206026 266134
rect 206262 265898 206346 266134
rect 206582 265898 206614 266134
rect 205994 239454 206614 265898
rect 205994 239218 206026 239454
rect 206262 239218 206346 239454
rect 206582 239218 206614 239454
rect 205994 239134 206614 239218
rect 205994 238898 206026 239134
rect 206262 238898 206346 239134
rect 206582 238898 206614 239134
rect 205994 212454 206614 238898
rect 205994 212218 206026 212454
rect 206262 212218 206346 212454
rect 206582 212218 206614 212454
rect 205994 212134 206614 212218
rect 205994 211898 206026 212134
rect 206262 211898 206346 212134
rect 206582 211898 206614 212134
rect 205994 185454 206614 211898
rect 205994 185218 206026 185454
rect 206262 185218 206346 185454
rect 206582 185218 206614 185454
rect 205994 185134 206614 185218
rect 205994 184898 206026 185134
rect 206262 184898 206346 185134
rect 206582 184898 206614 185134
rect 205994 158454 206614 184898
rect 205994 158218 206026 158454
rect 206262 158218 206346 158454
rect 206582 158218 206614 158454
rect 205994 158134 206614 158218
rect 205994 157898 206026 158134
rect 206262 157898 206346 158134
rect 206582 157898 206614 158134
rect 205994 131454 206614 157898
rect 205994 131218 206026 131454
rect 206262 131218 206346 131454
rect 206582 131218 206614 131454
rect 205994 131134 206614 131218
rect 205994 130898 206026 131134
rect 206262 130898 206346 131134
rect 206582 130898 206614 131134
rect 205994 104454 206614 130898
rect 205994 104218 206026 104454
rect 206262 104218 206346 104454
rect 206582 104218 206614 104454
rect 205994 104134 206614 104218
rect 205994 103898 206026 104134
rect 206262 103898 206346 104134
rect 206582 103898 206614 104134
rect 205994 77454 206614 103898
rect 205994 77218 206026 77454
rect 206262 77218 206346 77454
rect 206582 77218 206614 77454
rect 205994 77134 206614 77218
rect 205994 76898 206026 77134
rect 206262 76898 206346 77134
rect 206582 76898 206614 77134
rect 205994 69000 206614 76898
rect 209494 704838 210114 711590
rect 209494 704602 209526 704838
rect 209762 704602 209846 704838
rect 210082 704602 210114 704838
rect 209494 704518 210114 704602
rect 209494 704282 209526 704518
rect 209762 704282 209846 704518
rect 210082 704282 210114 704518
rect 209494 701829 210114 704282
rect 209494 701593 209526 701829
rect 209762 701593 209846 701829
rect 210082 701593 210114 701829
rect 209494 701509 210114 701593
rect 209494 701273 209526 701509
rect 209762 701273 209846 701509
rect 210082 701273 210114 701509
rect 209494 674829 210114 701273
rect 209494 674593 209526 674829
rect 209762 674593 209846 674829
rect 210082 674593 210114 674829
rect 209494 674509 210114 674593
rect 209494 674273 209526 674509
rect 209762 674273 209846 674509
rect 210082 674273 210114 674509
rect 209494 647829 210114 674273
rect 209494 647593 209526 647829
rect 209762 647593 209846 647829
rect 210082 647593 210114 647829
rect 209494 647509 210114 647593
rect 209494 647273 209526 647509
rect 209762 647273 209846 647509
rect 210082 647273 210114 647509
rect 209494 620829 210114 647273
rect 209494 620593 209526 620829
rect 209762 620593 209846 620829
rect 210082 620593 210114 620829
rect 209494 620509 210114 620593
rect 209494 620273 209526 620509
rect 209762 620273 209846 620509
rect 210082 620273 210114 620509
rect 209494 593829 210114 620273
rect 209494 593593 209526 593829
rect 209762 593593 209846 593829
rect 210082 593593 210114 593829
rect 209494 593509 210114 593593
rect 209494 593273 209526 593509
rect 209762 593273 209846 593509
rect 210082 593273 210114 593509
rect 209494 566829 210114 593273
rect 209494 566593 209526 566829
rect 209762 566593 209846 566829
rect 210082 566593 210114 566829
rect 209494 566509 210114 566593
rect 209494 566273 209526 566509
rect 209762 566273 209846 566509
rect 210082 566273 210114 566509
rect 209494 539829 210114 566273
rect 209494 539593 209526 539829
rect 209762 539593 209846 539829
rect 210082 539593 210114 539829
rect 209494 539509 210114 539593
rect 209494 539273 209526 539509
rect 209762 539273 209846 539509
rect 210082 539273 210114 539509
rect 209494 512829 210114 539273
rect 209494 512593 209526 512829
rect 209762 512593 209846 512829
rect 210082 512593 210114 512829
rect 209494 512509 210114 512593
rect 209494 512273 209526 512509
rect 209762 512273 209846 512509
rect 210082 512273 210114 512509
rect 209494 485829 210114 512273
rect 209494 485593 209526 485829
rect 209762 485593 209846 485829
rect 210082 485593 210114 485829
rect 209494 485509 210114 485593
rect 209494 485273 209526 485509
rect 209762 485273 209846 485509
rect 210082 485273 210114 485509
rect 209494 458829 210114 485273
rect 209494 458593 209526 458829
rect 209762 458593 209846 458829
rect 210082 458593 210114 458829
rect 209494 458509 210114 458593
rect 209494 458273 209526 458509
rect 209762 458273 209846 458509
rect 210082 458273 210114 458509
rect 209494 431829 210114 458273
rect 209494 431593 209526 431829
rect 209762 431593 209846 431829
rect 210082 431593 210114 431829
rect 209494 431509 210114 431593
rect 209494 431273 209526 431509
rect 209762 431273 209846 431509
rect 210082 431273 210114 431509
rect 209494 404829 210114 431273
rect 209494 404593 209526 404829
rect 209762 404593 209846 404829
rect 210082 404593 210114 404829
rect 209494 404509 210114 404593
rect 209494 404273 209526 404509
rect 209762 404273 209846 404509
rect 210082 404273 210114 404509
rect 209494 377829 210114 404273
rect 209494 377593 209526 377829
rect 209762 377593 209846 377829
rect 210082 377593 210114 377829
rect 209494 377509 210114 377593
rect 209494 377273 209526 377509
rect 209762 377273 209846 377509
rect 210082 377273 210114 377509
rect 209494 350829 210114 377273
rect 209494 350593 209526 350829
rect 209762 350593 209846 350829
rect 210082 350593 210114 350829
rect 209494 350509 210114 350593
rect 209494 350273 209526 350509
rect 209762 350273 209846 350509
rect 210082 350273 210114 350509
rect 209494 323829 210114 350273
rect 209494 323593 209526 323829
rect 209762 323593 209846 323829
rect 210082 323593 210114 323829
rect 209494 323509 210114 323593
rect 209494 323273 209526 323509
rect 209762 323273 209846 323509
rect 210082 323273 210114 323509
rect 209494 296829 210114 323273
rect 209494 296593 209526 296829
rect 209762 296593 209846 296829
rect 210082 296593 210114 296829
rect 209494 296509 210114 296593
rect 209494 296273 209526 296509
rect 209762 296273 209846 296509
rect 210082 296273 210114 296509
rect 209494 269829 210114 296273
rect 209494 269593 209526 269829
rect 209762 269593 209846 269829
rect 210082 269593 210114 269829
rect 209494 269509 210114 269593
rect 209494 269273 209526 269509
rect 209762 269273 209846 269509
rect 210082 269273 210114 269509
rect 209494 242829 210114 269273
rect 209494 242593 209526 242829
rect 209762 242593 209846 242829
rect 210082 242593 210114 242829
rect 209494 242509 210114 242593
rect 209494 242273 209526 242509
rect 209762 242273 209846 242509
rect 210082 242273 210114 242509
rect 209494 215829 210114 242273
rect 209494 215593 209526 215829
rect 209762 215593 209846 215829
rect 210082 215593 210114 215829
rect 209494 215509 210114 215593
rect 209494 215273 209526 215509
rect 209762 215273 209846 215509
rect 210082 215273 210114 215509
rect 209494 188829 210114 215273
rect 209494 188593 209526 188829
rect 209762 188593 209846 188829
rect 210082 188593 210114 188829
rect 209494 188509 210114 188593
rect 209494 188273 209526 188509
rect 209762 188273 209846 188509
rect 210082 188273 210114 188509
rect 209494 161829 210114 188273
rect 209494 161593 209526 161829
rect 209762 161593 209846 161829
rect 210082 161593 210114 161829
rect 209494 161509 210114 161593
rect 209494 161273 209526 161509
rect 209762 161273 209846 161509
rect 210082 161273 210114 161509
rect 209494 134829 210114 161273
rect 209494 134593 209526 134829
rect 209762 134593 209846 134829
rect 210082 134593 210114 134829
rect 209494 134509 210114 134593
rect 209494 134273 209526 134509
rect 209762 134273 209846 134509
rect 210082 134273 210114 134509
rect 209494 107829 210114 134273
rect 209494 107593 209526 107829
rect 209762 107593 209846 107829
rect 210082 107593 210114 107829
rect 209494 107509 210114 107593
rect 209494 107273 209526 107509
rect 209762 107273 209846 107509
rect 210082 107273 210114 107509
rect 209494 80829 210114 107273
rect 209494 80593 209526 80829
rect 209762 80593 209846 80829
rect 210082 80593 210114 80829
rect 209494 80509 210114 80593
rect 209494 80273 209526 80509
rect 209762 80273 209846 80509
rect 210082 80273 210114 80509
rect 209494 69000 210114 80273
rect 233994 705798 234614 711590
rect 233994 705562 234026 705798
rect 234262 705562 234346 705798
rect 234582 705562 234614 705798
rect 233994 705478 234614 705562
rect 233994 705242 234026 705478
rect 234262 705242 234346 705478
rect 234582 705242 234614 705478
rect 233994 698454 234614 705242
rect 233994 698218 234026 698454
rect 234262 698218 234346 698454
rect 234582 698218 234614 698454
rect 233994 698134 234614 698218
rect 233994 697898 234026 698134
rect 234262 697898 234346 698134
rect 234582 697898 234614 698134
rect 233994 671454 234614 697898
rect 233994 671218 234026 671454
rect 234262 671218 234346 671454
rect 234582 671218 234614 671454
rect 233994 671134 234614 671218
rect 233994 670898 234026 671134
rect 234262 670898 234346 671134
rect 234582 670898 234614 671134
rect 233994 644454 234614 670898
rect 233994 644218 234026 644454
rect 234262 644218 234346 644454
rect 234582 644218 234614 644454
rect 233994 644134 234614 644218
rect 233994 643898 234026 644134
rect 234262 643898 234346 644134
rect 234582 643898 234614 644134
rect 233994 617454 234614 643898
rect 233994 617218 234026 617454
rect 234262 617218 234346 617454
rect 234582 617218 234614 617454
rect 233994 617134 234614 617218
rect 233994 616898 234026 617134
rect 234262 616898 234346 617134
rect 234582 616898 234614 617134
rect 233994 590454 234614 616898
rect 233994 590218 234026 590454
rect 234262 590218 234346 590454
rect 234582 590218 234614 590454
rect 233994 590134 234614 590218
rect 233994 589898 234026 590134
rect 234262 589898 234346 590134
rect 234582 589898 234614 590134
rect 233994 563454 234614 589898
rect 233994 563218 234026 563454
rect 234262 563218 234346 563454
rect 234582 563218 234614 563454
rect 233994 563134 234614 563218
rect 233994 562898 234026 563134
rect 234262 562898 234346 563134
rect 234582 562898 234614 563134
rect 233994 536454 234614 562898
rect 233994 536218 234026 536454
rect 234262 536218 234346 536454
rect 234582 536218 234614 536454
rect 233994 536134 234614 536218
rect 233994 535898 234026 536134
rect 234262 535898 234346 536134
rect 234582 535898 234614 536134
rect 233994 509454 234614 535898
rect 233994 509218 234026 509454
rect 234262 509218 234346 509454
rect 234582 509218 234614 509454
rect 233994 509134 234614 509218
rect 233994 508898 234026 509134
rect 234262 508898 234346 509134
rect 234582 508898 234614 509134
rect 233994 482454 234614 508898
rect 233994 482218 234026 482454
rect 234262 482218 234346 482454
rect 234582 482218 234614 482454
rect 233994 482134 234614 482218
rect 233994 481898 234026 482134
rect 234262 481898 234346 482134
rect 234582 481898 234614 482134
rect 233994 455454 234614 481898
rect 233994 455218 234026 455454
rect 234262 455218 234346 455454
rect 234582 455218 234614 455454
rect 233994 455134 234614 455218
rect 233994 454898 234026 455134
rect 234262 454898 234346 455134
rect 234582 454898 234614 455134
rect 233994 428454 234614 454898
rect 233994 428218 234026 428454
rect 234262 428218 234346 428454
rect 234582 428218 234614 428454
rect 233994 428134 234614 428218
rect 233994 427898 234026 428134
rect 234262 427898 234346 428134
rect 234582 427898 234614 428134
rect 233994 401454 234614 427898
rect 233994 401218 234026 401454
rect 234262 401218 234346 401454
rect 234582 401218 234614 401454
rect 233994 401134 234614 401218
rect 233994 400898 234026 401134
rect 234262 400898 234346 401134
rect 234582 400898 234614 401134
rect 233994 374454 234614 400898
rect 233994 374218 234026 374454
rect 234262 374218 234346 374454
rect 234582 374218 234614 374454
rect 233994 374134 234614 374218
rect 233994 373898 234026 374134
rect 234262 373898 234346 374134
rect 234582 373898 234614 374134
rect 233994 347454 234614 373898
rect 233994 347218 234026 347454
rect 234262 347218 234346 347454
rect 234582 347218 234614 347454
rect 233994 347134 234614 347218
rect 233994 346898 234026 347134
rect 234262 346898 234346 347134
rect 234582 346898 234614 347134
rect 233994 320454 234614 346898
rect 233994 320218 234026 320454
rect 234262 320218 234346 320454
rect 234582 320218 234614 320454
rect 233994 320134 234614 320218
rect 233994 319898 234026 320134
rect 234262 319898 234346 320134
rect 234582 319898 234614 320134
rect 233994 293454 234614 319898
rect 233994 293218 234026 293454
rect 234262 293218 234346 293454
rect 234582 293218 234614 293454
rect 233994 293134 234614 293218
rect 233994 292898 234026 293134
rect 234262 292898 234346 293134
rect 234582 292898 234614 293134
rect 233994 266454 234614 292898
rect 233994 266218 234026 266454
rect 234262 266218 234346 266454
rect 234582 266218 234614 266454
rect 233994 266134 234614 266218
rect 233994 265898 234026 266134
rect 234262 265898 234346 266134
rect 234582 265898 234614 266134
rect 233994 239454 234614 265898
rect 233994 239218 234026 239454
rect 234262 239218 234346 239454
rect 234582 239218 234614 239454
rect 233994 239134 234614 239218
rect 233994 238898 234026 239134
rect 234262 238898 234346 239134
rect 234582 238898 234614 239134
rect 233994 212454 234614 238898
rect 233994 212218 234026 212454
rect 234262 212218 234346 212454
rect 234582 212218 234614 212454
rect 233994 212134 234614 212218
rect 233994 211898 234026 212134
rect 234262 211898 234346 212134
rect 234582 211898 234614 212134
rect 233994 185454 234614 211898
rect 233994 185218 234026 185454
rect 234262 185218 234346 185454
rect 234582 185218 234614 185454
rect 233994 185134 234614 185218
rect 233994 184898 234026 185134
rect 234262 184898 234346 185134
rect 234582 184898 234614 185134
rect 233994 158454 234614 184898
rect 233994 158218 234026 158454
rect 234262 158218 234346 158454
rect 234582 158218 234614 158454
rect 233994 158134 234614 158218
rect 233994 157898 234026 158134
rect 234262 157898 234346 158134
rect 234582 157898 234614 158134
rect 233994 131454 234614 157898
rect 233994 131218 234026 131454
rect 234262 131218 234346 131454
rect 234582 131218 234614 131454
rect 233994 131134 234614 131218
rect 233994 130898 234026 131134
rect 234262 130898 234346 131134
rect 234582 130898 234614 131134
rect 233994 104454 234614 130898
rect 233994 104218 234026 104454
rect 234262 104218 234346 104454
rect 234582 104218 234614 104454
rect 233994 104134 234614 104218
rect 233994 103898 234026 104134
rect 234262 103898 234346 104134
rect 234582 103898 234614 104134
rect 233994 77454 234614 103898
rect 233994 77218 234026 77454
rect 234262 77218 234346 77454
rect 234582 77218 234614 77454
rect 233994 77134 234614 77218
rect 233994 76898 234026 77134
rect 234262 76898 234346 77134
rect 234582 76898 234614 77134
rect 233994 69000 234614 76898
rect 237494 704838 238114 711590
rect 237494 704602 237526 704838
rect 237762 704602 237846 704838
rect 238082 704602 238114 704838
rect 237494 704518 238114 704602
rect 237494 704282 237526 704518
rect 237762 704282 237846 704518
rect 238082 704282 238114 704518
rect 237494 701829 238114 704282
rect 237494 701593 237526 701829
rect 237762 701593 237846 701829
rect 238082 701593 238114 701829
rect 237494 701509 238114 701593
rect 237494 701273 237526 701509
rect 237762 701273 237846 701509
rect 238082 701273 238114 701509
rect 237494 674829 238114 701273
rect 237494 674593 237526 674829
rect 237762 674593 237846 674829
rect 238082 674593 238114 674829
rect 237494 674509 238114 674593
rect 237494 674273 237526 674509
rect 237762 674273 237846 674509
rect 238082 674273 238114 674509
rect 237494 647829 238114 674273
rect 237494 647593 237526 647829
rect 237762 647593 237846 647829
rect 238082 647593 238114 647829
rect 237494 647509 238114 647593
rect 237494 647273 237526 647509
rect 237762 647273 237846 647509
rect 238082 647273 238114 647509
rect 237494 620829 238114 647273
rect 237494 620593 237526 620829
rect 237762 620593 237846 620829
rect 238082 620593 238114 620829
rect 237494 620509 238114 620593
rect 237494 620273 237526 620509
rect 237762 620273 237846 620509
rect 238082 620273 238114 620509
rect 237494 593829 238114 620273
rect 237494 593593 237526 593829
rect 237762 593593 237846 593829
rect 238082 593593 238114 593829
rect 237494 593509 238114 593593
rect 237494 593273 237526 593509
rect 237762 593273 237846 593509
rect 238082 593273 238114 593509
rect 237494 566829 238114 593273
rect 237494 566593 237526 566829
rect 237762 566593 237846 566829
rect 238082 566593 238114 566829
rect 237494 566509 238114 566593
rect 237494 566273 237526 566509
rect 237762 566273 237846 566509
rect 238082 566273 238114 566509
rect 237494 539829 238114 566273
rect 237494 539593 237526 539829
rect 237762 539593 237846 539829
rect 238082 539593 238114 539829
rect 237494 539509 238114 539593
rect 237494 539273 237526 539509
rect 237762 539273 237846 539509
rect 238082 539273 238114 539509
rect 237494 512829 238114 539273
rect 237494 512593 237526 512829
rect 237762 512593 237846 512829
rect 238082 512593 238114 512829
rect 237494 512509 238114 512593
rect 237494 512273 237526 512509
rect 237762 512273 237846 512509
rect 238082 512273 238114 512509
rect 237494 485829 238114 512273
rect 237494 485593 237526 485829
rect 237762 485593 237846 485829
rect 238082 485593 238114 485829
rect 237494 485509 238114 485593
rect 237494 485273 237526 485509
rect 237762 485273 237846 485509
rect 238082 485273 238114 485509
rect 237494 458829 238114 485273
rect 237494 458593 237526 458829
rect 237762 458593 237846 458829
rect 238082 458593 238114 458829
rect 237494 458509 238114 458593
rect 237494 458273 237526 458509
rect 237762 458273 237846 458509
rect 238082 458273 238114 458509
rect 237494 431829 238114 458273
rect 237494 431593 237526 431829
rect 237762 431593 237846 431829
rect 238082 431593 238114 431829
rect 237494 431509 238114 431593
rect 237494 431273 237526 431509
rect 237762 431273 237846 431509
rect 238082 431273 238114 431509
rect 237494 404829 238114 431273
rect 237494 404593 237526 404829
rect 237762 404593 237846 404829
rect 238082 404593 238114 404829
rect 237494 404509 238114 404593
rect 237494 404273 237526 404509
rect 237762 404273 237846 404509
rect 238082 404273 238114 404509
rect 237494 377829 238114 404273
rect 237494 377593 237526 377829
rect 237762 377593 237846 377829
rect 238082 377593 238114 377829
rect 237494 377509 238114 377593
rect 237494 377273 237526 377509
rect 237762 377273 237846 377509
rect 238082 377273 238114 377509
rect 237494 350829 238114 377273
rect 237494 350593 237526 350829
rect 237762 350593 237846 350829
rect 238082 350593 238114 350829
rect 237494 350509 238114 350593
rect 237494 350273 237526 350509
rect 237762 350273 237846 350509
rect 238082 350273 238114 350509
rect 237494 323829 238114 350273
rect 237494 323593 237526 323829
rect 237762 323593 237846 323829
rect 238082 323593 238114 323829
rect 237494 323509 238114 323593
rect 237494 323273 237526 323509
rect 237762 323273 237846 323509
rect 238082 323273 238114 323509
rect 237494 296829 238114 323273
rect 237494 296593 237526 296829
rect 237762 296593 237846 296829
rect 238082 296593 238114 296829
rect 237494 296509 238114 296593
rect 237494 296273 237526 296509
rect 237762 296273 237846 296509
rect 238082 296273 238114 296509
rect 237494 269829 238114 296273
rect 237494 269593 237526 269829
rect 237762 269593 237846 269829
rect 238082 269593 238114 269829
rect 237494 269509 238114 269593
rect 237494 269273 237526 269509
rect 237762 269273 237846 269509
rect 238082 269273 238114 269509
rect 237494 242829 238114 269273
rect 237494 242593 237526 242829
rect 237762 242593 237846 242829
rect 238082 242593 238114 242829
rect 237494 242509 238114 242593
rect 237494 242273 237526 242509
rect 237762 242273 237846 242509
rect 238082 242273 238114 242509
rect 237494 215829 238114 242273
rect 237494 215593 237526 215829
rect 237762 215593 237846 215829
rect 238082 215593 238114 215829
rect 237494 215509 238114 215593
rect 237494 215273 237526 215509
rect 237762 215273 237846 215509
rect 238082 215273 238114 215509
rect 237494 188829 238114 215273
rect 237494 188593 237526 188829
rect 237762 188593 237846 188829
rect 238082 188593 238114 188829
rect 237494 188509 238114 188593
rect 237494 188273 237526 188509
rect 237762 188273 237846 188509
rect 238082 188273 238114 188509
rect 237494 161829 238114 188273
rect 237494 161593 237526 161829
rect 237762 161593 237846 161829
rect 238082 161593 238114 161829
rect 237494 161509 238114 161593
rect 237494 161273 237526 161509
rect 237762 161273 237846 161509
rect 238082 161273 238114 161509
rect 237494 134829 238114 161273
rect 237494 134593 237526 134829
rect 237762 134593 237846 134829
rect 238082 134593 238114 134829
rect 237494 134509 238114 134593
rect 237494 134273 237526 134509
rect 237762 134273 237846 134509
rect 238082 134273 238114 134509
rect 237494 107829 238114 134273
rect 237494 107593 237526 107829
rect 237762 107593 237846 107829
rect 238082 107593 238114 107829
rect 237494 107509 238114 107593
rect 237494 107273 237526 107509
rect 237762 107273 237846 107509
rect 238082 107273 238114 107509
rect 237494 80829 238114 107273
rect 237494 80593 237526 80829
rect 237762 80593 237846 80829
rect 238082 80593 238114 80829
rect 237494 80509 238114 80593
rect 237494 80273 237526 80509
rect 237762 80273 237846 80509
rect 238082 80273 238114 80509
rect 237494 69000 238114 80273
rect 261994 705798 262614 711590
rect 261994 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 262614 705798
rect 261994 705478 262614 705562
rect 261994 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 262614 705478
rect 261994 698454 262614 705242
rect 261994 698218 262026 698454
rect 262262 698218 262346 698454
rect 262582 698218 262614 698454
rect 261994 698134 262614 698218
rect 261994 697898 262026 698134
rect 262262 697898 262346 698134
rect 262582 697898 262614 698134
rect 261994 671454 262614 697898
rect 261994 671218 262026 671454
rect 262262 671218 262346 671454
rect 262582 671218 262614 671454
rect 261994 671134 262614 671218
rect 261994 670898 262026 671134
rect 262262 670898 262346 671134
rect 262582 670898 262614 671134
rect 261994 644454 262614 670898
rect 261994 644218 262026 644454
rect 262262 644218 262346 644454
rect 262582 644218 262614 644454
rect 261994 644134 262614 644218
rect 261994 643898 262026 644134
rect 262262 643898 262346 644134
rect 262582 643898 262614 644134
rect 261994 617454 262614 643898
rect 261994 617218 262026 617454
rect 262262 617218 262346 617454
rect 262582 617218 262614 617454
rect 261994 617134 262614 617218
rect 261994 616898 262026 617134
rect 262262 616898 262346 617134
rect 262582 616898 262614 617134
rect 261994 590454 262614 616898
rect 261994 590218 262026 590454
rect 262262 590218 262346 590454
rect 262582 590218 262614 590454
rect 261994 590134 262614 590218
rect 261994 589898 262026 590134
rect 262262 589898 262346 590134
rect 262582 589898 262614 590134
rect 261994 563454 262614 589898
rect 261994 563218 262026 563454
rect 262262 563218 262346 563454
rect 262582 563218 262614 563454
rect 261994 563134 262614 563218
rect 261994 562898 262026 563134
rect 262262 562898 262346 563134
rect 262582 562898 262614 563134
rect 261994 536454 262614 562898
rect 261994 536218 262026 536454
rect 262262 536218 262346 536454
rect 262582 536218 262614 536454
rect 261994 536134 262614 536218
rect 261994 535898 262026 536134
rect 262262 535898 262346 536134
rect 262582 535898 262614 536134
rect 261994 509454 262614 535898
rect 261994 509218 262026 509454
rect 262262 509218 262346 509454
rect 262582 509218 262614 509454
rect 261994 509134 262614 509218
rect 261994 508898 262026 509134
rect 262262 508898 262346 509134
rect 262582 508898 262614 509134
rect 261994 482454 262614 508898
rect 261994 482218 262026 482454
rect 262262 482218 262346 482454
rect 262582 482218 262614 482454
rect 261994 482134 262614 482218
rect 261994 481898 262026 482134
rect 262262 481898 262346 482134
rect 262582 481898 262614 482134
rect 261994 455454 262614 481898
rect 261994 455218 262026 455454
rect 262262 455218 262346 455454
rect 262582 455218 262614 455454
rect 261994 455134 262614 455218
rect 261994 454898 262026 455134
rect 262262 454898 262346 455134
rect 262582 454898 262614 455134
rect 261994 428454 262614 454898
rect 261994 428218 262026 428454
rect 262262 428218 262346 428454
rect 262582 428218 262614 428454
rect 261994 428134 262614 428218
rect 261994 427898 262026 428134
rect 262262 427898 262346 428134
rect 262582 427898 262614 428134
rect 261994 401454 262614 427898
rect 261994 401218 262026 401454
rect 262262 401218 262346 401454
rect 262582 401218 262614 401454
rect 261994 401134 262614 401218
rect 261994 400898 262026 401134
rect 262262 400898 262346 401134
rect 262582 400898 262614 401134
rect 261994 374454 262614 400898
rect 261994 374218 262026 374454
rect 262262 374218 262346 374454
rect 262582 374218 262614 374454
rect 261994 374134 262614 374218
rect 261994 373898 262026 374134
rect 262262 373898 262346 374134
rect 262582 373898 262614 374134
rect 261994 347454 262614 373898
rect 261994 347218 262026 347454
rect 262262 347218 262346 347454
rect 262582 347218 262614 347454
rect 261994 347134 262614 347218
rect 261994 346898 262026 347134
rect 262262 346898 262346 347134
rect 262582 346898 262614 347134
rect 261994 320454 262614 346898
rect 261994 320218 262026 320454
rect 262262 320218 262346 320454
rect 262582 320218 262614 320454
rect 261994 320134 262614 320218
rect 261994 319898 262026 320134
rect 262262 319898 262346 320134
rect 262582 319898 262614 320134
rect 261994 293454 262614 319898
rect 261994 293218 262026 293454
rect 262262 293218 262346 293454
rect 262582 293218 262614 293454
rect 261994 293134 262614 293218
rect 261994 292898 262026 293134
rect 262262 292898 262346 293134
rect 262582 292898 262614 293134
rect 261994 266454 262614 292898
rect 261994 266218 262026 266454
rect 262262 266218 262346 266454
rect 262582 266218 262614 266454
rect 261994 266134 262614 266218
rect 261994 265898 262026 266134
rect 262262 265898 262346 266134
rect 262582 265898 262614 266134
rect 261994 239454 262614 265898
rect 261994 239218 262026 239454
rect 262262 239218 262346 239454
rect 262582 239218 262614 239454
rect 261994 239134 262614 239218
rect 261994 238898 262026 239134
rect 262262 238898 262346 239134
rect 262582 238898 262614 239134
rect 261994 212454 262614 238898
rect 261994 212218 262026 212454
rect 262262 212218 262346 212454
rect 262582 212218 262614 212454
rect 261994 212134 262614 212218
rect 261994 211898 262026 212134
rect 262262 211898 262346 212134
rect 262582 211898 262614 212134
rect 261994 185454 262614 211898
rect 261994 185218 262026 185454
rect 262262 185218 262346 185454
rect 262582 185218 262614 185454
rect 261994 185134 262614 185218
rect 261994 184898 262026 185134
rect 262262 184898 262346 185134
rect 262582 184898 262614 185134
rect 261994 158454 262614 184898
rect 261994 158218 262026 158454
rect 262262 158218 262346 158454
rect 262582 158218 262614 158454
rect 261994 158134 262614 158218
rect 261994 157898 262026 158134
rect 262262 157898 262346 158134
rect 262582 157898 262614 158134
rect 261994 131454 262614 157898
rect 261994 131218 262026 131454
rect 262262 131218 262346 131454
rect 262582 131218 262614 131454
rect 261994 131134 262614 131218
rect 261994 130898 262026 131134
rect 262262 130898 262346 131134
rect 262582 130898 262614 131134
rect 261994 104454 262614 130898
rect 261994 104218 262026 104454
rect 262262 104218 262346 104454
rect 262582 104218 262614 104454
rect 261994 104134 262614 104218
rect 261994 103898 262026 104134
rect 262262 103898 262346 104134
rect 262582 103898 262614 104134
rect 261994 77454 262614 103898
rect 261994 77218 262026 77454
rect 262262 77218 262346 77454
rect 262582 77218 262614 77454
rect 261994 77134 262614 77218
rect 261994 76898 262026 77134
rect 262262 76898 262346 77134
rect 262582 76898 262614 77134
rect 261994 69000 262614 76898
rect 265494 704838 266114 711590
rect 265494 704602 265526 704838
rect 265762 704602 265846 704838
rect 266082 704602 266114 704838
rect 265494 704518 266114 704602
rect 265494 704282 265526 704518
rect 265762 704282 265846 704518
rect 266082 704282 266114 704518
rect 265494 701829 266114 704282
rect 265494 701593 265526 701829
rect 265762 701593 265846 701829
rect 266082 701593 266114 701829
rect 265494 701509 266114 701593
rect 265494 701273 265526 701509
rect 265762 701273 265846 701509
rect 266082 701273 266114 701509
rect 265494 674829 266114 701273
rect 265494 674593 265526 674829
rect 265762 674593 265846 674829
rect 266082 674593 266114 674829
rect 265494 674509 266114 674593
rect 265494 674273 265526 674509
rect 265762 674273 265846 674509
rect 266082 674273 266114 674509
rect 265494 647829 266114 674273
rect 265494 647593 265526 647829
rect 265762 647593 265846 647829
rect 266082 647593 266114 647829
rect 265494 647509 266114 647593
rect 265494 647273 265526 647509
rect 265762 647273 265846 647509
rect 266082 647273 266114 647509
rect 265494 620829 266114 647273
rect 265494 620593 265526 620829
rect 265762 620593 265846 620829
rect 266082 620593 266114 620829
rect 265494 620509 266114 620593
rect 265494 620273 265526 620509
rect 265762 620273 265846 620509
rect 266082 620273 266114 620509
rect 265494 593829 266114 620273
rect 265494 593593 265526 593829
rect 265762 593593 265846 593829
rect 266082 593593 266114 593829
rect 265494 593509 266114 593593
rect 265494 593273 265526 593509
rect 265762 593273 265846 593509
rect 266082 593273 266114 593509
rect 265494 566829 266114 593273
rect 265494 566593 265526 566829
rect 265762 566593 265846 566829
rect 266082 566593 266114 566829
rect 265494 566509 266114 566593
rect 265494 566273 265526 566509
rect 265762 566273 265846 566509
rect 266082 566273 266114 566509
rect 265494 539829 266114 566273
rect 265494 539593 265526 539829
rect 265762 539593 265846 539829
rect 266082 539593 266114 539829
rect 265494 539509 266114 539593
rect 265494 539273 265526 539509
rect 265762 539273 265846 539509
rect 266082 539273 266114 539509
rect 265494 512829 266114 539273
rect 265494 512593 265526 512829
rect 265762 512593 265846 512829
rect 266082 512593 266114 512829
rect 265494 512509 266114 512593
rect 265494 512273 265526 512509
rect 265762 512273 265846 512509
rect 266082 512273 266114 512509
rect 265494 485829 266114 512273
rect 265494 485593 265526 485829
rect 265762 485593 265846 485829
rect 266082 485593 266114 485829
rect 265494 485509 266114 485593
rect 265494 485273 265526 485509
rect 265762 485273 265846 485509
rect 266082 485273 266114 485509
rect 265494 458829 266114 485273
rect 265494 458593 265526 458829
rect 265762 458593 265846 458829
rect 266082 458593 266114 458829
rect 265494 458509 266114 458593
rect 265494 458273 265526 458509
rect 265762 458273 265846 458509
rect 266082 458273 266114 458509
rect 265494 431829 266114 458273
rect 265494 431593 265526 431829
rect 265762 431593 265846 431829
rect 266082 431593 266114 431829
rect 265494 431509 266114 431593
rect 265494 431273 265526 431509
rect 265762 431273 265846 431509
rect 266082 431273 266114 431509
rect 265494 404829 266114 431273
rect 265494 404593 265526 404829
rect 265762 404593 265846 404829
rect 266082 404593 266114 404829
rect 265494 404509 266114 404593
rect 265494 404273 265526 404509
rect 265762 404273 265846 404509
rect 266082 404273 266114 404509
rect 265494 377829 266114 404273
rect 265494 377593 265526 377829
rect 265762 377593 265846 377829
rect 266082 377593 266114 377829
rect 265494 377509 266114 377593
rect 265494 377273 265526 377509
rect 265762 377273 265846 377509
rect 266082 377273 266114 377509
rect 265494 350829 266114 377273
rect 265494 350593 265526 350829
rect 265762 350593 265846 350829
rect 266082 350593 266114 350829
rect 265494 350509 266114 350593
rect 265494 350273 265526 350509
rect 265762 350273 265846 350509
rect 266082 350273 266114 350509
rect 265494 323829 266114 350273
rect 265494 323593 265526 323829
rect 265762 323593 265846 323829
rect 266082 323593 266114 323829
rect 265494 323509 266114 323593
rect 265494 323273 265526 323509
rect 265762 323273 265846 323509
rect 266082 323273 266114 323509
rect 265494 296829 266114 323273
rect 265494 296593 265526 296829
rect 265762 296593 265846 296829
rect 266082 296593 266114 296829
rect 265494 296509 266114 296593
rect 265494 296273 265526 296509
rect 265762 296273 265846 296509
rect 266082 296273 266114 296509
rect 265494 269829 266114 296273
rect 265494 269593 265526 269829
rect 265762 269593 265846 269829
rect 266082 269593 266114 269829
rect 265494 269509 266114 269593
rect 265494 269273 265526 269509
rect 265762 269273 265846 269509
rect 266082 269273 266114 269509
rect 265494 242829 266114 269273
rect 265494 242593 265526 242829
rect 265762 242593 265846 242829
rect 266082 242593 266114 242829
rect 265494 242509 266114 242593
rect 265494 242273 265526 242509
rect 265762 242273 265846 242509
rect 266082 242273 266114 242509
rect 265494 215829 266114 242273
rect 265494 215593 265526 215829
rect 265762 215593 265846 215829
rect 266082 215593 266114 215829
rect 265494 215509 266114 215593
rect 265494 215273 265526 215509
rect 265762 215273 265846 215509
rect 266082 215273 266114 215509
rect 265494 188829 266114 215273
rect 265494 188593 265526 188829
rect 265762 188593 265846 188829
rect 266082 188593 266114 188829
rect 265494 188509 266114 188593
rect 265494 188273 265526 188509
rect 265762 188273 265846 188509
rect 266082 188273 266114 188509
rect 265494 161829 266114 188273
rect 265494 161593 265526 161829
rect 265762 161593 265846 161829
rect 266082 161593 266114 161829
rect 265494 161509 266114 161593
rect 265494 161273 265526 161509
rect 265762 161273 265846 161509
rect 266082 161273 266114 161509
rect 265494 134829 266114 161273
rect 265494 134593 265526 134829
rect 265762 134593 265846 134829
rect 266082 134593 266114 134829
rect 265494 134509 266114 134593
rect 265494 134273 265526 134509
rect 265762 134273 265846 134509
rect 266082 134273 266114 134509
rect 265494 107829 266114 134273
rect 265494 107593 265526 107829
rect 265762 107593 265846 107829
rect 266082 107593 266114 107829
rect 265494 107509 266114 107593
rect 265494 107273 265526 107509
rect 265762 107273 265846 107509
rect 266082 107273 266114 107509
rect 265494 80829 266114 107273
rect 265494 80593 265526 80829
rect 265762 80593 265846 80829
rect 266082 80593 266114 80829
rect 265494 80509 266114 80593
rect 265494 80273 265526 80509
rect 265762 80273 265846 80509
rect 266082 80273 266114 80509
rect 265494 69000 266114 80273
rect 289994 705798 290614 711590
rect 289994 705562 290026 705798
rect 290262 705562 290346 705798
rect 290582 705562 290614 705798
rect 289994 705478 290614 705562
rect 289994 705242 290026 705478
rect 290262 705242 290346 705478
rect 290582 705242 290614 705478
rect 289994 698454 290614 705242
rect 289994 698218 290026 698454
rect 290262 698218 290346 698454
rect 290582 698218 290614 698454
rect 289994 698134 290614 698218
rect 289994 697898 290026 698134
rect 290262 697898 290346 698134
rect 290582 697898 290614 698134
rect 289994 671454 290614 697898
rect 289994 671218 290026 671454
rect 290262 671218 290346 671454
rect 290582 671218 290614 671454
rect 289994 671134 290614 671218
rect 289994 670898 290026 671134
rect 290262 670898 290346 671134
rect 290582 670898 290614 671134
rect 289994 644454 290614 670898
rect 289994 644218 290026 644454
rect 290262 644218 290346 644454
rect 290582 644218 290614 644454
rect 289994 644134 290614 644218
rect 289994 643898 290026 644134
rect 290262 643898 290346 644134
rect 290582 643898 290614 644134
rect 289994 617454 290614 643898
rect 289994 617218 290026 617454
rect 290262 617218 290346 617454
rect 290582 617218 290614 617454
rect 289994 617134 290614 617218
rect 289994 616898 290026 617134
rect 290262 616898 290346 617134
rect 290582 616898 290614 617134
rect 289994 590454 290614 616898
rect 289994 590218 290026 590454
rect 290262 590218 290346 590454
rect 290582 590218 290614 590454
rect 289994 590134 290614 590218
rect 289994 589898 290026 590134
rect 290262 589898 290346 590134
rect 290582 589898 290614 590134
rect 289994 563454 290614 589898
rect 289994 563218 290026 563454
rect 290262 563218 290346 563454
rect 290582 563218 290614 563454
rect 289994 563134 290614 563218
rect 289994 562898 290026 563134
rect 290262 562898 290346 563134
rect 290582 562898 290614 563134
rect 289994 536454 290614 562898
rect 289994 536218 290026 536454
rect 290262 536218 290346 536454
rect 290582 536218 290614 536454
rect 289994 536134 290614 536218
rect 289994 535898 290026 536134
rect 290262 535898 290346 536134
rect 290582 535898 290614 536134
rect 289994 509454 290614 535898
rect 289994 509218 290026 509454
rect 290262 509218 290346 509454
rect 290582 509218 290614 509454
rect 289994 509134 290614 509218
rect 289994 508898 290026 509134
rect 290262 508898 290346 509134
rect 290582 508898 290614 509134
rect 289994 482454 290614 508898
rect 289994 482218 290026 482454
rect 290262 482218 290346 482454
rect 290582 482218 290614 482454
rect 289994 482134 290614 482218
rect 289994 481898 290026 482134
rect 290262 481898 290346 482134
rect 290582 481898 290614 482134
rect 289994 455454 290614 481898
rect 289994 455218 290026 455454
rect 290262 455218 290346 455454
rect 290582 455218 290614 455454
rect 289994 455134 290614 455218
rect 289994 454898 290026 455134
rect 290262 454898 290346 455134
rect 290582 454898 290614 455134
rect 289994 428454 290614 454898
rect 289994 428218 290026 428454
rect 290262 428218 290346 428454
rect 290582 428218 290614 428454
rect 289994 428134 290614 428218
rect 289994 427898 290026 428134
rect 290262 427898 290346 428134
rect 290582 427898 290614 428134
rect 289994 401454 290614 427898
rect 289994 401218 290026 401454
rect 290262 401218 290346 401454
rect 290582 401218 290614 401454
rect 289994 401134 290614 401218
rect 289994 400898 290026 401134
rect 290262 400898 290346 401134
rect 290582 400898 290614 401134
rect 289994 374454 290614 400898
rect 289994 374218 290026 374454
rect 290262 374218 290346 374454
rect 290582 374218 290614 374454
rect 289994 374134 290614 374218
rect 289994 373898 290026 374134
rect 290262 373898 290346 374134
rect 290582 373898 290614 374134
rect 289994 347454 290614 373898
rect 289994 347218 290026 347454
rect 290262 347218 290346 347454
rect 290582 347218 290614 347454
rect 289994 347134 290614 347218
rect 289994 346898 290026 347134
rect 290262 346898 290346 347134
rect 290582 346898 290614 347134
rect 289994 320454 290614 346898
rect 289994 320218 290026 320454
rect 290262 320218 290346 320454
rect 290582 320218 290614 320454
rect 289994 320134 290614 320218
rect 289994 319898 290026 320134
rect 290262 319898 290346 320134
rect 290582 319898 290614 320134
rect 289994 293454 290614 319898
rect 289994 293218 290026 293454
rect 290262 293218 290346 293454
rect 290582 293218 290614 293454
rect 289994 293134 290614 293218
rect 289994 292898 290026 293134
rect 290262 292898 290346 293134
rect 290582 292898 290614 293134
rect 289994 266454 290614 292898
rect 289994 266218 290026 266454
rect 290262 266218 290346 266454
rect 290582 266218 290614 266454
rect 289994 266134 290614 266218
rect 289994 265898 290026 266134
rect 290262 265898 290346 266134
rect 290582 265898 290614 266134
rect 289994 239454 290614 265898
rect 289994 239218 290026 239454
rect 290262 239218 290346 239454
rect 290582 239218 290614 239454
rect 289994 239134 290614 239218
rect 289994 238898 290026 239134
rect 290262 238898 290346 239134
rect 290582 238898 290614 239134
rect 289994 212454 290614 238898
rect 289994 212218 290026 212454
rect 290262 212218 290346 212454
rect 290582 212218 290614 212454
rect 289994 212134 290614 212218
rect 289994 211898 290026 212134
rect 290262 211898 290346 212134
rect 290582 211898 290614 212134
rect 289994 185454 290614 211898
rect 289994 185218 290026 185454
rect 290262 185218 290346 185454
rect 290582 185218 290614 185454
rect 289994 185134 290614 185218
rect 289994 184898 290026 185134
rect 290262 184898 290346 185134
rect 290582 184898 290614 185134
rect 289994 158454 290614 184898
rect 289994 158218 290026 158454
rect 290262 158218 290346 158454
rect 290582 158218 290614 158454
rect 289994 158134 290614 158218
rect 289994 157898 290026 158134
rect 290262 157898 290346 158134
rect 290582 157898 290614 158134
rect 289994 131454 290614 157898
rect 289994 131218 290026 131454
rect 290262 131218 290346 131454
rect 290582 131218 290614 131454
rect 289994 131134 290614 131218
rect 289994 130898 290026 131134
rect 290262 130898 290346 131134
rect 290582 130898 290614 131134
rect 289994 104454 290614 130898
rect 289994 104218 290026 104454
rect 290262 104218 290346 104454
rect 290582 104218 290614 104454
rect 289994 104134 290614 104218
rect 289994 103898 290026 104134
rect 290262 103898 290346 104134
rect 290582 103898 290614 104134
rect 289994 77454 290614 103898
rect 289994 77218 290026 77454
rect 290262 77218 290346 77454
rect 290582 77218 290614 77454
rect 289994 77134 290614 77218
rect 289994 76898 290026 77134
rect 290262 76898 290346 77134
rect 290582 76898 290614 77134
rect 289994 69000 290614 76898
rect 293494 704838 294114 711590
rect 293494 704602 293526 704838
rect 293762 704602 293846 704838
rect 294082 704602 294114 704838
rect 293494 704518 294114 704602
rect 293494 704282 293526 704518
rect 293762 704282 293846 704518
rect 294082 704282 294114 704518
rect 293494 701829 294114 704282
rect 293494 701593 293526 701829
rect 293762 701593 293846 701829
rect 294082 701593 294114 701829
rect 293494 701509 294114 701593
rect 293494 701273 293526 701509
rect 293762 701273 293846 701509
rect 294082 701273 294114 701509
rect 293494 674829 294114 701273
rect 293494 674593 293526 674829
rect 293762 674593 293846 674829
rect 294082 674593 294114 674829
rect 293494 674509 294114 674593
rect 293494 674273 293526 674509
rect 293762 674273 293846 674509
rect 294082 674273 294114 674509
rect 293494 647829 294114 674273
rect 293494 647593 293526 647829
rect 293762 647593 293846 647829
rect 294082 647593 294114 647829
rect 293494 647509 294114 647593
rect 293494 647273 293526 647509
rect 293762 647273 293846 647509
rect 294082 647273 294114 647509
rect 293494 620829 294114 647273
rect 293494 620593 293526 620829
rect 293762 620593 293846 620829
rect 294082 620593 294114 620829
rect 293494 620509 294114 620593
rect 293494 620273 293526 620509
rect 293762 620273 293846 620509
rect 294082 620273 294114 620509
rect 293494 593829 294114 620273
rect 293494 593593 293526 593829
rect 293762 593593 293846 593829
rect 294082 593593 294114 593829
rect 293494 593509 294114 593593
rect 293494 593273 293526 593509
rect 293762 593273 293846 593509
rect 294082 593273 294114 593509
rect 293494 566829 294114 593273
rect 293494 566593 293526 566829
rect 293762 566593 293846 566829
rect 294082 566593 294114 566829
rect 293494 566509 294114 566593
rect 293494 566273 293526 566509
rect 293762 566273 293846 566509
rect 294082 566273 294114 566509
rect 293494 539829 294114 566273
rect 293494 539593 293526 539829
rect 293762 539593 293846 539829
rect 294082 539593 294114 539829
rect 293494 539509 294114 539593
rect 293494 539273 293526 539509
rect 293762 539273 293846 539509
rect 294082 539273 294114 539509
rect 293494 512829 294114 539273
rect 293494 512593 293526 512829
rect 293762 512593 293846 512829
rect 294082 512593 294114 512829
rect 293494 512509 294114 512593
rect 293494 512273 293526 512509
rect 293762 512273 293846 512509
rect 294082 512273 294114 512509
rect 293494 485829 294114 512273
rect 293494 485593 293526 485829
rect 293762 485593 293846 485829
rect 294082 485593 294114 485829
rect 293494 485509 294114 485593
rect 293494 485273 293526 485509
rect 293762 485273 293846 485509
rect 294082 485273 294114 485509
rect 293494 458829 294114 485273
rect 293494 458593 293526 458829
rect 293762 458593 293846 458829
rect 294082 458593 294114 458829
rect 293494 458509 294114 458593
rect 293494 458273 293526 458509
rect 293762 458273 293846 458509
rect 294082 458273 294114 458509
rect 293494 431829 294114 458273
rect 293494 431593 293526 431829
rect 293762 431593 293846 431829
rect 294082 431593 294114 431829
rect 293494 431509 294114 431593
rect 293494 431273 293526 431509
rect 293762 431273 293846 431509
rect 294082 431273 294114 431509
rect 293494 404829 294114 431273
rect 293494 404593 293526 404829
rect 293762 404593 293846 404829
rect 294082 404593 294114 404829
rect 293494 404509 294114 404593
rect 293494 404273 293526 404509
rect 293762 404273 293846 404509
rect 294082 404273 294114 404509
rect 293494 377829 294114 404273
rect 293494 377593 293526 377829
rect 293762 377593 293846 377829
rect 294082 377593 294114 377829
rect 293494 377509 294114 377593
rect 293494 377273 293526 377509
rect 293762 377273 293846 377509
rect 294082 377273 294114 377509
rect 293494 350829 294114 377273
rect 293494 350593 293526 350829
rect 293762 350593 293846 350829
rect 294082 350593 294114 350829
rect 293494 350509 294114 350593
rect 293494 350273 293526 350509
rect 293762 350273 293846 350509
rect 294082 350273 294114 350509
rect 293494 323829 294114 350273
rect 293494 323593 293526 323829
rect 293762 323593 293846 323829
rect 294082 323593 294114 323829
rect 293494 323509 294114 323593
rect 293494 323273 293526 323509
rect 293762 323273 293846 323509
rect 294082 323273 294114 323509
rect 293494 296829 294114 323273
rect 293494 296593 293526 296829
rect 293762 296593 293846 296829
rect 294082 296593 294114 296829
rect 293494 296509 294114 296593
rect 293494 296273 293526 296509
rect 293762 296273 293846 296509
rect 294082 296273 294114 296509
rect 293494 269829 294114 296273
rect 293494 269593 293526 269829
rect 293762 269593 293846 269829
rect 294082 269593 294114 269829
rect 293494 269509 294114 269593
rect 293494 269273 293526 269509
rect 293762 269273 293846 269509
rect 294082 269273 294114 269509
rect 293494 242829 294114 269273
rect 293494 242593 293526 242829
rect 293762 242593 293846 242829
rect 294082 242593 294114 242829
rect 293494 242509 294114 242593
rect 293494 242273 293526 242509
rect 293762 242273 293846 242509
rect 294082 242273 294114 242509
rect 293494 215829 294114 242273
rect 293494 215593 293526 215829
rect 293762 215593 293846 215829
rect 294082 215593 294114 215829
rect 293494 215509 294114 215593
rect 293494 215273 293526 215509
rect 293762 215273 293846 215509
rect 294082 215273 294114 215509
rect 293494 188829 294114 215273
rect 293494 188593 293526 188829
rect 293762 188593 293846 188829
rect 294082 188593 294114 188829
rect 293494 188509 294114 188593
rect 293494 188273 293526 188509
rect 293762 188273 293846 188509
rect 294082 188273 294114 188509
rect 293494 161829 294114 188273
rect 293494 161593 293526 161829
rect 293762 161593 293846 161829
rect 294082 161593 294114 161829
rect 293494 161509 294114 161593
rect 293494 161273 293526 161509
rect 293762 161273 293846 161509
rect 294082 161273 294114 161509
rect 293494 134829 294114 161273
rect 293494 134593 293526 134829
rect 293762 134593 293846 134829
rect 294082 134593 294114 134829
rect 293494 134509 294114 134593
rect 293494 134273 293526 134509
rect 293762 134273 293846 134509
rect 294082 134273 294114 134509
rect 293494 107829 294114 134273
rect 293494 107593 293526 107829
rect 293762 107593 293846 107829
rect 294082 107593 294114 107829
rect 293494 107509 294114 107593
rect 293494 107273 293526 107509
rect 293762 107273 293846 107509
rect 294082 107273 294114 107509
rect 293494 80829 294114 107273
rect 293494 80593 293526 80829
rect 293762 80593 293846 80829
rect 294082 80593 294114 80829
rect 293494 80509 294114 80593
rect 293494 80273 293526 80509
rect 293762 80273 293846 80509
rect 294082 80273 294114 80509
rect 293494 69000 294114 80273
rect 317994 705798 318614 711590
rect 317994 705562 318026 705798
rect 318262 705562 318346 705798
rect 318582 705562 318614 705798
rect 317994 705478 318614 705562
rect 317994 705242 318026 705478
rect 318262 705242 318346 705478
rect 318582 705242 318614 705478
rect 317994 698454 318614 705242
rect 317994 698218 318026 698454
rect 318262 698218 318346 698454
rect 318582 698218 318614 698454
rect 317994 698134 318614 698218
rect 317994 697898 318026 698134
rect 318262 697898 318346 698134
rect 318582 697898 318614 698134
rect 317994 671454 318614 697898
rect 317994 671218 318026 671454
rect 318262 671218 318346 671454
rect 318582 671218 318614 671454
rect 317994 671134 318614 671218
rect 317994 670898 318026 671134
rect 318262 670898 318346 671134
rect 318582 670898 318614 671134
rect 317994 644454 318614 670898
rect 317994 644218 318026 644454
rect 318262 644218 318346 644454
rect 318582 644218 318614 644454
rect 317994 644134 318614 644218
rect 317994 643898 318026 644134
rect 318262 643898 318346 644134
rect 318582 643898 318614 644134
rect 317994 617454 318614 643898
rect 317994 617218 318026 617454
rect 318262 617218 318346 617454
rect 318582 617218 318614 617454
rect 317994 617134 318614 617218
rect 317994 616898 318026 617134
rect 318262 616898 318346 617134
rect 318582 616898 318614 617134
rect 317994 590454 318614 616898
rect 317994 590218 318026 590454
rect 318262 590218 318346 590454
rect 318582 590218 318614 590454
rect 317994 590134 318614 590218
rect 317994 589898 318026 590134
rect 318262 589898 318346 590134
rect 318582 589898 318614 590134
rect 317994 563454 318614 589898
rect 317994 563218 318026 563454
rect 318262 563218 318346 563454
rect 318582 563218 318614 563454
rect 317994 563134 318614 563218
rect 317994 562898 318026 563134
rect 318262 562898 318346 563134
rect 318582 562898 318614 563134
rect 317994 536454 318614 562898
rect 317994 536218 318026 536454
rect 318262 536218 318346 536454
rect 318582 536218 318614 536454
rect 317994 536134 318614 536218
rect 317994 535898 318026 536134
rect 318262 535898 318346 536134
rect 318582 535898 318614 536134
rect 317994 509454 318614 535898
rect 317994 509218 318026 509454
rect 318262 509218 318346 509454
rect 318582 509218 318614 509454
rect 317994 509134 318614 509218
rect 317994 508898 318026 509134
rect 318262 508898 318346 509134
rect 318582 508898 318614 509134
rect 317994 482454 318614 508898
rect 317994 482218 318026 482454
rect 318262 482218 318346 482454
rect 318582 482218 318614 482454
rect 317994 482134 318614 482218
rect 317994 481898 318026 482134
rect 318262 481898 318346 482134
rect 318582 481898 318614 482134
rect 317994 455454 318614 481898
rect 317994 455218 318026 455454
rect 318262 455218 318346 455454
rect 318582 455218 318614 455454
rect 317994 455134 318614 455218
rect 317994 454898 318026 455134
rect 318262 454898 318346 455134
rect 318582 454898 318614 455134
rect 317994 428454 318614 454898
rect 317994 428218 318026 428454
rect 318262 428218 318346 428454
rect 318582 428218 318614 428454
rect 317994 428134 318614 428218
rect 317994 427898 318026 428134
rect 318262 427898 318346 428134
rect 318582 427898 318614 428134
rect 317994 401454 318614 427898
rect 317994 401218 318026 401454
rect 318262 401218 318346 401454
rect 318582 401218 318614 401454
rect 317994 401134 318614 401218
rect 317994 400898 318026 401134
rect 318262 400898 318346 401134
rect 318582 400898 318614 401134
rect 317994 374454 318614 400898
rect 317994 374218 318026 374454
rect 318262 374218 318346 374454
rect 318582 374218 318614 374454
rect 317994 374134 318614 374218
rect 317994 373898 318026 374134
rect 318262 373898 318346 374134
rect 318582 373898 318614 374134
rect 317994 347454 318614 373898
rect 317994 347218 318026 347454
rect 318262 347218 318346 347454
rect 318582 347218 318614 347454
rect 317994 347134 318614 347218
rect 317994 346898 318026 347134
rect 318262 346898 318346 347134
rect 318582 346898 318614 347134
rect 317994 320454 318614 346898
rect 317994 320218 318026 320454
rect 318262 320218 318346 320454
rect 318582 320218 318614 320454
rect 317994 320134 318614 320218
rect 317994 319898 318026 320134
rect 318262 319898 318346 320134
rect 318582 319898 318614 320134
rect 317994 293454 318614 319898
rect 317994 293218 318026 293454
rect 318262 293218 318346 293454
rect 318582 293218 318614 293454
rect 317994 293134 318614 293218
rect 317994 292898 318026 293134
rect 318262 292898 318346 293134
rect 318582 292898 318614 293134
rect 317994 266454 318614 292898
rect 317994 266218 318026 266454
rect 318262 266218 318346 266454
rect 318582 266218 318614 266454
rect 317994 266134 318614 266218
rect 317994 265898 318026 266134
rect 318262 265898 318346 266134
rect 318582 265898 318614 266134
rect 317994 239454 318614 265898
rect 317994 239218 318026 239454
rect 318262 239218 318346 239454
rect 318582 239218 318614 239454
rect 317994 239134 318614 239218
rect 317994 238898 318026 239134
rect 318262 238898 318346 239134
rect 318582 238898 318614 239134
rect 317994 212454 318614 238898
rect 317994 212218 318026 212454
rect 318262 212218 318346 212454
rect 318582 212218 318614 212454
rect 317994 212134 318614 212218
rect 317994 211898 318026 212134
rect 318262 211898 318346 212134
rect 318582 211898 318614 212134
rect 317994 185454 318614 211898
rect 317994 185218 318026 185454
rect 318262 185218 318346 185454
rect 318582 185218 318614 185454
rect 317994 185134 318614 185218
rect 317994 184898 318026 185134
rect 318262 184898 318346 185134
rect 318582 184898 318614 185134
rect 317994 158454 318614 184898
rect 317994 158218 318026 158454
rect 318262 158218 318346 158454
rect 318582 158218 318614 158454
rect 317994 158134 318614 158218
rect 317994 157898 318026 158134
rect 318262 157898 318346 158134
rect 318582 157898 318614 158134
rect 317994 131454 318614 157898
rect 317994 131218 318026 131454
rect 318262 131218 318346 131454
rect 318582 131218 318614 131454
rect 317994 131134 318614 131218
rect 317994 130898 318026 131134
rect 318262 130898 318346 131134
rect 318582 130898 318614 131134
rect 317994 104454 318614 130898
rect 317994 104218 318026 104454
rect 318262 104218 318346 104454
rect 318582 104218 318614 104454
rect 317994 104134 318614 104218
rect 317994 103898 318026 104134
rect 318262 103898 318346 104134
rect 318582 103898 318614 104134
rect 317994 77454 318614 103898
rect 317994 77218 318026 77454
rect 318262 77218 318346 77454
rect 318582 77218 318614 77454
rect 317994 77134 318614 77218
rect 317994 76898 318026 77134
rect 318262 76898 318346 77134
rect 318582 76898 318614 77134
rect 317994 69000 318614 76898
rect 321494 704838 322114 711590
rect 321494 704602 321526 704838
rect 321762 704602 321846 704838
rect 322082 704602 322114 704838
rect 321494 704518 322114 704602
rect 321494 704282 321526 704518
rect 321762 704282 321846 704518
rect 322082 704282 322114 704518
rect 321494 701829 322114 704282
rect 321494 701593 321526 701829
rect 321762 701593 321846 701829
rect 322082 701593 322114 701829
rect 321494 701509 322114 701593
rect 321494 701273 321526 701509
rect 321762 701273 321846 701509
rect 322082 701273 322114 701509
rect 321494 674829 322114 701273
rect 321494 674593 321526 674829
rect 321762 674593 321846 674829
rect 322082 674593 322114 674829
rect 321494 674509 322114 674593
rect 321494 674273 321526 674509
rect 321762 674273 321846 674509
rect 322082 674273 322114 674509
rect 321494 647829 322114 674273
rect 321494 647593 321526 647829
rect 321762 647593 321846 647829
rect 322082 647593 322114 647829
rect 321494 647509 322114 647593
rect 321494 647273 321526 647509
rect 321762 647273 321846 647509
rect 322082 647273 322114 647509
rect 321494 620829 322114 647273
rect 321494 620593 321526 620829
rect 321762 620593 321846 620829
rect 322082 620593 322114 620829
rect 321494 620509 322114 620593
rect 321494 620273 321526 620509
rect 321762 620273 321846 620509
rect 322082 620273 322114 620509
rect 321494 593829 322114 620273
rect 321494 593593 321526 593829
rect 321762 593593 321846 593829
rect 322082 593593 322114 593829
rect 321494 593509 322114 593593
rect 321494 593273 321526 593509
rect 321762 593273 321846 593509
rect 322082 593273 322114 593509
rect 321494 566829 322114 593273
rect 321494 566593 321526 566829
rect 321762 566593 321846 566829
rect 322082 566593 322114 566829
rect 321494 566509 322114 566593
rect 321494 566273 321526 566509
rect 321762 566273 321846 566509
rect 322082 566273 322114 566509
rect 321494 539829 322114 566273
rect 321494 539593 321526 539829
rect 321762 539593 321846 539829
rect 322082 539593 322114 539829
rect 321494 539509 322114 539593
rect 321494 539273 321526 539509
rect 321762 539273 321846 539509
rect 322082 539273 322114 539509
rect 321494 512829 322114 539273
rect 321494 512593 321526 512829
rect 321762 512593 321846 512829
rect 322082 512593 322114 512829
rect 321494 512509 322114 512593
rect 321494 512273 321526 512509
rect 321762 512273 321846 512509
rect 322082 512273 322114 512509
rect 321494 485829 322114 512273
rect 321494 485593 321526 485829
rect 321762 485593 321846 485829
rect 322082 485593 322114 485829
rect 321494 485509 322114 485593
rect 321494 485273 321526 485509
rect 321762 485273 321846 485509
rect 322082 485273 322114 485509
rect 321494 458829 322114 485273
rect 321494 458593 321526 458829
rect 321762 458593 321846 458829
rect 322082 458593 322114 458829
rect 321494 458509 322114 458593
rect 321494 458273 321526 458509
rect 321762 458273 321846 458509
rect 322082 458273 322114 458509
rect 321494 431829 322114 458273
rect 321494 431593 321526 431829
rect 321762 431593 321846 431829
rect 322082 431593 322114 431829
rect 321494 431509 322114 431593
rect 321494 431273 321526 431509
rect 321762 431273 321846 431509
rect 322082 431273 322114 431509
rect 321494 404829 322114 431273
rect 321494 404593 321526 404829
rect 321762 404593 321846 404829
rect 322082 404593 322114 404829
rect 321494 404509 322114 404593
rect 321494 404273 321526 404509
rect 321762 404273 321846 404509
rect 322082 404273 322114 404509
rect 321494 377829 322114 404273
rect 321494 377593 321526 377829
rect 321762 377593 321846 377829
rect 322082 377593 322114 377829
rect 321494 377509 322114 377593
rect 321494 377273 321526 377509
rect 321762 377273 321846 377509
rect 322082 377273 322114 377509
rect 321494 350829 322114 377273
rect 321494 350593 321526 350829
rect 321762 350593 321846 350829
rect 322082 350593 322114 350829
rect 321494 350509 322114 350593
rect 321494 350273 321526 350509
rect 321762 350273 321846 350509
rect 322082 350273 322114 350509
rect 321494 323829 322114 350273
rect 321494 323593 321526 323829
rect 321762 323593 321846 323829
rect 322082 323593 322114 323829
rect 321494 323509 322114 323593
rect 321494 323273 321526 323509
rect 321762 323273 321846 323509
rect 322082 323273 322114 323509
rect 321494 296829 322114 323273
rect 321494 296593 321526 296829
rect 321762 296593 321846 296829
rect 322082 296593 322114 296829
rect 321494 296509 322114 296593
rect 321494 296273 321526 296509
rect 321762 296273 321846 296509
rect 322082 296273 322114 296509
rect 321494 269829 322114 296273
rect 321494 269593 321526 269829
rect 321762 269593 321846 269829
rect 322082 269593 322114 269829
rect 321494 269509 322114 269593
rect 321494 269273 321526 269509
rect 321762 269273 321846 269509
rect 322082 269273 322114 269509
rect 321494 242829 322114 269273
rect 321494 242593 321526 242829
rect 321762 242593 321846 242829
rect 322082 242593 322114 242829
rect 321494 242509 322114 242593
rect 321494 242273 321526 242509
rect 321762 242273 321846 242509
rect 322082 242273 322114 242509
rect 321494 215829 322114 242273
rect 321494 215593 321526 215829
rect 321762 215593 321846 215829
rect 322082 215593 322114 215829
rect 321494 215509 322114 215593
rect 321494 215273 321526 215509
rect 321762 215273 321846 215509
rect 322082 215273 322114 215509
rect 321494 188829 322114 215273
rect 321494 188593 321526 188829
rect 321762 188593 321846 188829
rect 322082 188593 322114 188829
rect 321494 188509 322114 188593
rect 321494 188273 321526 188509
rect 321762 188273 321846 188509
rect 322082 188273 322114 188509
rect 321494 161829 322114 188273
rect 321494 161593 321526 161829
rect 321762 161593 321846 161829
rect 322082 161593 322114 161829
rect 321494 161509 322114 161593
rect 321494 161273 321526 161509
rect 321762 161273 321846 161509
rect 322082 161273 322114 161509
rect 321494 134829 322114 161273
rect 321494 134593 321526 134829
rect 321762 134593 321846 134829
rect 322082 134593 322114 134829
rect 321494 134509 322114 134593
rect 321494 134273 321526 134509
rect 321762 134273 321846 134509
rect 322082 134273 322114 134509
rect 321494 107829 322114 134273
rect 321494 107593 321526 107829
rect 321762 107593 321846 107829
rect 322082 107593 322114 107829
rect 321494 107509 322114 107593
rect 321494 107273 321526 107509
rect 321762 107273 321846 107509
rect 322082 107273 322114 107509
rect 321494 80829 322114 107273
rect 321494 80593 321526 80829
rect 321762 80593 321846 80829
rect 322082 80593 322114 80829
rect 321494 80509 322114 80593
rect 321494 80273 321526 80509
rect 321762 80273 321846 80509
rect 322082 80273 322114 80509
rect 321494 69000 322114 80273
rect 345994 705798 346614 711590
rect 345994 705562 346026 705798
rect 346262 705562 346346 705798
rect 346582 705562 346614 705798
rect 345994 705478 346614 705562
rect 345994 705242 346026 705478
rect 346262 705242 346346 705478
rect 346582 705242 346614 705478
rect 345994 698454 346614 705242
rect 345994 698218 346026 698454
rect 346262 698218 346346 698454
rect 346582 698218 346614 698454
rect 345994 698134 346614 698218
rect 345994 697898 346026 698134
rect 346262 697898 346346 698134
rect 346582 697898 346614 698134
rect 345994 671454 346614 697898
rect 345994 671218 346026 671454
rect 346262 671218 346346 671454
rect 346582 671218 346614 671454
rect 345994 671134 346614 671218
rect 345994 670898 346026 671134
rect 346262 670898 346346 671134
rect 346582 670898 346614 671134
rect 345994 644454 346614 670898
rect 345994 644218 346026 644454
rect 346262 644218 346346 644454
rect 346582 644218 346614 644454
rect 345994 644134 346614 644218
rect 345994 643898 346026 644134
rect 346262 643898 346346 644134
rect 346582 643898 346614 644134
rect 345994 617454 346614 643898
rect 345994 617218 346026 617454
rect 346262 617218 346346 617454
rect 346582 617218 346614 617454
rect 345994 617134 346614 617218
rect 345994 616898 346026 617134
rect 346262 616898 346346 617134
rect 346582 616898 346614 617134
rect 345994 590454 346614 616898
rect 345994 590218 346026 590454
rect 346262 590218 346346 590454
rect 346582 590218 346614 590454
rect 345994 590134 346614 590218
rect 345994 589898 346026 590134
rect 346262 589898 346346 590134
rect 346582 589898 346614 590134
rect 345994 563454 346614 589898
rect 345994 563218 346026 563454
rect 346262 563218 346346 563454
rect 346582 563218 346614 563454
rect 345994 563134 346614 563218
rect 345994 562898 346026 563134
rect 346262 562898 346346 563134
rect 346582 562898 346614 563134
rect 345994 536454 346614 562898
rect 345994 536218 346026 536454
rect 346262 536218 346346 536454
rect 346582 536218 346614 536454
rect 345994 536134 346614 536218
rect 345994 535898 346026 536134
rect 346262 535898 346346 536134
rect 346582 535898 346614 536134
rect 345994 509454 346614 535898
rect 345994 509218 346026 509454
rect 346262 509218 346346 509454
rect 346582 509218 346614 509454
rect 345994 509134 346614 509218
rect 345994 508898 346026 509134
rect 346262 508898 346346 509134
rect 346582 508898 346614 509134
rect 345994 482454 346614 508898
rect 345994 482218 346026 482454
rect 346262 482218 346346 482454
rect 346582 482218 346614 482454
rect 345994 482134 346614 482218
rect 345994 481898 346026 482134
rect 346262 481898 346346 482134
rect 346582 481898 346614 482134
rect 345994 455454 346614 481898
rect 345994 455218 346026 455454
rect 346262 455218 346346 455454
rect 346582 455218 346614 455454
rect 345994 455134 346614 455218
rect 345994 454898 346026 455134
rect 346262 454898 346346 455134
rect 346582 454898 346614 455134
rect 345994 428454 346614 454898
rect 345994 428218 346026 428454
rect 346262 428218 346346 428454
rect 346582 428218 346614 428454
rect 345994 428134 346614 428218
rect 345994 427898 346026 428134
rect 346262 427898 346346 428134
rect 346582 427898 346614 428134
rect 345994 401454 346614 427898
rect 345994 401218 346026 401454
rect 346262 401218 346346 401454
rect 346582 401218 346614 401454
rect 345994 401134 346614 401218
rect 345994 400898 346026 401134
rect 346262 400898 346346 401134
rect 346582 400898 346614 401134
rect 345994 374454 346614 400898
rect 345994 374218 346026 374454
rect 346262 374218 346346 374454
rect 346582 374218 346614 374454
rect 345994 374134 346614 374218
rect 345994 373898 346026 374134
rect 346262 373898 346346 374134
rect 346582 373898 346614 374134
rect 345994 347454 346614 373898
rect 345994 347218 346026 347454
rect 346262 347218 346346 347454
rect 346582 347218 346614 347454
rect 345994 347134 346614 347218
rect 345994 346898 346026 347134
rect 346262 346898 346346 347134
rect 346582 346898 346614 347134
rect 345994 320454 346614 346898
rect 345994 320218 346026 320454
rect 346262 320218 346346 320454
rect 346582 320218 346614 320454
rect 345994 320134 346614 320218
rect 345994 319898 346026 320134
rect 346262 319898 346346 320134
rect 346582 319898 346614 320134
rect 345994 293454 346614 319898
rect 345994 293218 346026 293454
rect 346262 293218 346346 293454
rect 346582 293218 346614 293454
rect 345994 293134 346614 293218
rect 345994 292898 346026 293134
rect 346262 292898 346346 293134
rect 346582 292898 346614 293134
rect 345994 266454 346614 292898
rect 345994 266218 346026 266454
rect 346262 266218 346346 266454
rect 346582 266218 346614 266454
rect 345994 266134 346614 266218
rect 345994 265898 346026 266134
rect 346262 265898 346346 266134
rect 346582 265898 346614 266134
rect 345994 239454 346614 265898
rect 345994 239218 346026 239454
rect 346262 239218 346346 239454
rect 346582 239218 346614 239454
rect 345994 239134 346614 239218
rect 345994 238898 346026 239134
rect 346262 238898 346346 239134
rect 346582 238898 346614 239134
rect 345994 212454 346614 238898
rect 345994 212218 346026 212454
rect 346262 212218 346346 212454
rect 346582 212218 346614 212454
rect 345994 212134 346614 212218
rect 345994 211898 346026 212134
rect 346262 211898 346346 212134
rect 346582 211898 346614 212134
rect 345994 185454 346614 211898
rect 345994 185218 346026 185454
rect 346262 185218 346346 185454
rect 346582 185218 346614 185454
rect 345994 185134 346614 185218
rect 345994 184898 346026 185134
rect 346262 184898 346346 185134
rect 346582 184898 346614 185134
rect 345994 158454 346614 184898
rect 345994 158218 346026 158454
rect 346262 158218 346346 158454
rect 346582 158218 346614 158454
rect 345994 158134 346614 158218
rect 345994 157898 346026 158134
rect 346262 157898 346346 158134
rect 346582 157898 346614 158134
rect 345994 131454 346614 157898
rect 345994 131218 346026 131454
rect 346262 131218 346346 131454
rect 346582 131218 346614 131454
rect 345994 131134 346614 131218
rect 345994 130898 346026 131134
rect 346262 130898 346346 131134
rect 346582 130898 346614 131134
rect 345994 104454 346614 130898
rect 345994 104218 346026 104454
rect 346262 104218 346346 104454
rect 346582 104218 346614 104454
rect 345994 104134 346614 104218
rect 345994 103898 346026 104134
rect 346262 103898 346346 104134
rect 346582 103898 346614 104134
rect 345994 77454 346614 103898
rect 345994 77218 346026 77454
rect 346262 77218 346346 77454
rect 346582 77218 346614 77454
rect 345994 77134 346614 77218
rect 345994 76898 346026 77134
rect 346262 76898 346346 77134
rect 346582 76898 346614 77134
rect 345994 69000 346614 76898
rect 349494 704838 350114 711590
rect 349494 704602 349526 704838
rect 349762 704602 349846 704838
rect 350082 704602 350114 704838
rect 349494 704518 350114 704602
rect 349494 704282 349526 704518
rect 349762 704282 349846 704518
rect 350082 704282 350114 704518
rect 349494 701829 350114 704282
rect 349494 701593 349526 701829
rect 349762 701593 349846 701829
rect 350082 701593 350114 701829
rect 349494 701509 350114 701593
rect 349494 701273 349526 701509
rect 349762 701273 349846 701509
rect 350082 701273 350114 701509
rect 349494 674829 350114 701273
rect 349494 674593 349526 674829
rect 349762 674593 349846 674829
rect 350082 674593 350114 674829
rect 349494 674509 350114 674593
rect 349494 674273 349526 674509
rect 349762 674273 349846 674509
rect 350082 674273 350114 674509
rect 349494 647829 350114 674273
rect 349494 647593 349526 647829
rect 349762 647593 349846 647829
rect 350082 647593 350114 647829
rect 349494 647509 350114 647593
rect 349494 647273 349526 647509
rect 349762 647273 349846 647509
rect 350082 647273 350114 647509
rect 349494 620829 350114 647273
rect 349494 620593 349526 620829
rect 349762 620593 349846 620829
rect 350082 620593 350114 620829
rect 349494 620509 350114 620593
rect 349494 620273 349526 620509
rect 349762 620273 349846 620509
rect 350082 620273 350114 620509
rect 349494 593829 350114 620273
rect 349494 593593 349526 593829
rect 349762 593593 349846 593829
rect 350082 593593 350114 593829
rect 349494 593509 350114 593593
rect 349494 593273 349526 593509
rect 349762 593273 349846 593509
rect 350082 593273 350114 593509
rect 349494 566829 350114 593273
rect 349494 566593 349526 566829
rect 349762 566593 349846 566829
rect 350082 566593 350114 566829
rect 349494 566509 350114 566593
rect 349494 566273 349526 566509
rect 349762 566273 349846 566509
rect 350082 566273 350114 566509
rect 349494 539829 350114 566273
rect 349494 539593 349526 539829
rect 349762 539593 349846 539829
rect 350082 539593 350114 539829
rect 349494 539509 350114 539593
rect 349494 539273 349526 539509
rect 349762 539273 349846 539509
rect 350082 539273 350114 539509
rect 349494 512829 350114 539273
rect 349494 512593 349526 512829
rect 349762 512593 349846 512829
rect 350082 512593 350114 512829
rect 349494 512509 350114 512593
rect 349494 512273 349526 512509
rect 349762 512273 349846 512509
rect 350082 512273 350114 512509
rect 349494 485829 350114 512273
rect 349494 485593 349526 485829
rect 349762 485593 349846 485829
rect 350082 485593 350114 485829
rect 349494 485509 350114 485593
rect 349494 485273 349526 485509
rect 349762 485273 349846 485509
rect 350082 485273 350114 485509
rect 349494 458829 350114 485273
rect 349494 458593 349526 458829
rect 349762 458593 349846 458829
rect 350082 458593 350114 458829
rect 349494 458509 350114 458593
rect 349494 458273 349526 458509
rect 349762 458273 349846 458509
rect 350082 458273 350114 458509
rect 349494 431829 350114 458273
rect 349494 431593 349526 431829
rect 349762 431593 349846 431829
rect 350082 431593 350114 431829
rect 349494 431509 350114 431593
rect 349494 431273 349526 431509
rect 349762 431273 349846 431509
rect 350082 431273 350114 431509
rect 349494 404829 350114 431273
rect 349494 404593 349526 404829
rect 349762 404593 349846 404829
rect 350082 404593 350114 404829
rect 349494 404509 350114 404593
rect 349494 404273 349526 404509
rect 349762 404273 349846 404509
rect 350082 404273 350114 404509
rect 349494 377829 350114 404273
rect 349494 377593 349526 377829
rect 349762 377593 349846 377829
rect 350082 377593 350114 377829
rect 349494 377509 350114 377593
rect 349494 377273 349526 377509
rect 349762 377273 349846 377509
rect 350082 377273 350114 377509
rect 349494 350829 350114 377273
rect 349494 350593 349526 350829
rect 349762 350593 349846 350829
rect 350082 350593 350114 350829
rect 349494 350509 350114 350593
rect 349494 350273 349526 350509
rect 349762 350273 349846 350509
rect 350082 350273 350114 350509
rect 349494 323829 350114 350273
rect 349494 323593 349526 323829
rect 349762 323593 349846 323829
rect 350082 323593 350114 323829
rect 349494 323509 350114 323593
rect 349494 323273 349526 323509
rect 349762 323273 349846 323509
rect 350082 323273 350114 323509
rect 349494 296829 350114 323273
rect 349494 296593 349526 296829
rect 349762 296593 349846 296829
rect 350082 296593 350114 296829
rect 349494 296509 350114 296593
rect 349494 296273 349526 296509
rect 349762 296273 349846 296509
rect 350082 296273 350114 296509
rect 349494 269829 350114 296273
rect 349494 269593 349526 269829
rect 349762 269593 349846 269829
rect 350082 269593 350114 269829
rect 349494 269509 350114 269593
rect 349494 269273 349526 269509
rect 349762 269273 349846 269509
rect 350082 269273 350114 269509
rect 349494 242829 350114 269273
rect 349494 242593 349526 242829
rect 349762 242593 349846 242829
rect 350082 242593 350114 242829
rect 349494 242509 350114 242593
rect 349494 242273 349526 242509
rect 349762 242273 349846 242509
rect 350082 242273 350114 242509
rect 349494 215829 350114 242273
rect 349494 215593 349526 215829
rect 349762 215593 349846 215829
rect 350082 215593 350114 215829
rect 349494 215509 350114 215593
rect 349494 215273 349526 215509
rect 349762 215273 349846 215509
rect 350082 215273 350114 215509
rect 349494 188829 350114 215273
rect 349494 188593 349526 188829
rect 349762 188593 349846 188829
rect 350082 188593 350114 188829
rect 349494 188509 350114 188593
rect 349494 188273 349526 188509
rect 349762 188273 349846 188509
rect 350082 188273 350114 188509
rect 349494 161829 350114 188273
rect 349494 161593 349526 161829
rect 349762 161593 349846 161829
rect 350082 161593 350114 161829
rect 349494 161509 350114 161593
rect 349494 161273 349526 161509
rect 349762 161273 349846 161509
rect 350082 161273 350114 161509
rect 349494 134829 350114 161273
rect 349494 134593 349526 134829
rect 349762 134593 349846 134829
rect 350082 134593 350114 134829
rect 349494 134509 350114 134593
rect 349494 134273 349526 134509
rect 349762 134273 349846 134509
rect 350082 134273 350114 134509
rect 349494 107829 350114 134273
rect 349494 107593 349526 107829
rect 349762 107593 349846 107829
rect 350082 107593 350114 107829
rect 349494 107509 350114 107593
rect 349494 107273 349526 107509
rect 349762 107273 349846 107509
rect 350082 107273 350114 107509
rect 349494 80829 350114 107273
rect 349494 80593 349526 80829
rect 349762 80593 349846 80829
rect 350082 80593 350114 80829
rect 349494 80509 350114 80593
rect 349494 80273 349526 80509
rect 349762 80273 349846 80509
rect 350082 80273 350114 80509
rect 349494 69000 350114 80273
rect 373994 705798 374614 711590
rect 373994 705562 374026 705798
rect 374262 705562 374346 705798
rect 374582 705562 374614 705798
rect 373994 705478 374614 705562
rect 373994 705242 374026 705478
rect 374262 705242 374346 705478
rect 374582 705242 374614 705478
rect 373994 698454 374614 705242
rect 373994 698218 374026 698454
rect 374262 698218 374346 698454
rect 374582 698218 374614 698454
rect 373994 698134 374614 698218
rect 373994 697898 374026 698134
rect 374262 697898 374346 698134
rect 374582 697898 374614 698134
rect 373994 671454 374614 697898
rect 373994 671218 374026 671454
rect 374262 671218 374346 671454
rect 374582 671218 374614 671454
rect 373994 671134 374614 671218
rect 373994 670898 374026 671134
rect 374262 670898 374346 671134
rect 374582 670898 374614 671134
rect 373994 644454 374614 670898
rect 373994 644218 374026 644454
rect 374262 644218 374346 644454
rect 374582 644218 374614 644454
rect 373994 644134 374614 644218
rect 373994 643898 374026 644134
rect 374262 643898 374346 644134
rect 374582 643898 374614 644134
rect 373994 617454 374614 643898
rect 373994 617218 374026 617454
rect 374262 617218 374346 617454
rect 374582 617218 374614 617454
rect 373994 617134 374614 617218
rect 373994 616898 374026 617134
rect 374262 616898 374346 617134
rect 374582 616898 374614 617134
rect 373994 590454 374614 616898
rect 373994 590218 374026 590454
rect 374262 590218 374346 590454
rect 374582 590218 374614 590454
rect 373994 590134 374614 590218
rect 373994 589898 374026 590134
rect 374262 589898 374346 590134
rect 374582 589898 374614 590134
rect 373994 563454 374614 589898
rect 373994 563218 374026 563454
rect 374262 563218 374346 563454
rect 374582 563218 374614 563454
rect 373994 563134 374614 563218
rect 373994 562898 374026 563134
rect 374262 562898 374346 563134
rect 374582 562898 374614 563134
rect 373994 536454 374614 562898
rect 373994 536218 374026 536454
rect 374262 536218 374346 536454
rect 374582 536218 374614 536454
rect 373994 536134 374614 536218
rect 373994 535898 374026 536134
rect 374262 535898 374346 536134
rect 374582 535898 374614 536134
rect 373994 509454 374614 535898
rect 373994 509218 374026 509454
rect 374262 509218 374346 509454
rect 374582 509218 374614 509454
rect 373994 509134 374614 509218
rect 373994 508898 374026 509134
rect 374262 508898 374346 509134
rect 374582 508898 374614 509134
rect 373994 482454 374614 508898
rect 373994 482218 374026 482454
rect 374262 482218 374346 482454
rect 374582 482218 374614 482454
rect 373994 482134 374614 482218
rect 373994 481898 374026 482134
rect 374262 481898 374346 482134
rect 374582 481898 374614 482134
rect 373994 455454 374614 481898
rect 373994 455218 374026 455454
rect 374262 455218 374346 455454
rect 374582 455218 374614 455454
rect 373994 455134 374614 455218
rect 373994 454898 374026 455134
rect 374262 454898 374346 455134
rect 374582 454898 374614 455134
rect 373994 428454 374614 454898
rect 373994 428218 374026 428454
rect 374262 428218 374346 428454
rect 374582 428218 374614 428454
rect 373994 428134 374614 428218
rect 373994 427898 374026 428134
rect 374262 427898 374346 428134
rect 374582 427898 374614 428134
rect 373994 401454 374614 427898
rect 373994 401218 374026 401454
rect 374262 401218 374346 401454
rect 374582 401218 374614 401454
rect 373994 401134 374614 401218
rect 373994 400898 374026 401134
rect 374262 400898 374346 401134
rect 374582 400898 374614 401134
rect 373994 374454 374614 400898
rect 373994 374218 374026 374454
rect 374262 374218 374346 374454
rect 374582 374218 374614 374454
rect 373994 374134 374614 374218
rect 373994 373898 374026 374134
rect 374262 373898 374346 374134
rect 374582 373898 374614 374134
rect 373994 347454 374614 373898
rect 373994 347218 374026 347454
rect 374262 347218 374346 347454
rect 374582 347218 374614 347454
rect 373994 347134 374614 347218
rect 373994 346898 374026 347134
rect 374262 346898 374346 347134
rect 374582 346898 374614 347134
rect 373994 320454 374614 346898
rect 373994 320218 374026 320454
rect 374262 320218 374346 320454
rect 374582 320218 374614 320454
rect 373994 320134 374614 320218
rect 373994 319898 374026 320134
rect 374262 319898 374346 320134
rect 374582 319898 374614 320134
rect 373994 293454 374614 319898
rect 373994 293218 374026 293454
rect 374262 293218 374346 293454
rect 374582 293218 374614 293454
rect 373994 293134 374614 293218
rect 373994 292898 374026 293134
rect 374262 292898 374346 293134
rect 374582 292898 374614 293134
rect 373994 266454 374614 292898
rect 373994 266218 374026 266454
rect 374262 266218 374346 266454
rect 374582 266218 374614 266454
rect 373994 266134 374614 266218
rect 373994 265898 374026 266134
rect 374262 265898 374346 266134
rect 374582 265898 374614 266134
rect 373994 239454 374614 265898
rect 373994 239218 374026 239454
rect 374262 239218 374346 239454
rect 374582 239218 374614 239454
rect 373994 239134 374614 239218
rect 373994 238898 374026 239134
rect 374262 238898 374346 239134
rect 374582 238898 374614 239134
rect 373994 212454 374614 238898
rect 373994 212218 374026 212454
rect 374262 212218 374346 212454
rect 374582 212218 374614 212454
rect 373994 212134 374614 212218
rect 373994 211898 374026 212134
rect 374262 211898 374346 212134
rect 374582 211898 374614 212134
rect 373994 185454 374614 211898
rect 373994 185218 374026 185454
rect 374262 185218 374346 185454
rect 374582 185218 374614 185454
rect 373994 185134 374614 185218
rect 373994 184898 374026 185134
rect 374262 184898 374346 185134
rect 374582 184898 374614 185134
rect 373994 158454 374614 184898
rect 373994 158218 374026 158454
rect 374262 158218 374346 158454
rect 374582 158218 374614 158454
rect 373994 158134 374614 158218
rect 373994 157898 374026 158134
rect 374262 157898 374346 158134
rect 374582 157898 374614 158134
rect 373994 131454 374614 157898
rect 373994 131218 374026 131454
rect 374262 131218 374346 131454
rect 374582 131218 374614 131454
rect 373994 131134 374614 131218
rect 373994 130898 374026 131134
rect 374262 130898 374346 131134
rect 374582 130898 374614 131134
rect 373994 104454 374614 130898
rect 373994 104218 374026 104454
rect 374262 104218 374346 104454
rect 374582 104218 374614 104454
rect 373994 104134 374614 104218
rect 373994 103898 374026 104134
rect 374262 103898 374346 104134
rect 374582 103898 374614 104134
rect 373994 77454 374614 103898
rect 373994 77218 374026 77454
rect 374262 77218 374346 77454
rect 374582 77218 374614 77454
rect 373994 77134 374614 77218
rect 373994 76898 374026 77134
rect 374262 76898 374346 77134
rect 374582 76898 374614 77134
rect 373994 69000 374614 76898
rect 377494 704838 378114 711590
rect 377494 704602 377526 704838
rect 377762 704602 377846 704838
rect 378082 704602 378114 704838
rect 377494 704518 378114 704602
rect 377494 704282 377526 704518
rect 377762 704282 377846 704518
rect 378082 704282 378114 704518
rect 377494 701829 378114 704282
rect 377494 701593 377526 701829
rect 377762 701593 377846 701829
rect 378082 701593 378114 701829
rect 377494 701509 378114 701593
rect 377494 701273 377526 701509
rect 377762 701273 377846 701509
rect 378082 701273 378114 701509
rect 377494 674829 378114 701273
rect 401994 705798 402614 711590
rect 401994 705562 402026 705798
rect 402262 705562 402346 705798
rect 402582 705562 402614 705798
rect 401994 705478 402614 705562
rect 401994 705242 402026 705478
rect 402262 705242 402346 705478
rect 402582 705242 402614 705478
rect 397683 699820 397749 699821
rect 397683 699756 397684 699820
rect 397748 699756 397749 699820
rect 397683 699755 397749 699756
rect 377494 674593 377526 674829
rect 377762 674593 377846 674829
rect 378082 674593 378114 674829
rect 377494 674509 378114 674593
rect 377494 674273 377526 674509
rect 377762 674273 377846 674509
rect 378082 674273 378114 674509
rect 377494 647829 378114 674273
rect 377494 647593 377526 647829
rect 377762 647593 377846 647829
rect 378082 647593 378114 647829
rect 377494 647509 378114 647593
rect 377494 647273 377526 647509
rect 377762 647273 377846 647509
rect 378082 647273 378114 647509
rect 377494 620829 378114 647273
rect 377494 620593 377526 620829
rect 377762 620593 377846 620829
rect 378082 620593 378114 620829
rect 377494 620509 378114 620593
rect 377494 620273 377526 620509
rect 377762 620273 377846 620509
rect 378082 620273 378114 620509
rect 377494 593829 378114 620273
rect 377494 593593 377526 593829
rect 377762 593593 377846 593829
rect 378082 593593 378114 593829
rect 377494 593509 378114 593593
rect 377494 593273 377526 593509
rect 377762 593273 377846 593509
rect 378082 593273 378114 593509
rect 377494 566829 378114 593273
rect 377494 566593 377526 566829
rect 377762 566593 377846 566829
rect 378082 566593 378114 566829
rect 377494 566509 378114 566593
rect 377494 566273 377526 566509
rect 377762 566273 377846 566509
rect 378082 566273 378114 566509
rect 377494 539829 378114 566273
rect 377494 539593 377526 539829
rect 377762 539593 377846 539829
rect 378082 539593 378114 539829
rect 377494 539509 378114 539593
rect 377494 539273 377526 539509
rect 377762 539273 377846 539509
rect 378082 539273 378114 539509
rect 377494 512829 378114 539273
rect 377494 512593 377526 512829
rect 377762 512593 377846 512829
rect 378082 512593 378114 512829
rect 377494 512509 378114 512593
rect 377494 512273 377526 512509
rect 377762 512273 377846 512509
rect 378082 512273 378114 512509
rect 377494 485829 378114 512273
rect 377494 485593 377526 485829
rect 377762 485593 377846 485829
rect 378082 485593 378114 485829
rect 377494 485509 378114 485593
rect 377494 485273 377526 485509
rect 377762 485273 377846 485509
rect 378082 485273 378114 485509
rect 377494 458829 378114 485273
rect 377494 458593 377526 458829
rect 377762 458593 377846 458829
rect 378082 458593 378114 458829
rect 377494 458509 378114 458593
rect 377494 458273 377526 458509
rect 377762 458273 377846 458509
rect 378082 458273 378114 458509
rect 377494 431829 378114 458273
rect 377494 431593 377526 431829
rect 377762 431593 377846 431829
rect 378082 431593 378114 431829
rect 377494 431509 378114 431593
rect 377494 431273 377526 431509
rect 377762 431273 377846 431509
rect 378082 431273 378114 431509
rect 377494 404829 378114 431273
rect 377494 404593 377526 404829
rect 377762 404593 377846 404829
rect 378082 404593 378114 404829
rect 377494 404509 378114 404593
rect 377494 404273 377526 404509
rect 377762 404273 377846 404509
rect 378082 404273 378114 404509
rect 377494 377829 378114 404273
rect 377494 377593 377526 377829
rect 377762 377593 377846 377829
rect 378082 377593 378114 377829
rect 377494 377509 378114 377593
rect 377494 377273 377526 377509
rect 377762 377273 377846 377509
rect 378082 377273 378114 377509
rect 377494 350829 378114 377273
rect 377494 350593 377526 350829
rect 377762 350593 377846 350829
rect 378082 350593 378114 350829
rect 377494 350509 378114 350593
rect 377494 350273 377526 350509
rect 377762 350273 377846 350509
rect 378082 350273 378114 350509
rect 377494 323829 378114 350273
rect 377494 323593 377526 323829
rect 377762 323593 377846 323829
rect 378082 323593 378114 323829
rect 377494 323509 378114 323593
rect 377494 323273 377526 323509
rect 377762 323273 377846 323509
rect 378082 323273 378114 323509
rect 377494 296829 378114 323273
rect 377494 296593 377526 296829
rect 377762 296593 377846 296829
rect 378082 296593 378114 296829
rect 377494 296509 378114 296593
rect 377494 296273 377526 296509
rect 377762 296273 377846 296509
rect 378082 296273 378114 296509
rect 377494 269829 378114 296273
rect 377494 269593 377526 269829
rect 377762 269593 377846 269829
rect 378082 269593 378114 269829
rect 377494 269509 378114 269593
rect 377494 269273 377526 269509
rect 377762 269273 377846 269509
rect 378082 269273 378114 269509
rect 377494 242829 378114 269273
rect 377494 242593 377526 242829
rect 377762 242593 377846 242829
rect 378082 242593 378114 242829
rect 377494 242509 378114 242593
rect 377494 242273 377526 242509
rect 377762 242273 377846 242509
rect 378082 242273 378114 242509
rect 377494 215829 378114 242273
rect 377494 215593 377526 215829
rect 377762 215593 377846 215829
rect 378082 215593 378114 215829
rect 377494 215509 378114 215593
rect 377494 215273 377526 215509
rect 377762 215273 377846 215509
rect 378082 215273 378114 215509
rect 377494 188829 378114 215273
rect 377494 188593 377526 188829
rect 377762 188593 377846 188829
rect 378082 188593 378114 188829
rect 377494 188509 378114 188593
rect 377494 188273 377526 188509
rect 377762 188273 377846 188509
rect 378082 188273 378114 188509
rect 377494 161829 378114 188273
rect 377494 161593 377526 161829
rect 377762 161593 377846 161829
rect 378082 161593 378114 161829
rect 377494 161509 378114 161593
rect 377494 161273 377526 161509
rect 377762 161273 377846 161509
rect 378082 161273 378114 161509
rect 377494 134829 378114 161273
rect 377494 134593 377526 134829
rect 377762 134593 377846 134829
rect 378082 134593 378114 134829
rect 377494 134509 378114 134593
rect 377494 134273 377526 134509
rect 377762 134273 377846 134509
rect 378082 134273 378114 134509
rect 377494 107829 378114 134273
rect 377494 107593 377526 107829
rect 377762 107593 377846 107829
rect 378082 107593 378114 107829
rect 377494 107509 378114 107593
rect 377494 107273 377526 107509
rect 377762 107273 377846 107509
rect 378082 107273 378114 107509
rect 377494 80829 378114 107273
rect 377494 80593 377526 80829
rect 377762 80593 377846 80829
rect 378082 80593 378114 80829
rect 377494 80509 378114 80593
rect 377494 80273 377526 80509
rect 377762 80273 377846 80509
rect 378082 80273 378114 80509
rect 377494 69000 378114 80273
rect 249011 65652 249077 65653
rect 249011 65588 249012 65652
rect 249076 65588 249077 65652
rect 249011 65587 249077 65588
rect 277899 65652 277965 65653
rect 277899 65588 277900 65652
rect 277964 65588 277965 65652
rect 277899 65587 277965 65588
rect 306971 65652 307037 65653
rect 306971 65588 306972 65652
rect 307036 65588 307037 65652
rect 306971 65587 307037 65588
rect 335859 65652 335925 65653
rect 335859 65588 335860 65652
rect 335924 65588 335925 65652
rect 335859 65587 335925 65588
rect 364931 65652 364997 65653
rect 364931 65588 364932 65652
rect 364996 65588 364997 65652
rect 364931 65587 364997 65588
rect 393819 65652 393885 65653
rect 393819 65588 393820 65652
rect 393884 65588 393885 65652
rect 393819 65587 393885 65588
rect 181494 53593 181526 53829
rect 181762 53593 181846 53829
rect 182082 53593 182114 53829
rect 181494 53509 182114 53593
rect 181494 53273 181526 53509
rect 181762 53273 181846 53509
rect 182082 53273 182114 53509
rect 181494 42000 182114 53273
rect 192918 53829 193238 53861
rect 192918 53593 192960 53829
rect 193196 53593 193238 53829
rect 192918 53509 193238 53593
rect 192918 53273 192960 53509
rect 193196 53273 193238 53509
rect 192918 53241 193238 53273
rect 196866 53829 197186 53861
rect 196866 53593 196908 53829
rect 197144 53593 197186 53829
rect 196866 53509 197186 53593
rect 196866 53273 196908 53509
rect 197144 53273 197186 53509
rect 196866 53241 197186 53273
rect 200814 53829 201134 53861
rect 200814 53593 200856 53829
rect 201092 53593 201134 53829
rect 200814 53509 201134 53593
rect 200814 53273 200856 53509
rect 201092 53273 201134 53509
rect 200814 53241 201134 53273
rect 204762 53829 205082 53861
rect 204762 53593 204804 53829
rect 205040 53593 205082 53829
rect 204762 53509 205082 53593
rect 204762 53273 204804 53509
rect 205040 53273 205082 53509
rect 204762 53241 205082 53273
rect 213218 53829 213538 53861
rect 213218 53593 213260 53829
rect 213496 53593 213538 53829
rect 213218 53509 213538 53593
rect 213218 53273 213260 53509
rect 213496 53273 213538 53509
rect 213218 53241 213538 53273
rect 214166 53829 214486 53861
rect 214166 53593 214208 53829
rect 214444 53593 214486 53829
rect 214166 53509 214486 53593
rect 214166 53273 214208 53509
rect 214444 53273 214486 53509
rect 214166 53241 214486 53273
rect 215114 53829 215434 53861
rect 215114 53593 215156 53829
rect 215392 53593 215434 53829
rect 215114 53509 215434 53593
rect 215114 53273 215156 53509
rect 215392 53273 215434 53509
rect 215114 53241 215434 53273
rect 216062 53829 216382 53861
rect 216062 53593 216104 53829
rect 216340 53593 216382 53829
rect 216062 53509 216382 53593
rect 216062 53273 216104 53509
rect 216340 53273 216382 53509
rect 216062 53241 216382 53273
rect 221918 53829 222238 53861
rect 221918 53593 221960 53829
rect 222196 53593 222238 53829
rect 221918 53509 222238 53593
rect 221918 53273 221960 53509
rect 222196 53273 222238 53509
rect 221918 53241 222238 53273
rect 225866 53829 226186 53861
rect 225866 53593 225908 53829
rect 226144 53593 226186 53829
rect 225866 53509 226186 53593
rect 225866 53273 225908 53509
rect 226144 53273 226186 53509
rect 225866 53241 226186 53273
rect 229814 53829 230134 53861
rect 229814 53593 229856 53829
rect 230092 53593 230134 53829
rect 229814 53509 230134 53593
rect 229814 53273 229856 53509
rect 230092 53273 230134 53509
rect 229814 53241 230134 53273
rect 233762 53829 234082 53861
rect 233762 53593 233804 53829
rect 234040 53593 234082 53829
rect 233762 53509 234082 53593
rect 233762 53273 233804 53509
rect 234040 53273 234082 53509
rect 233762 53241 234082 53273
rect 242218 53829 242538 53861
rect 242218 53593 242260 53829
rect 242496 53593 242538 53829
rect 242218 53509 242538 53593
rect 242218 53273 242260 53509
rect 242496 53273 242538 53509
rect 242218 53241 242538 53273
rect 243166 53829 243486 53861
rect 243166 53593 243208 53829
rect 243444 53593 243486 53829
rect 243166 53509 243486 53593
rect 243166 53273 243208 53509
rect 243444 53273 243486 53509
rect 243166 53241 243486 53273
rect 244114 53829 244434 53861
rect 244114 53593 244156 53829
rect 244392 53593 244434 53829
rect 244114 53509 244434 53593
rect 244114 53273 244156 53509
rect 244392 53273 244434 53509
rect 244114 53241 244434 53273
rect 245062 53829 245382 53861
rect 245062 53593 245104 53829
rect 245340 53593 245382 53829
rect 245062 53509 245382 53593
rect 245062 53273 245104 53509
rect 245340 53273 245382 53509
rect 245062 53241 245382 53273
rect 194892 50454 195212 50486
rect 194892 50218 194934 50454
rect 195170 50218 195212 50454
rect 194892 50134 195212 50218
rect 194892 49898 194934 50134
rect 195170 49898 195212 50134
rect 194892 49866 195212 49898
rect 198840 50454 199160 50486
rect 198840 50218 198882 50454
rect 199118 50218 199160 50454
rect 198840 50134 199160 50218
rect 198840 49898 198882 50134
rect 199118 49898 199160 50134
rect 198840 49866 199160 49898
rect 202788 50454 203108 50486
rect 202788 50218 202830 50454
rect 203066 50218 203108 50454
rect 202788 50134 203108 50218
rect 202788 49898 202830 50134
rect 203066 49898 203108 50134
rect 202788 49866 203108 49898
rect 213692 50454 214012 50486
rect 213692 50218 213734 50454
rect 213970 50218 214012 50454
rect 213692 50134 214012 50218
rect 213692 49898 213734 50134
rect 213970 49898 214012 50134
rect 213692 49866 214012 49898
rect 214640 50454 214960 50486
rect 214640 50218 214682 50454
rect 214918 50218 214960 50454
rect 214640 50134 214960 50218
rect 214640 49898 214682 50134
rect 214918 49898 214960 50134
rect 214640 49866 214960 49898
rect 215588 50454 215908 50486
rect 215588 50218 215630 50454
rect 215866 50218 215908 50454
rect 215588 50134 215908 50218
rect 215588 49898 215630 50134
rect 215866 49898 215908 50134
rect 215588 49866 215908 49898
rect 223892 50454 224212 50486
rect 223892 50218 223934 50454
rect 224170 50218 224212 50454
rect 223892 50134 224212 50218
rect 223892 49898 223934 50134
rect 224170 49898 224212 50134
rect 223892 49866 224212 49898
rect 227840 50454 228160 50486
rect 227840 50218 227882 50454
rect 228118 50218 228160 50454
rect 227840 50134 228160 50218
rect 227840 49898 227882 50134
rect 228118 49898 228160 50134
rect 227840 49866 228160 49898
rect 231788 50454 232108 50486
rect 231788 50218 231830 50454
rect 232066 50218 232108 50454
rect 231788 50134 232108 50218
rect 231788 49898 231830 50134
rect 232066 49898 232108 50134
rect 231788 49866 232108 49898
rect 242692 50454 243012 50486
rect 242692 50218 242734 50454
rect 242970 50218 243012 50454
rect 242692 50134 243012 50218
rect 242692 49898 242734 50134
rect 242970 49898 243012 50134
rect 242692 49866 243012 49898
rect 243640 50454 243960 50486
rect 243640 50218 243682 50454
rect 243918 50218 243960 50454
rect 243640 50134 243960 50218
rect 243640 49898 243682 50134
rect 243918 49898 243960 50134
rect 243640 49866 243960 49898
rect 244588 50454 244908 50486
rect 244588 50218 244630 50454
rect 244866 50218 244908 50454
rect 244588 50134 244908 50218
rect 244588 49898 244630 50134
rect 244866 49898 244908 50134
rect 244588 49866 244908 49898
rect 249014 43349 249074 65587
rect 250918 53829 251238 53861
rect 250918 53593 250960 53829
rect 251196 53593 251238 53829
rect 250918 53509 251238 53593
rect 250918 53273 250960 53509
rect 251196 53273 251238 53509
rect 250918 53241 251238 53273
rect 254866 53829 255186 53861
rect 254866 53593 254908 53829
rect 255144 53593 255186 53829
rect 254866 53509 255186 53593
rect 254866 53273 254908 53509
rect 255144 53273 255186 53509
rect 254866 53241 255186 53273
rect 258814 53829 259134 53861
rect 258814 53593 258856 53829
rect 259092 53593 259134 53829
rect 258814 53509 259134 53593
rect 258814 53273 258856 53509
rect 259092 53273 259134 53509
rect 258814 53241 259134 53273
rect 262762 53829 263082 53861
rect 262762 53593 262804 53829
rect 263040 53593 263082 53829
rect 262762 53509 263082 53593
rect 262762 53273 262804 53509
rect 263040 53273 263082 53509
rect 262762 53241 263082 53273
rect 271218 53829 271538 53861
rect 271218 53593 271260 53829
rect 271496 53593 271538 53829
rect 271218 53509 271538 53593
rect 271218 53273 271260 53509
rect 271496 53273 271538 53509
rect 271218 53241 271538 53273
rect 272166 53829 272486 53861
rect 272166 53593 272208 53829
rect 272444 53593 272486 53829
rect 272166 53509 272486 53593
rect 272166 53273 272208 53509
rect 272444 53273 272486 53509
rect 272166 53241 272486 53273
rect 273114 53829 273434 53861
rect 273114 53593 273156 53829
rect 273392 53593 273434 53829
rect 273114 53509 273434 53593
rect 273114 53273 273156 53509
rect 273392 53273 273434 53509
rect 273114 53241 273434 53273
rect 274062 53829 274382 53861
rect 274062 53593 274104 53829
rect 274340 53593 274382 53829
rect 274062 53509 274382 53593
rect 274062 53273 274104 53509
rect 274340 53273 274382 53509
rect 274062 53241 274382 53273
rect 252892 50454 253212 50486
rect 252892 50218 252934 50454
rect 253170 50218 253212 50454
rect 252892 50134 253212 50218
rect 252892 49898 252934 50134
rect 253170 49898 253212 50134
rect 252892 49866 253212 49898
rect 256840 50454 257160 50486
rect 256840 50218 256882 50454
rect 257118 50218 257160 50454
rect 256840 50134 257160 50218
rect 256840 49898 256882 50134
rect 257118 49898 257160 50134
rect 256840 49866 257160 49898
rect 260788 50454 261108 50486
rect 260788 50218 260830 50454
rect 261066 50218 261108 50454
rect 260788 50134 261108 50218
rect 260788 49898 260830 50134
rect 261066 49898 261108 50134
rect 260788 49866 261108 49898
rect 271692 50454 272012 50486
rect 271692 50218 271734 50454
rect 271970 50218 272012 50454
rect 271692 50134 272012 50218
rect 271692 49898 271734 50134
rect 271970 49898 272012 50134
rect 271692 49866 272012 49898
rect 272640 50454 272960 50486
rect 272640 50218 272682 50454
rect 272918 50218 272960 50454
rect 272640 50134 272960 50218
rect 272640 49898 272682 50134
rect 272918 49898 272960 50134
rect 272640 49866 272960 49898
rect 273588 50454 273908 50486
rect 273588 50218 273630 50454
rect 273866 50218 273908 50454
rect 273588 50134 273908 50218
rect 273588 49898 273630 50134
rect 273866 49898 273908 50134
rect 273588 49866 273908 49898
rect 277902 43621 277962 65587
rect 279918 53829 280238 53861
rect 279918 53593 279960 53829
rect 280196 53593 280238 53829
rect 279918 53509 280238 53593
rect 279918 53273 279960 53509
rect 280196 53273 280238 53509
rect 279918 53241 280238 53273
rect 283866 53829 284186 53861
rect 283866 53593 283908 53829
rect 284144 53593 284186 53829
rect 283866 53509 284186 53593
rect 283866 53273 283908 53509
rect 284144 53273 284186 53509
rect 283866 53241 284186 53273
rect 287814 53829 288134 53861
rect 287814 53593 287856 53829
rect 288092 53593 288134 53829
rect 287814 53509 288134 53593
rect 287814 53273 287856 53509
rect 288092 53273 288134 53509
rect 287814 53241 288134 53273
rect 291762 53829 292082 53861
rect 291762 53593 291804 53829
rect 292040 53593 292082 53829
rect 291762 53509 292082 53593
rect 291762 53273 291804 53509
rect 292040 53273 292082 53509
rect 291762 53241 292082 53273
rect 300218 53829 300538 53861
rect 300218 53593 300260 53829
rect 300496 53593 300538 53829
rect 300218 53509 300538 53593
rect 300218 53273 300260 53509
rect 300496 53273 300538 53509
rect 300218 53241 300538 53273
rect 301166 53829 301486 53861
rect 301166 53593 301208 53829
rect 301444 53593 301486 53829
rect 301166 53509 301486 53593
rect 301166 53273 301208 53509
rect 301444 53273 301486 53509
rect 301166 53241 301486 53273
rect 302114 53829 302434 53861
rect 302114 53593 302156 53829
rect 302392 53593 302434 53829
rect 302114 53509 302434 53593
rect 302114 53273 302156 53509
rect 302392 53273 302434 53509
rect 302114 53241 302434 53273
rect 303062 53829 303382 53861
rect 303062 53593 303104 53829
rect 303340 53593 303382 53829
rect 303062 53509 303382 53593
rect 303062 53273 303104 53509
rect 303340 53273 303382 53509
rect 303062 53241 303382 53273
rect 281892 50454 282212 50486
rect 281892 50218 281934 50454
rect 282170 50218 282212 50454
rect 281892 50134 282212 50218
rect 281892 49898 281934 50134
rect 282170 49898 282212 50134
rect 281892 49866 282212 49898
rect 285840 50454 286160 50486
rect 285840 50218 285882 50454
rect 286118 50218 286160 50454
rect 285840 50134 286160 50218
rect 285840 49898 285882 50134
rect 286118 49898 286160 50134
rect 285840 49866 286160 49898
rect 289788 50454 290108 50486
rect 289788 50218 289830 50454
rect 290066 50218 290108 50454
rect 289788 50134 290108 50218
rect 289788 49898 289830 50134
rect 290066 49898 290108 50134
rect 289788 49866 290108 49898
rect 300692 50454 301012 50486
rect 300692 50218 300734 50454
rect 300970 50218 301012 50454
rect 300692 50134 301012 50218
rect 300692 49898 300734 50134
rect 300970 49898 301012 50134
rect 300692 49866 301012 49898
rect 301640 50454 301960 50486
rect 301640 50218 301682 50454
rect 301918 50218 301960 50454
rect 301640 50134 301960 50218
rect 301640 49898 301682 50134
rect 301918 49898 301960 50134
rect 301640 49866 301960 49898
rect 302588 50454 302908 50486
rect 302588 50218 302630 50454
rect 302866 50218 302908 50454
rect 302588 50134 302908 50218
rect 302588 49898 302630 50134
rect 302866 49898 302908 50134
rect 302588 49866 302908 49898
rect 306974 43621 307034 65587
rect 308918 53829 309238 53861
rect 308918 53593 308960 53829
rect 309196 53593 309238 53829
rect 308918 53509 309238 53593
rect 308918 53273 308960 53509
rect 309196 53273 309238 53509
rect 308918 53241 309238 53273
rect 312866 53829 313186 53861
rect 312866 53593 312908 53829
rect 313144 53593 313186 53829
rect 312866 53509 313186 53593
rect 312866 53273 312908 53509
rect 313144 53273 313186 53509
rect 312866 53241 313186 53273
rect 316814 53829 317134 53861
rect 316814 53593 316856 53829
rect 317092 53593 317134 53829
rect 316814 53509 317134 53593
rect 316814 53273 316856 53509
rect 317092 53273 317134 53509
rect 316814 53241 317134 53273
rect 320762 53829 321082 53861
rect 320762 53593 320804 53829
rect 321040 53593 321082 53829
rect 320762 53509 321082 53593
rect 320762 53273 320804 53509
rect 321040 53273 321082 53509
rect 320762 53241 321082 53273
rect 329218 53829 329538 53861
rect 329218 53593 329260 53829
rect 329496 53593 329538 53829
rect 329218 53509 329538 53593
rect 329218 53273 329260 53509
rect 329496 53273 329538 53509
rect 329218 53241 329538 53273
rect 330166 53829 330486 53861
rect 330166 53593 330208 53829
rect 330444 53593 330486 53829
rect 330166 53509 330486 53593
rect 330166 53273 330208 53509
rect 330444 53273 330486 53509
rect 330166 53241 330486 53273
rect 331114 53829 331434 53861
rect 331114 53593 331156 53829
rect 331392 53593 331434 53829
rect 331114 53509 331434 53593
rect 331114 53273 331156 53509
rect 331392 53273 331434 53509
rect 331114 53241 331434 53273
rect 332062 53829 332382 53861
rect 332062 53593 332104 53829
rect 332340 53593 332382 53829
rect 332062 53509 332382 53593
rect 332062 53273 332104 53509
rect 332340 53273 332382 53509
rect 332062 53241 332382 53273
rect 310892 50454 311212 50486
rect 310892 50218 310934 50454
rect 311170 50218 311212 50454
rect 310892 50134 311212 50218
rect 310892 49898 310934 50134
rect 311170 49898 311212 50134
rect 310892 49866 311212 49898
rect 314840 50454 315160 50486
rect 314840 50218 314882 50454
rect 315118 50218 315160 50454
rect 314840 50134 315160 50218
rect 314840 49898 314882 50134
rect 315118 49898 315160 50134
rect 314840 49866 315160 49898
rect 318788 50454 319108 50486
rect 318788 50218 318830 50454
rect 319066 50218 319108 50454
rect 318788 50134 319108 50218
rect 318788 49898 318830 50134
rect 319066 49898 319108 50134
rect 318788 49866 319108 49898
rect 329692 50454 330012 50486
rect 329692 50218 329734 50454
rect 329970 50218 330012 50454
rect 329692 50134 330012 50218
rect 329692 49898 329734 50134
rect 329970 49898 330012 50134
rect 329692 49866 330012 49898
rect 330640 50454 330960 50486
rect 330640 50218 330682 50454
rect 330918 50218 330960 50454
rect 330640 50134 330960 50218
rect 330640 49898 330682 50134
rect 330918 49898 330960 50134
rect 330640 49866 330960 49898
rect 331588 50454 331908 50486
rect 331588 50218 331630 50454
rect 331866 50218 331908 50454
rect 331588 50134 331908 50218
rect 331588 49898 331630 50134
rect 331866 49898 331908 50134
rect 331588 49866 331908 49898
rect 335862 43621 335922 65587
rect 337918 53829 338238 53861
rect 337918 53593 337960 53829
rect 338196 53593 338238 53829
rect 337918 53509 338238 53593
rect 337918 53273 337960 53509
rect 338196 53273 338238 53509
rect 337918 53241 338238 53273
rect 341866 53829 342186 53861
rect 341866 53593 341908 53829
rect 342144 53593 342186 53829
rect 341866 53509 342186 53593
rect 341866 53273 341908 53509
rect 342144 53273 342186 53509
rect 341866 53241 342186 53273
rect 345814 53829 346134 53861
rect 345814 53593 345856 53829
rect 346092 53593 346134 53829
rect 345814 53509 346134 53593
rect 345814 53273 345856 53509
rect 346092 53273 346134 53509
rect 345814 53241 346134 53273
rect 349762 53829 350082 53861
rect 349762 53593 349804 53829
rect 350040 53593 350082 53829
rect 349762 53509 350082 53593
rect 349762 53273 349804 53509
rect 350040 53273 350082 53509
rect 349762 53241 350082 53273
rect 358218 53829 358538 53861
rect 358218 53593 358260 53829
rect 358496 53593 358538 53829
rect 358218 53509 358538 53593
rect 358218 53273 358260 53509
rect 358496 53273 358538 53509
rect 358218 53241 358538 53273
rect 359166 53829 359486 53861
rect 359166 53593 359208 53829
rect 359444 53593 359486 53829
rect 359166 53509 359486 53593
rect 359166 53273 359208 53509
rect 359444 53273 359486 53509
rect 359166 53241 359486 53273
rect 360114 53829 360434 53861
rect 360114 53593 360156 53829
rect 360392 53593 360434 53829
rect 360114 53509 360434 53593
rect 360114 53273 360156 53509
rect 360392 53273 360434 53509
rect 360114 53241 360434 53273
rect 361062 53829 361382 53861
rect 361062 53593 361104 53829
rect 361340 53593 361382 53829
rect 361062 53509 361382 53593
rect 361062 53273 361104 53509
rect 361340 53273 361382 53509
rect 361062 53241 361382 53273
rect 339892 50454 340212 50486
rect 339892 50218 339934 50454
rect 340170 50218 340212 50454
rect 339892 50134 340212 50218
rect 339892 49898 339934 50134
rect 340170 49898 340212 50134
rect 339892 49866 340212 49898
rect 343840 50454 344160 50486
rect 343840 50218 343882 50454
rect 344118 50218 344160 50454
rect 343840 50134 344160 50218
rect 343840 49898 343882 50134
rect 344118 49898 344160 50134
rect 343840 49866 344160 49898
rect 347788 50454 348108 50486
rect 347788 50218 347830 50454
rect 348066 50218 348108 50454
rect 347788 50134 348108 50218
rect 347788 49898 347830 50134
rect 348066 49898 348108 50134
rect 347788 49866 348108 49898
rect 358692 50454 359012 50486
rect 358692 50218 358734 50454
rect 358970 50218 359012 50454
rect 358692 50134 359012 50218
rect 358692 49898 358734 50134
rect 358970 49898 359012 50134
rect 358692 49866 359012 49898
rect 359640 50454 359960 50486
rect 359640 50218 359682 50454
rect 359918 50218 359960 50454
rect 359640 50134 359960 50218
rect 359640 49898 359682 50134
rect 359918 49898 359960 50134
rect 359640 49866 359960 49898
rect 360588 50454 360908 50486
rect 360588 50218 360630 50454
rect 360866 50218 360908 50454
rect 360588 50134 360908 50218
rect 360588 49898 360630 50134
rect 360866 49898 360908 50134
rect 360588 49866 360908 49898
rect 364934 43621 364994 65587
rect 366918 53829 367238 53861
rect 366918 53593 366960 53829
rect 367196 53593 367238 53829
rect 366918 53509 367238 53593
rect 366918 53273 366960 53509
rect 367196 53273 367238 53509
rect 366918 53241 367238 53273
rect 370866 53829 371186 53861
rect 370866 53593 370908 53829
rect 371144 53593 371186 53829
rect 370866 53509 371186 53593
rect 370866 53273 370908 53509
rect 371144 53273 371186 53509
rect 370866 53241 371186 53273
rect 374814 53829 375134 53861
rect 374814 53593 374856 53829
rect 375092 53593 375134 53829
rect 374814 53509 375134 53593
rect 374814 53273 374856 53509
rect 375092 53273 375134 53509
rect 374814 53241 375134 53273
rect 378762 53829 379082 53861
rect 378762 53593 378804 53829
rect 379040 53593 379082 53829
rect 378762 53509 379082 53593
rect 378762 53273 378804 53509
rect 379040 53273 379082 53509
rect 378762 53241 379082 53273
rect 387218 53829 387538 53861
rect 387218 53593 387260 53829
rect 387496 53593 387538 53829
rect 387218 53509 387538 53593
rect 387218 53273 387260 53509
rect 387496 53273 387538 53509
rect 387218 53241 387538 53273
rect 388166 53829 388486 53861
rect 388166 53593 388208 53829
rect 388444 53593 388486 53829
rect 388166 53509 388486 53593
rect 388166 53273 388208 53509
rect 388444 53273 388486 53509
rect 388166 53241 388486 53273
rect 389114 53829 389434 53861
rect 389114 53593 389156 53829
rect 389392 53593 389434 53829
rect 389114 53509 389434 53593
rect 389114 53273 389156 53509
rect 389392 53273 389434 53509
rect 389114 53241 389434 53273
rect 390062 53829 390382 53861
rect 390062 53593 390104 53829
rect 390340 53593 390382 53829
rect 390062 53509 390382 53593
rect 390062 53273 390104 53509
rect 390340 53273 390382 53509
rect 390062 53241 390382 53273
rect 368892 50454 369212 50486
rect 368892 50218 368934 50454
rect 369170 50218 369212 50454
rect 368892 50134 369212 50218
rect 368892 49898 368934 50134
rect 369170 49898 369212 50134
rect 368892 49866 369212 49898
rect 372840 50454 373160 50486
rect 372840 50218 372882 50454
rect 373118 50218 373160 50454
rect 372840 50134 373160 50218
rect 372840 49898 372882 50134
rect 373118 49898 373160 50134
rect 372840 49866 373160 49898
rect 376788 50454 377108 50486
rect 376788 50218 376830 50454
rect 377066 50218 377108 50454
rect 376788 50134 377108 50218
rect 376788 49898 376830 50134
rect 377066 49898 377108 50134
rect 376788 49866 377108 49898
rect 387692 50454 388012 50486
rect 387692 50218 387734 50454
rect 387970 50218 388012 50454
rect 387692 50134 388012 50218
rect 387692 49898 387734 50134
rect 387970 49898 388012 50134
rect 387692 49866 388012 49898
rect 388640 50454 388960 50486
rect 388640 50218 388682 50454
rect 388918 50218 388960 50454
rect 388640 50134 388960 50218
rect 388640 49898 388682 50134
rect 388918 49898 388960 50134
rect 388640 49866 388960 49898
rect 389588 50454 389908 50486
rect 389588 50218 389630 50454
rect 389866 50218 389908 50454
rect 389588 50134 389908 50218
rect 389588 49898 389630 50134
rect 389866 49898 389908 50134
rect 389588 49866 389908 49898
rect 393822 43621 393882 65587
rect 395918 53829 396238 53861
rect 395918 53593 395960 53829
rect 396196 53593 396238 53829
rect 395918 53509 396238 53593
rect 395918 53273 395960 53509
rect 396196 53273 396238 53509
rect 395918 53241 396238 53273
rect 277899 43620 277965 43621
rect 277899 43556 277900 43620
rect 277964 43556 277965 43620
rect 277899 43555 277965 43556
rect 306971 43620 307037 43621
rect 306971 43556 306972 43620
rect 307036 43556 307037 43620
rect 306971 43555 307037 43556
rect 335859 43620 335925 43621
rect 335859 43556 335860 43620
rect 335924 43556 335925 43620
rect 335859 43555 335925 43556
rect 364931 43620 364997 43621
rect 364931 43556 364932 43620
rect 364996 43556 364997 43620
rect 364931 43555 364997 43556
rect 393819 43620 393885 43621
rect 393819 43556 393820 43620
rect 393884 43556 393885 43620
rect 393819 43555 393885 43556
rect 249011 43348 249077 43349
rect 249011 43284 249012 43348
rect 249076 43284 249077 43348
rect 249011 43283 249077 43284
rect 171118 26829 171438 26861
rect 171118 26593 171160 26829
rect 171396 26593 171438 26829
rect 171118 26509 171438 26593
rect 171118 26273 171160 26509
rect 171396 26273 171438 26509
rect 171118 26241 171438 26273
rect 175066 26829 175386 26861
rect 175066 26593 175108 26829
rect 175344 26593 175386 26829
rect 175066 26509 175386 26593
rect 175066 26273 175108 26509
rect 175344 26273 175386 26509
rect 175066 26241 175386 26273
rect 179014 26829 179334 26861
rect 179014 26593 179056 26829
rect 179292 26593 179334 26829
rect 179014 26509 179334 26593
rect 179014 26273 179056 26509
rect 179292 26273 179334 26509
rect 179014 26241 179334 26273
rect 182962 26829 183282 26861
rect 182962 26593 183004 26829
rect 183240 26593 183282 26829
rect 182962 26509 183282 26593
rect 182962 26273 183004 26509
rect 183240 26273 183282 26509
rect 182962 26241 183282 26273
rect 191418 26829 191738 26861
rect 191418 26593 191460 26829
rect 191696 26593 191738 26829
rect 191418 26509 191738 26593
rect 191418 26273 191460 26509
rect 191696 26273 191738 26509
rect 191418 26241 191738 26273
rect 192366 26829 192686 26861
rect 192366 26593 192408 26829
rect 192644 26593 192686 26829
rect 192366 26509 192686 26593
rect 192366 26273 192408 26509
rect 192644 26273 192686 26509
rect 192366 26241 192686 26273
rect 193314 26829 193634 26861
rect 193314 26593 193356 26829
rect 193592 26593 193634 26829
rect 193314 26509 193634 26593
rect 193314 26273 193356 26509
rect 193592 26273 193634 26509
rect 193314 26241 193634 26273
rect 194262 26829 194582 26861
rect 194262 26593 194304 26829
rect 194540 26593 194582 26829
rect 194262 26509 194582 26593
rect 194262 26273 194304 26509
rect 194540 26273 194582 26509
rect 194262 26241 194582 26273
rect 200118 26829 200438 26861
rect 200118 26593 200160 26829
rect 200396 26593 200438 26829
rect 200118 26509 200438 26593
rect 200118 26273 200160 26509
rect 200396 26273 200438 26509
rect 200118 26241 200438 26273
rect 204066 26829 204386 26861
rect 204066 26593 204108 26829
rect 204344 26593 204386 26829
rect 204066 26509 204386 26593
rect 204066 26273 204108 26509
rect 204344 26273 204386 26509
rect 204066 26241 204386 26273
rect 208014 26829 208334 26861
rect 208014 26593 208056 26829
rect 208292 26593 208334 26829
rect 208014 26509 208334 26593
rect 208014 26273 208056 26509
rect 208292 26273 208334 26509
rect 208014 26241 208334 26273
rect 211962 26829 212282 26861
rect 211962 26593 212004 26829
rect 212240 26593 212282 26829
rect 211962 26509 212282 26593
rect 211962 26273 212004 26509
rect 212240 26273 212282 26509
rect 211962 26241 212282 26273
rect 220418 26829 220738 26861
rect 220418 26593 220460 26829
rect 220696 26593 220738 26829
rect 220418 26509 220738 26593
rect 220418 26273 220460 26509
rect 220696 26273 220738 26509
rect 220418 26241 220738 26273
rect 221366 26829 221686 26861
rect 221366 26593 221408 26829
rect 221644 26593 221686 26829
rect 221366 26509 221686 26593
rect 221366 26273 221408 26509
rect 221644 26273 221686 26509
rect 221366 26241 221686 26273
rect 222314 26829 222634 26861
rect 222314 26593 222356 26829
rect 222592 26593 222634 26829
rect 222314 26509 222634 26593
rect 222314 26273 222356 26509
rect 222592 26273 222634 26509
rect 222314 26241 222634 26273
rect 223262 26829 223582 26861
rect 223262 26593 223304 26829
rect 223540 26593 223582 26829
rect 223262 26509 223582 26593
rect 223262 26273 223304 26509
rect 223540 26273 223582 26509
rect 223262 26241 223582 26273
rect 229118 26829 229438 26861
rect 229118 26593 229160 26829
rect 229396 26593 229438 26829
rect 229118 26509 229438 26593
rect 229118 26273 229160 26509
rect 229396 26273 229438 26509
rect 229118 26241 229438 26273
rect 233066 26829 233386 26861
rect 233066 26593 233108 26829
rect 233344 26593 233386 26829
rect 233066 26509 233386 26593
rect 233066 26273 233108 26509
rect 233344 26273 233386 26509
rect 233066 26241 233386 26273
rect 237014 26829 237334 26861
rect 237014 26593 237056 26829
rect 237292 26593 237334 26829
rect 237014 26509 237334 26593
rect 237014 26273 237056 26509
rect 237292 26273 237334 26509
rect 237014 26241 237334 26273
rect 240962 26829 241282 26861
rect 240962 26593 241004 26829
rect 241240 26593 241282 26829
rect 240962 26509 241282 26593
rect 240962 26273 241004 26509
rect 241240 26273 241282 26509
rect 240962 26241 241282 26273
rect 249418 26829 249738 26861
rect 249418 26593 249460 26829
rect 249696 26593 249738 26829
rect 249418 26509 249738 26593
rect 249418 26273 249460 26509
rect 249696 26273 249738 26509
rect 249418 26241 249738 26273
rect 250366 26829 250686 26861
rect 250366 26593 250408 26829
rect 250644 26593 250686 26829
rect 250366 26509 250686 26593
rect 250366 26273 250408 26509
rect 250644 26273 250686 26509
rect 250366 26241 250686 26273
rect 251314 26829 251634 26861
rect 251314 26593 251356 26829
rect 251592 26593 251634 26829
rect 251314 26509 251634 26593
rect 251314 26273 251356 26509
rect 251592 26273 251634 26509
rect 251314 26241 251634 26273
rect 252262 26829 252582 26861
rect 252262 26593 252304 26829
rect 252540 26593 252582 26829
rect 252262 26509 252582 26593
rect 252262 26273 252304 26509
rect 252540 26273 252582 26509
rect 252262 26241 252582 26273
rect 258118 26829 258438 26861
rect 258118 26593 258160 26829
rect 258396 26593 258438 26829
rect 258118 26509 258438 26593
rect 258118 26273 258160 26509
rect 258396 26273 258438 26509
rect 258118 26241 258438 26273
rect 262066 26829 262386 26861
rect 262066 26593 262108 26829
rect 262344 26593 262386 26829
rect 262066 26509 262386 26593
rect 262066 26273 262108 26509
rect 262344 26273 262386 26509
rect 262066 26241 262386 26273
rect 266014 26829 266334 26861
rect 266014 26593 266056 26829
rect 266292 26593 266334 26829
rect 266014 26509 266334 26593
rect 266014 26273 266056 26509
rect 266292 26273 266334 26509
rect 266014 26241 266334 26273
rect 269962 26829 270282 26861
rect 269962 26593 270004 26829
rect 270240 26593 270282 26829
rect 269962 26509 270282 26593
rect 269962 26273 270004 26509
rect 270240 26273 270282 26509
rect 269962 26241 270282 26273
rect 278418 26829 278738 26861
rect 278418 26593 278460 26829
rect 278696 26593 278738 26829
rect 278418 26509 278738 26593
rect 278418 26273 278460 26509
rect 278696 26273 278738 26509
rect 278418 26241 278738 26273
rect 279366 26829 279686 26861
rect 279366 26593 279408 26829
rect 279644 26593 279686 26829
rect 279366 26509 279686 26593
rect 279366 26273 279408 26509
rect 279644 26273 279686 26509
rect 279366 26241 279686 26273
rect 280314 26829 280634 26861
rect 280314 26593 280356 26829
rect 280592 26593 280634 26829
rect 280314 26509 280634 26593
rect 280314 26273 280356 26509
rect 280592 26273 280634 26509
rect 280314 26241 280634 26273
rect 281262 26829 281582 26861
rect 281262 26593 281304 26829
rect 281540 26593 281582 26829
rect 281262 26509 281582 26593
rect 281262 26273 281304 26509
rect 281540 26273 281582 26509
rect 281262 26241 281582 26273
rect 287118 26829 287438 26861
rect 287118 26593 287160 26829
rect 287396 26593 287438 26829
rect 287118 26509 287438 26593
rect 287118 26273 287160 26509
rect 287396 26273 287438 26509
rect 287118 26241 287438 26273
rect 291066 26829 291386 26861
rect 291066 26593 291108 26829
rect 291344 26593 291386 26829
rect 291066 26509 291386 26593
rect 291066 26273 291108 26509
rect 291344 26273 291386 26509
rect 291066 26241 291386 26273
rect 295014 26829 295334 26861
rect 295014 26593 295056 26829
rect 295292 26593 295334 26829
rect 295014 26509 295334 26593
rect 295014 26273 295056 26509
rect 295292 26273 295334 26509
rect 295014 26241 295334 26273
rect 298962 26829 299282 26861
rect 298962 26593 299004 26829
rect 299240 26593 299282 26829
rect 298962 26509 299282 26593
rect 298962 26273 299004 26509
rect 299240 26273 299282 26509
rect 298962 26241 299282 26273
rect 307418 26829 307738 26861
rect 307418 26593 307460 26829
rect 307696 26593 307738 26829
rect 307418 26509 307738 26593
rect 307418 26273 307460 26509
rect 307696 26273 307738 26509
rect 307418 26241 307738 26273
rect 308366 26829 308686 26861
rect 308366 26593 308408 26829
rect 308644 26593 308686 26829
rect 308366 26509 308686 26593
rect 308366 26273 308408 26509
rect 308644 26273 308686 26509
rect 308366 26241 308686 26273
rect 309314 26829 309634 26861
rect 309314 26593 309356 26829
rect 309592 26593 309634 26829
rect 309314 26509 309634 26593
rect 309314 26273 309356 26509
rect 309592 26273 309634 26509
rect 309314 26241 309634 26273
rect 310262 26829 310582 26861
rect 310262 26593 310304 26829
rect 310540 26593 310582 26829
rect 310262 26509 310582 26593
rect 310262 26273 310304 26509
rect 310540 26273 310582 26509
rect 310262 26241 310582 26273
rect 316118 26829 316438 26861
rect 316118 26593 316160 26829
rect 316396 26593 316438 26829
rect 316118 26509 316438 26593
rect 316118 26273 316160 26509
rect 316396 26273 316438 26509
rect 316118 26241 316438 26273
rect 320066 26829 320386 26861
rect 320066 26593 320108 26829
rect 320344 26593 320386 26829
rect 320066 26509 320386 26593
rect 320066 26273 320108 26509
rect 320344 26273 320386 26509
rect 320066 26241 320386 26273
rect 324014 26829 324334 26861
rect 324014 26593 324056 26829
rect 324292 26593 324334 26829
rect 324014 26509 324334 26593
rect 324014 26273 324056 26509
rect 324292 26273 324334 26509
rect 324014 26241 324334 26273
rect 327962 26829 328282 26861
rect 327962 26593 328004 26829
rect 328240 26593 328282 26829
rect 327962 26509 328282 26593
rect 327962 26273 328004 26509
rect 328240 26273 328282 26509
rect 327962 26241 328282 26273
rect 336418 26829 336738 26861
rect 336418 26593 336460 26829
rect 336696 26593 336738 26829
rect 336418 26509 336738 26593
rect 336418 26273 336460 26509
rect 336696 26273 336738 26509
rect 336418 26241 336738 26273
rect 337366 26829 337686 26861
rect 337366 26593 337408 26829
rect 337644 26593 337686 26829
rect 337366 26509 337686 26593
rect 337366 26273 337408 26509
rect 337644 26273 337686 26509
rect 337366 26241 337686 26273
rect 338314 26829 338634 26861
rect 338314 26593 338356 26829
rect 338592 26593 338634 26829
rect 338314 26509 338634 26593
rect 338314 26273 338356 26509
rect 338592 26273 338634 26509
rect 338314 26241 338634 26273
rect 339262 26829 339582 26861
rect 339262 26593 339304 26829
rect 339540 26593 339582 26829
rect 339262 26509 339582 26593
rect 339262 26273 339304 26509
rect 339540 26273 339582 26509
rect 339262 26241 339582 26273
rect 345118 26829 345438 26861
rect 345118 26593 345160 26829
rect 345396 26593 345438 26829
rect 345118 26509 345438 26593
rect 345118 26273 345160 26509
rect 345396 26273 345438 26509
rect 345118 26241 345438 26273
rect 349066 26829 349386 26861
rect 349066 26593 349108 26829
rect 349344 26593 349386 26829
rect 349066 26509 349386 26593
rect 349066 26273 349108 26509
rect 349344 26273 349386 26509
rect 349066 26241 349386 26273
rect 353014 26829 353334 26861
rect 353014 26593 353056 26829
rect 353292 26593 353334 26829
rect 353014 26509 353334 26593
rect 353014 26273 353056 26509
rect 353292 26273 353334 26509
rect 353014 26241 353334 26273
rect 356962 26829 357282 26861
rect 356962 26593 357004 26829
rect 357240 26593 357282 26829
rect 356962 26509 357282 26593
rect 356962 26273 357004 26509
rect 357240 26273 357282 26509
rect 356962 26241 357282 26273
rect 365418 26829 365738 26861
rect 365418 26593 365460 26829
rect 365696 26593 365738 26829
rect 365418 26509 365738 26593
rect 365418 26273 365460 26509
rect 365696 26273 365738 26509
rect 365418 26241 365738 26273
rect 366366 26829 366686 26861
rect 366366 26593 366408 26829
rect 366644 26593 366686 26829
rect 366366 26509 366686 26593
rect 366366 26273 366408 26509
rect 366644 26273 366686 26509
rect 366366 26241 366686 26273
rect 367314 26829 367634 26861
rect 367314 26593 367356 26829
rect 367592 26593 367634 26829
rect 367314 26509 367634 26593
rect 367314 26273 367356 26509
rect 367592 26273 367634 26509
rect 367314 26241 367634 26273
rect 368262 26829 368582 26861
rect 368262 26593 368304 26829
rect 368540 26593 368582 26829
rect 368262 26509 368582 26593
rect 368262 26273 368304 26509
rect 368540 26273 368582 26509
rect 368262 26241 368582 26273
rect 374118 26829 374438 26861
rect 374118 26593 374160 26829
rect 374396 26593 374438 26829
rect 374118 26509 374438 26593
rect 374118 26273 374160 26509
rect 374396 26273 374438 26509
rect 374118 26241 374438 26273
rect 378066 26829 378386 26861
rect 378066 26593 378108 26829
rect 378344 26593 378386 26829
rect 378066 26509 378386 26593
rect 378066 26273 378108 26509
rect 378344 26273 378386 26509
rect 378066 26241 378386 26273
rect 382014 26829 382334 26861
rect 382014 26593 382056 26829
rect 382292 26593 382334 26829
rect 382014 26509 382334 26593
rect 382014 26273 382056 26509
rect 382292 26273 382334 26509
rect 382014 26241 382334 26273
rect 385962 26829 386282 26861
rect 385962 26593 386004 26829
rect 386240 26593 386282 26829
rect 385962 26509 386282 26593
rect 385962 26273 386004 26509
rect 386240 26273 386282 26509
rect 385962 26241 386282 26273
rect 394418 26829 394738 26861
rect 394418 26593 394460 26829
rect 394696 26593 394738 26829
rect 394418 26509 394738 26593
rect 394418 26273 394460 26509
rect 394696 26273 394738 26509
rect 394418 26241 394738 26273
rect 395366 26829 395686 26861
rect 395366 26593 395408 26829
rect 395644 26593 395686 26829
rect 395366 26509 395686 26593
rect 395366 26273 395408 26509
rect 395644 26273 395686 26509
rect 395366 26241 395686 26273
rect 396314 26829 396634 26861
rect 396314 26593 396356 26829
rect 396592 26593 396634 26829
rect 396314 26509 396634 26593
rect 396314 26273 396356 26509
rect 396592 26273 396634 26509
rect 396314 26241 396634 26273
rect 397262 26829 397582 26861
rect 397262 26593 397304 26829
rect 397540 26593 397582 26829
rect 397262 26509 397582 26593
rect 397262 26273 397304 26509
rect 397540 26273 397582 26509
rect 397262 26241 397582 26273
rect 173092 23454 173412 23486
rect 173092 23218 173134 23454
rect 173370 23218 173412 23454
rect 173092 23134 173412 23218
rect 173092 22898 173134 23134
rect 173370 22898 173412 23134
rect 173092 22866 173412 22898
rect 177040 23454 177360 23486
rect 177040 23218 177082 23454
rect 177318 23218 177360 23454
rect 177040 23134 177360 23218
rect 177040 22898 177082 23134
rect 177318 22898 177360 23134
rect 177040 22866 177360 22898
rect 180988 23454 181308 23486
rect 180988 23218 181030 23454
rect 181266 23218 181308 23454
rect 180988 23134 181308 23218
rect 180988 22898 181030 23134
rect 181266 22898 181308 23134
rect 180988 22866 181308 22898
rect 191892 23454 192212 23486
rect 191892 23218 191934 23454
rect 192170 23218 192212 23454
rect 191892 23134 192212 23218
rect 191892 22898 191934 23134
rect 192170 22898 192212 23134
rect 191892 22866 192212 22898
rect 192840 23454 193160 23486
rect 192840 23218 192882 23454
rect 193118 23218 193160 23454
rect 192840 23134 193160 23218
rect 192840 22898 192882 23134
rect 193118 22898 193160 23134
rect 192840 22866 193160 22898
rect 193788 23454 194108 23486
rect 193788 23218 193830 23454
rect 194066 23218 194108 23454
rect 193788 23134 194108 23218
rect 193788 22898 193830 23134
rect 194066 22898 194108 23134
rect 193788 22866 194108 22898
rect 202092 23454 202412 23486
rect 202092 23218 202134 23454
rect 202370 23218 202412 23454
rect 202092 23134 202412 23218
rect 202092 22898 202134 23134
rect 202370 22898 202412 23134
rect 202092 22866 202412 22898
rect 206040 23454 206360 23486
rect 206040 23218 206082 23454
rect 206318 23218 206360 23454
rect 206040 23134 206360 23218
rect 206040 22898 206082 23134
rect 206318 22898 206360 23134
rect 206040 22866 206360 22898
rect 209988 23454 210308 23486
rect 209988 23218 210030 23454
rect 210266 23218 210308 23454
rect 209988 23134 210308 23218
rect 209988 22898 210030 23134
rect 210266 22898 210308 23134
rect 209988 22866 210308 22898
rect 220892 23454 221212 23486
rect 220892 23218 220934 23454
rect 221170 23218 221212 23454
rect 220892 23134 221212 23218
rect 220892 22898 220934 23134
rect 221170 22898 221212 23134
rect 220892 22866 221212 22898
rect 221840 23454 222160 23486
rect 221840 23218 221882 23454
rect 222118 23218 222160 23454
rect 221840 23134 222160 23218
rect 221840 22898 221882 23134
rect 222118 22898 222160 23134
rect 221840 22866 222160 22898
rect 222788 23454 223108 23486
rect 222788 23218 222830 23454
rect 223066 23218 223108 23454
rect 222788 23134 223108 23218
rect 222788 22898 222830 23134
rect 223066 22898 223108 23134
rect 222788 22866 223108 22898
rect 231092 23454 231412 23486
rect 231092 23218 231134 23454
rect 231370 23218 231412 23454
rect 231092 23134 231412 23218
rect 231092 22898 231134 23134
rect 231370 22898 231412 23134
rect 231092 22866 231412 22898
rect 235040 23454 235360 23486
rect 235040 23218 235082 23454
rect 235318 23218 235360 23454
rect 235040 23134 235360 23218
rect 235040 22898 235082 23134
rect 235318 22898 235360 23134
rect 235040 22866 235360 22898
rect 238988 23454 239308 23486
rect 238988 23218 239030 23454
rect 239266 23218 239308 23454
rect 238988 23134 239308 23218
rect 238988 22898 239030 23134
rect 239266 22898 239308 23134
rect 238988 22866 239308 22898
rect 249892 23454 250212 23486
rect 249892 23218 249934 23454
rect 250170 23218 250212 23454
rect 249892 23134 250212 23218
rect 249892 22898 249934 23134
rect 250170 22898 250212 23134
rect 249892 22866 250212 22898
rect 250840 23454 251160 23486
rect 250840 23218 250882 23454
rect 251118 23218 251160 23454
rect 250840 23134 251160 23218
rect 250840 22898 250882 23134
rect 251118 22898 251160 23134
rect 250840 22866 251160 22898
rect 251788 23454 252108 23486
rect 251788 23218 251830 23454
rect 252066 23218 252108 23454
rect 251788 23134 252108 23218
rect 251788 22898 251830 23134
rect 252066 22898 252108 23134
rect 251788 22866 252108 22898
rect 260092 23454 260412 23486
rect 260092 23218 260134 23454
rect 260370 23218 260412 23454
rect 260092 23134 260412 23218
rect 260092 22898 260134 23134
rect 260370 22898 260412 23134
rect 260092 22866 260412 22898
rect 264040 23454 264360 23486
rect 264040 23218 264082 23454
rect 264318 23218 264360 23454
rect 264040 23134 264360 23218
rect 264040 22898 264082 23134
rect 264318 22898 264360 23134
rect 264040 22866 264360 22898
rect 267988 23454 268308 23486
rect 267988 23218 268030 23454
rect 268266 23218 268308 23454
rect 267988 23134 268308 23218
rect 267988 22898 268030 23134
rect 268266 22898 268308 23134
rect 267988 22866 268308 22898
rect 278892 23454 279212 23486
rect 278892 23218 278934 23454
rect 279170 23218 279212 23454
rect 278892 23134 279212 23218
rect 278892 22898 278934 23134
rect 279170 22898 279212 23134
rect 278892 22866 279212 22898
rect 279840 23454 280160 23486
rect 279840 23218 279882 23454
rect 280118 23218 280160 23454
rect 279840 23134 280160 23218
rect 279840 22898 279882 23134
rect 280118 22898 280160 23134
rect 279840 22866 280160 22898
rect 280788 23454 281108 23486
rect 280788 23218 280830 23454
rect 281066 23218 281108 23454
rect 280788 23134 281108 23218
rect 280788 22898 280830 23134
rect 281066 22898 281108 23134
rect 280788 22866 281108 22898
rect 289092 23454 289412 23486
rect 289092 23218 289134 23454
rect 289370 23218 289412 23454
rect 289092 23134 289412 23218
rect 289092 22898 289134 23134
rect 289370 22898 289412 23134
rect 289092 22866 289412 22898
rect 293040 23454 293360 23486
rect 293040 23218 293082 23454
rect 293318 23218 293360 23454
rect 293040 23134 293360 23218
rect 293040 22898 293082 23134
rect 293318 22898 293360 23134
rect 293040 22866 293360 22898
rect 296988 23454 297308 23486
rect 296988 23218 297030 23454
rect 297266 23218 297308 23454
rect 296988 23134 297308 23218
rect 296988 22898 297030 23134
rect 297266 22898 297308 23134
rect 296988 22866 297308 22898
rect 307892 23454 308212 23486
rect 307892 23218 307934 23454
rect 308170 23218 308212 23454
rect 307892 23134 308212 23218
rect 307892 22898 307934 23134
rect 308170 22898 308212 23134
rect 307892 22866 308212 22898
rect 308840 23454 309160 23486
rect 308840 23218 308882 23454
rect 309118 23218 309160 23454
rect 308840 23134 309160 23218
rect 308840 22898 308882 23134
rect 309118 22898 309160 23134
rect 308840 22866 309160 22898
rect 309788 23454 310108 23486
rect 309788 23218 309830 23454
rect 310066 23218 310108 23454
rect 309788 23134 310108 23218
rect 309788 22898 309830 23134
rect 310066 22898 310108 23134
rect 309788 22866 310108 22898
rect 318092 23454 318412 23486
rect 318092 23218 318134 23454
rect 318370 23218 318412 23454
rect 318092 23134 318412 23218
rect 318092 22898 318134 23134
rect 318370 22898 318412 23134
rect 318092 22866 318412 22898
rect 322040 23454 322360 23486
rect 322040 23218 322082 23454
rect 322318 23218 322360 23454
rect 322040 23134 322360 23218
rect 322040 22898 322082 23134
rect 322318 22898 322360 23134
rect 322040 22866 322360 22898
rect 325988 23454 326308 23486
rect 325988 23218 326030 23454
rect 326266 23218 326308 23454
rect 325988 23134 326308 23218
rect 325988 22898 326030 23134
rect 326266 22898 326308 23134
rect 325988 22866 326308 22898
rect 336892 23454 337212 23486
rect 336892 23218 336934 23454
rect 337170 23218 337212 23454
rect 336892 23134 337212 23218
rect 336892 22898 336934 23134
rect 337170 22898 337212 23134
rect 336892 22866 337212 22898
rect 337840 23454 338160 23486
rect 337840 23218 337882 23454
rect 338118 23218 338160 23454
rect 337840 23134 338160 23218
rect 337840 22898 337882 23134
rect 338118 22898 338160 23134
rect 337840 22866 338160 22898
rect 338788 23454 339108 23486
rect 338788 23218 338830 23454
rect 339066 23218 339108 23454
rect 338788 23134 339108 23218
rect 338788 22898 338830 23134
rect 339066 22898 339108 23134
rect 338788 22866 339108 22898
rect 347092 23454 347412 23486
rect 347092 23218 347134 23454
rect 347370 23218 347412 23454
rect 347092 23134 347412 23218
rect 347092 22898 347134 23134
rect 347370 22898 347412 23134
rect 347092 22866 347412 22898
rect 351040 23454 351360 23486
rect 351040 23218 351082 23454
rect 351318 23218 351360 23454
rect 351040 23134 351360 23218
rect 351040 22898 351082 23134
rect 351318 22898 351360 23134
rect 351040 22866 351360 22898
rect 354988 23454 355308 23486
rect 354988 23218 355030 23454
rect 355266 23218 355308 23454
rect 354988 23134 355308 23218
rect 354988 22898 355030 23134
rect 355266 22898 355308 23134
rect 354988 22866 355308 22898
rect 365892 23454 366212 23486
rect 365892 23218 365934 23454
rect 366170 23218 366212 23454
rect 365892 23134 366212 23218
rect 365892 22898 365934 23134
rect 366170 22898 366212 23134
rect 365892 22866 366212 22898
rect 366840 23454 367160 23486
rect 366840 23218 366882 23454
rect 367118 23218 367160 23454
rect 366840 23134 367160 23218
rect 366840 22898 366882 23134
rect 367118 22898 367160 23134
rect 366840 22866 367160 22898
rect 367788 23454 368108 23486
rect 367788 23218 367830 23454
rect 368066 23218 368108 23454
rect 367788 23134 368108 23218
rect 367788 22898 367830 23134
rect 368066 22898 368108 23134
rect 367788 22866 368108 22898
rect 376092 23454 376412 23486
rect 376092 23218 376134 23454
rect 376370 23218 376412 23454
rect 376092 23134 376412 23218
rect 376092 22898 376134 23134
rect 376370 22898 376412 23134
rect 376092 22866 376412 22898
rect 380040 23454 380360 23486
rect 380040 23218 380082 23454
rect 380318 23218 380360 23454
rect 380040 23134 380360 23218
rect 380040 22898 380082 23134
rect 380318 22898 380360 23134
rect 380040 22866 380360 22898
rect 383988 23454 384308 23486
rect 383988 23218 384030 23454
rect 384266 23218 384308 23454
rect 383988 23134 384308 23218
rect 383988 22898 384030 23134
rect 384266 22898 384308 23134
rect 383988 22866 384308 22898
rect 394892 23454 395212 23486
rect 394892 23218 394934 23454
rect 395170 23218 395212 23454
rect 394892 23134 395212 23218
rect 394892 22898 394934 23134
rect 395170 22898 395212 23134
rect 394892 22866 395212 22898
rect 395840 23454 396160 23486
rect 395840 23218 395882 23454
rect 396118 23218 396160 23454
rect 395840 23134 396160 23218
rect 395840 22898 395882 23134
rect 396118 22898 396160 23134
rect 395840 22866 396160 22898
rect 396788 23454 397108 23486
rect 396788 23218 396830 23454
rect 397066 23218 397108 23454
rect 396788 23134 397108 23218
rect 396788 22898 396830 23134
rect 397066 22898 397108 23134
rect 396788 22866 397108 22898
rect 397686 13293 397746 699755
rect 401994 698454 402614 705242
rect 401994 698218 402026 698454
rect 402262 698218 402346 698454
rect 402582 698218 402614 698454
rect 401994 698134 402614 698218
rect 401994 697898 402026 698134
rect 402262 697898 402346 698134
rect 402582 697898 402614 698134
rect 401994 671454 402614 697898
rect 401994 671218 402026 671454
rect 402262 671218 402346 671454
rect 402582 671218 402614 671454
rect 401994 671134 402614 671218
rect 401994 670898 402026 671134
rect 402262 670898 402346 671134
rect 402582 670898 402614 671134
rect 401994 644454 402614 670898
rect 401994 644218 402026 644454
rect 402262 644218 402346 644454
rect 402582 644218 402614 644454
rect 401994 644134 402614 644218
rect 401994 643898 402026 644134
rect 402262 643898 402346 644134
rect 402582 643898 402614 644134
rect 401994 617454 402614 643898
rect 401994 617218 402026 617454
rect 402262 617218 402346 617454
rect 402582 617218 402614 617454
rect 401994 617134 402614 617218
rect 401994 616898 402026 617134
rect 402262 616898 402346 617134
rect 402582 616898 402614 617134
rect 401994 590454 402614 616898
rect 401994 590218 402026 590454
rect 402262 590218 402346 590454
rect 402582 590218 402614 590454
rect 401994 590134 402614 590218
rect 401994 589898 402026 590134
rect 402262 589898 402346 590134
rect 402582 589898 402614 590134
rect 401994 563454 402614 589898
rect 401994 563218 402026 563454
rect 402262 563218 402346 563454
rect 402582 563218 402614 563454
rect 401994 563134 402614 563218
rect 401994 562898 402026 563134
rect 402262 562898 402346 563134
rect 402582 562898 402614 563134
rect 401994 536454 402614 562898
rect 401994 536218 402026 536454
rect 402262 536218 402346 536454
rect 402582 536218 402614 536454
rect 401994 536134 402614 536218
rect 401994 535898 402026 536134
rect 402262 535898 402346 536134
rect 402582 535898 402614 536134
rect 401994 509454 402614 535898
rect 401994 509218 402026 509454
rect 402262 509218 402346 509454
rect 402582 509218 402614 509454
rect 401994 509134 402614 509218
rect 401994 508898 402026 509134
rect 402262 508898 402346 509134
rect 402582 508898 402614 509134
rect 401994 482454 402614 508898
rect 401994 482218 402026 482454
rect 402262 482218 402346 482454
rect 402582 482218 402614 482454
rect 401994 482134 402614 482218
rect 401994 481898 402026 482134
rect 402262 481898 402346 482134
rect 402582 481898 402614 482134
rect 401994 455454 402614 481898
rect 401994 455218 402026 455454
rect 402262 455218 402346 455454
rect 402582 455218 402614 455454
rect 401994 455134 402614 455218
rect 401994 454898 402026 455134
rect 402262 454898 402346 455134
rect 402582 454898 402614 455134
rect 401994 428454 402614 454898
rect 401994 428218 402026 428454
rect 402262 428218 402346 428454
rect 402582 428218 402614 428454
rect 401994 428134 402614 428218
rect 401994 427898 402026 428134
rect 402262 427898 402346 428134
rect 402582 427898 402614 428134
rect 401994 401454 402614 427898
rect 401994 401218 402026 401454
rect 402262 401218 402346 401454
rect 402582 401218 402614 401454
rect 401994 401134 402614 401218
rect 401994 400898 402026 401134
rect 402262 400898 402346 401134
rect 402582 400898 402614 401134
rect 401994 374454 402614 400898
rect 401994 374218 402026 374454
rect 402262 374218 402346 374454
rect 402582 374218 402614 374454
rect 401994 374134 402614 374218
rect 401994 373898 402026 374134
rect 402262 373898 402346 374134
rect 402582 373898 402614 374134
rect 401994 347454 402614 373898
rect 401994 347218 402026 347454
rect 402262 347218 402346 347454
rect 402582 347218 402614 347454
rect 401994 347134 402614 347218
rect 401994 346898 402026 347134
rect 402262 346898 402346 347134
rect 402582 346898 402614 347134
rect 401994 320454 402614 346898
rect 401994 320218 402026 320454
rect 402262 320218 402346 320454
rect 402582 320218 402614 320454
rect 401994 320134 402614 320218
rect 401994 319898 402026 320134
rect 402262 319898 402346 320134
rect 402582 319898 402614 320134
rect 401994 293454 402614 319898
rect 401994 293218 402026 293454
rect 402262 293218 402346 293454
rect 402582 293218 402614 293454
rect 401994 293134 402614 293218
rect 401994 292898 402026 293134
rect 402262 292898 402346 293134
rect 402582 292898 402614 293134
rect 401994 266454 402614 292898
rect 401994 266218 402026 266454
rect 402262 266218 402346 266454
rect 402582 266218 402614 266454
rect 401994 266134 402614 266218
rect 401994 265898 402026 266134
rect 402262 265898 402346 266134
rect 402582 265898 402614 266134
rect 401994 239454 402614 265898
rect 401994 239218 402026 239454
rect 402262 239218 402346 239454
rect 402582 239218 402614 239454
rect 401994 239134 402614 239218
rect 401994 238898 402026 239134
rect 402262 238898 402346 239134
rect 402582 238898 402614 239134
rect 401994 212454 402614 238898
rect 401994 212218 402026 212454
rect 402262 212218 402346 212454
rect 402582 212218 402614 212454
rect 401994 212134 402614 212218
rect 401994 211898 402026 212134
rect 402262 211898 402346 212134
rect 402582 211898 402614 212134
rect 401994 185454 402614 211898
rect 401994 185218 402026 185454
rect 402262 185218 402346 185454
rect 402582 185218 402614 185454
rect 401994 185134 402614 185218
rect 401994 184898 402026 185134
rect 402262 184898 402346 185134
rect 402582 184898 402614 185134
rect 401994 158454 402614 184898
rect 401994 158218 402026 158454
rect 402262 158218 402346 158454
rect 402582 158218 402614 158454
rect 401994 158134 402614 158218
rect 401994 157898 402026 158134
rect 402262 157898 402346 158134
rect 402582 157898 402614 158134
rect 401994 131454 402614 157898
rect 401994 131218 402026 131454
rect 402262 131218 402346 131454
rect 402582 131218 402614 131454
rect 401994 131134 402614 131218
rect 401994 130898 402026 131134
rect 402262 130898 402346 131134
rect 402582 130898 402614 131134
rect 401994 104454 402614 130898
rect 401994 104218 402026 104454
rect 402262 104218 402346 104454
rect 402582 104218 402614 104454
rect 401994 104134 402614 104218
rect 401994 103898 402026 104134
rect 402262 103898 402346 104134
rect 402582 103898 402614 104134
rect 401994 77454 402614 103898
rect 401994 77218 402026 77454
rect 402262 77218 402346 77454
rect 402582 77218 402614 77454
rect 401994 77134 402614 77218
rect 401994 76898 402026 77134
rect 402262 76898 402346 77134
rect 402582 76898 402614 77134
rect 401994 69000 402614 76898
rect 405494 704838 406114 711590
rect 405494 704602 405526 704838
rect 405762 704602 405846 704838
rect 406082 704602 406114 704838
rect 405494 704518 406114 704602
rect 405494 704282 405526 704518
rect 405762 704282 405846 704518
rect 406082 704282 406114 704518
rect 405494 701829 406114 704282
rect 405494 701593 405526 701829
rect 405762 701593 405846 701829
rect 406082 701593 406114 701829
rect 405494 701509 406114 701593
rect 405494 701273 405526 701509
rect 405762 701273 405846 701509
rect 406082 701273 406114 701509
rect 405494 674829 406114 701273
rect 429994 705798 430614 711590
rect 429994 705562 430026 705798
rect 430262 705562 430346 705798
rect 430582 705562 430614 705798
rect 429994 705478 430614 705562
rect 429994 705242 430026 705478
rect 430262 705242 430346 705478
rect 430582 705242 430614 705478
rect 429331 699820 429397 699821
rect 429331 699756 429332 699820
rect 429396 699756 429397 699820
rect 429331 699755 429397 699756
rect 405494 674593 405526 674829
rect 405762 674593 405846 674829
rect 406082 674593 406114 674829
rect 405494 674509 406114 674593
rect 405494 674273 405526 674509
rect 405762 674273 405846 674509
rect 406082 674273 406114 674509
rect 405494 647829 406114 674273
rect 405494 647593 405526 647829
rect 405762 647593 405846 647829
rect 406082 647593 406114 647829
rect 405494 647509 406114 647593
rect 405494 647273 405526 647509
rect 405762 647273 405846 647509
rect 406082 647273 406114 647509
rect 405494 620829 406114 647273
rect 405494 620593 405526 620829
rect 405762 620593 405846 620829
rect 406082 620593 406114 620829
rect 405494 620509 406114 620593
rect 405494 620273 405526 620509
rect 405762 620273 405846 620509
rect 406082 620273 406114 620509
rect 405494 593829 406114 620273
rect 405494 593593 405526 593829
rect 405762 593593 405846 593829
rect 406082 593593 406114 593829
rect 405494 593509 406114 593593
rect 405494 593273 405526 593509
rect 405762 593273 405846 593509
rect 406082 593273 406114 593509
rect 405494 566829 406114 593273
rect 405494 566593 405526 566829
rect 405762 566593 405846 566829
rect 406082 566593 406114 566829
rect 405494 566509 406114 566593
rect 405494 566273 405526 566509
rect 405762 566273 405846 566509
rect 406082 566273 406114 566509
rect 405494 539829 406114 566273
rect 405494 539593 405526 539829
rect 405762 539593 405846 539829
rect 406082 539593 406114 539829
rect 405494 539509 406114 539593
rect 405494 539273 405526 539509
rect 405762 539273 405846 539509
rect 406082 539273 406114 539509
rect 405494 512829 406114 539273
rect 405494 512593 405526 512829
rect 405762 512593 405846 512829
rect 406082 512593 406114 512829
rect 405494 512509 406114 512593
rect 405494 512273 405526 512509
rect 405762 512273 405846 512509
rect 406082 512273 406114 512509
rect 405494 485829 406114 512273
rect 405494 485593 405526 485829
rect 405762 485593 405846 485829
rect 406082 485593 406114 485829
rect 405494 485509 406114 485593
rect 405494 485273 405526 485509
rect 405762 485273 405846 485509
rect 406082 485273 406114 485509
rect 405494 458829 406114 485273
rect 405494 458593 405526 458829
rect 405762 458593 405846 458829
rect 406082 458593 406114 458829
rect 405494 458509 406114 458593
rect 405494 458273 405526 458509
rect 405762 458273 405846 458509
rect 406082 458273 406114 458509
rect 405494 431829 406114 458273
rect 405494 431593 405526 431829
rect 405762 431593 405846 431829
rect 406082 431593 406114 431829
rect 405494 431509 406114 431593
rect 405494 431273 405526 431509
rect 405762 431273 405846 431509
rect 406082 431273 406114 431509
rect 405494 404829 406114 431273
rect 405494 404593 405526 404829
rect 405762 404593 405846 404829
rect 406082 404593 406114 404829
rect 405494 404509 406114 404593
rect 405494 404273 405526 404509
rect 405762 404273 405846 404509
rect 406082 404273 406114 404509
rect 405494 377829 406114 404273
rect 405494 377593 405526 377829
rect 405762 377593 405846 377829
rect 406082 377593 406114 377829
rect 405494 377509 406114 377593
rect 405494 377273 405526 377509
rect 405762 377273 405846 377509
rect 406082 377273 406114 377509
rect 405494 350829 406114 377273
rect 405494 350593 405526 350829
rect 405762 350593 405846 350829
rect 406082 350593 406114 350829
rect 405494 350509 406114 350593
rect 405494 350273 405526 350509
rect 405762 350273 405846 350509
rect 406082 350273 406114 350509
rect 405494 323829 406114 350273
rect 405494 323593 405526 323829
rect 405762 323593 405846 323829
rect 406082 323593 406114 323829
rect 405494 323509 406114 323593
rect 405494 323273 405526 323509
rect 405762 323273 405846 323509
rect 406082 323273 406114 323509
rect 405494 296829 406114 323273
rect 405494 296593 405526 296829
rect 405762 296593 405846 296829
rect 406082 296593 406114 296829
rect 405494 296509 406114 296593
rect 405494 296273 405526 296509
rect 405762 296273 405846 296509
rect 406082 296273 406114 296509
rect 405494 269829 406114 296273
rect 405494 269593 405526 269829
rect 405762 269593 405846 269829
rect 406082 269593 406114 269829
rect 405494 269509 406114 269593
rect 405494 269273 405526 269509
rect 405762 269273 405846 269509
rect 406082 269273 406114 269509
rect 405494 242829 406114 269273
rect 405494 242593 405526 242829
rect 405762 242593 405846 242829
rect 406082 242593 406114 242829
rect 405494 242509 406114 242593
rect 405494 242273 405526 242509
rect 405762 242273 405846 242509
rect 406082 242273 406114 242509
rect 405494 215829 406114 242273
rect 405494 215593 405526 215829
rect 405762 215593 405846 215829
rect 406082 215593 406114 215829
rect 405494 215509 406114 215593
rect 405494 215273 405526 215509
rect 405762 215273 405846 215509
rect 406082 215273 406114 215509
rect 405494 188829 406114 215273
rect 405494 188593 405526 188829
rect 405762 188593 405846 188829
rect 406082 188593 406114 188829
rect 405494 188509 406114 188593
rect 405494 188273 405526 188509
rect 405762 188273 405846 188509
rect 406082 188273 406114 188509
rect 405494 161829 406114 188273
rect 405494 161593 405526 161829
rect 405762 161593 405846 161829
rect 406082 161593 406114 161829
rect 405494 161509 406114 161593
rect 405494 161273 405526 161509
rect 405762 161273 405846 161509
rect 406082 161273 406114 161509
rect 405494 134829 406114 161273
rect 405494 134593 405526 134829
rect 405762 134593 405846 134829
rect 406082 134593 406114 134829
rect 405494 134509 406114 134593
rect 405494 134273 405526 134509
rect 405762 134273 405846 134509
rect 406082 134273 406114 134509
rect 405494 107829 406114 134273
rect 405494 107593 405526 107829
rect 405762 107593 405846 107829
rect 406082 107593 406114 107829
rect 405494 107509 406114 107593
rect 405494 107273 405526 107509
rect 405762 107273 405846 107509
rect 406082 107273 406114 107509
rect 405494 80829 406114 107273
rect 405494 80593 405526 80829
rect 405762 80593 405846 80829
rect 406082 80593 406114 80829
rect 405494 80509 406114 80593
rect 405494 80273 405526 80509
rect 405762 80273 405846 80509
rect 406082 80273 406114 80509
rect 405494 69000 406114 80273
rect 422891 65652 422957 65653
rect 422891 65588 422892 65652
rect 422956 65588 422957 65652
rect 422891 65587 422957 65588
rect 399866 53829 400186 53861
rect 399866 53593 399908 53829
rect 400144 53593 400186 53829
rect 399866 53509 400186 53593
rect 399866 53273 399908 53509
rect 400144 53273 400186 53509
rect 399866 53241 400186 53273
rect 403814 53829 404134 53861
rect 403814 53593 403856 53829
rect 404092 53593 404134 53829
rect 403814 53509 404134 53593
rect 403814 53273 403856 53509
rect 404092 53273 404134 53509
rect 403814 53241 404134 53273
rect 407762 53829 408082 53861
rect 407762 53593 407804 53829
rect 408040 53593 408082 53829
rect 407762 53509 408082 53593
rect 407762 53273 407804 53509
rect 408040 53273 408082 53509
rect 407762 53241 408082 53273
rect 416218 53829 416538 53861
rect 416218 53593 416260 53829
rect 416496 53593 416538 53829
rect 416218 53509 416538 53593
rect 416218 53273 416260 53509
rect 416496 53273 416538 53509
rect 416218 53241 416538 53273
rect 417166 53829 417486 53861
rect 417166 53593 417208 53829
rect 417444 53593 417486 53829
rect 417166 53509 417486 53593
rect 417166 53273 417208 53509
rect 417444 53273 417486 53509
rect 417166 53241 417486 53273
rect 418114 53829 418434 53861
rect 418114 53593 418156 53829
rect 418392 53593 418434 53829
rect 418114 53509 418434 53593
rect 418114 53273 418156 53509
rect 418392 53273 418434 53509
rect 418114 53241 418434 53273
rect 419062 53829 419382 53861
rect 419062 53593 419104 53829
rect 419340 53593 419382 53829
rect 419062 53509 419382 53593
rect 419062 53273 419104 53509
rect 419340 53273 419382 53509
rect 419062 53241 419382 53273
rect 397892 50454 398212 50486
rect 397892 50218 397934 50454
rect 398170 50218 398212 50454
rect 397892 50134 398212 50218
rect 397892 49898 397934 50134
rect 398170 49898 398212 50134
rect 397892 49866 398212 49898
rect 401840 50454 402160 50486
rect 401840 50218 401882 50454
rect 402118 50218 402160 50454
rect 401840 50134 402160 50218
rect 401840 49898 401882 50134
rect 402118 49898 402160 50134
rect 401840 49866 402160 49898
rect 405788 50454 406108 50486
rect 405788 50218 405830 50454
rect 406066 50218 406108 50454
rect 405788 50134 406108 50218
rect 405788 49898 405830 50134
rect 406066 49898 406108 50134
rect 405788 49866 406108 49898
rect 416692 50454 417012 50486
rect 416692 50218 416734 50454
rect 416970 50218 417012 50454
rect 416692 50134 417012 50218
rect 416692 49898 416734 50134
rect 416970 49898 417012 50134
rect 416692 49866 417012 49898
rect 417640 50454 417960 50486
rect 417640 50218 417682 50454
rect 417918 50218 417960 50454
rect 417640 50134 417960 50218
rect 417640 49898 417682 50134
rect 417918 49898 417960 50134
rect 417640 49866 417960 49898
rect 418588 50454 418908 50486
rect 418588 50218 418630 50454
rect 418866 50218 418908 50454
rect 418588 50134 418908 50218
rect 418588 49898 418630 50134
rect 418866 49898 418908 50134
rect 418588 49866 418908 49898
rect 422894 43621 422954 65587
rect 424918 53829 425238 53861
rect 424918 53593 424960 53829
rect 425196 53593 425238 53829
rect 424918 53509 425238 53593
rect 424918 53273 424960 53509
rect 425196 53273 425238 53509
rect 424918 53241 425238 53273
rect 428866 53829 429186 53861
rect 428866 53593 428908 53829
rect 429144 53593 429186 53829
rect 428866 53509 429186 53593
rect 428866 53273 428908 53509
rect 429144 53273 429186 53509
rect 428866 53241 429186 53273
rect 426892 50454 427212 50486
rect 426892 50218 426934 50454
rect 427170 50218 427212 50454
rect 426892 50134 427212 50218
rect 426892 49898 426934 50134
rect 427170 49898 427212 50134
rect 426892 49866 427212 49898
rect 422891 43620 422957 43621
rect 422891 43556 422892 43620
rect 422956 43556 422957 43620
rect 422891 43555 422957 43556
rect 403118 26829 403438 26861
rect 403118 26593 403160 26829
rect 403396 26593 403438 26829
rect 403118 26509 403438 26593
rect 403118 26273 403160 26509
rect 403396 26273 403438 26509
rect 403118 26241 403438 26273
rect 407066 26829 407386 26861
rect 407066 26593 407108 26829
rect 407344 26593 407386 26829
rect 407066 26509 407386 26593
rect 407066 26273 407108 26509
rect 407344 26273 407386 26509
rect 407066 26241 407386 26273
rect 411014 26829 411334 26861
rect 411014 26593 411056 26829
rect 411292 26593 411334 26829
rect 411014 26509 411334 26593
rect 411014 26273 411056 26509
rect 411292 26273 411334 26509
rect 411014 26241 411334 26273
rect 414962 26829 415282 26861
rect 414962 26593 415004 26829
rect 415240 26593 415282 26829
rect 414962 26509 415282 26593
rect 414962 26273 415004 26509
rect 415240 26273 415282 26509
rect 414962 26241 415282 26273
rect 423418 26829 423738 26861
rect 423418 26593 423460 26829
rect 423696 26593 423738 26829
rect 423418 26509 423738 26593
rect 423418 26273 423460 26509
rect 423696 26273 423738 26509
rect 423418 26241 423738 26273
rect 424366 26829 424686 26861
rect 424366 26593 424408 26829
rect 424644 26593 424686 26829
rect 424366 26509 424686 26593
rect 424366 26273 424408 26509
rect 424644 26273 424686 26509
rect 424366 26241 424686 26273
rect 425314 26829 425634 26861
rect 425314 26593 425356 26829
rect 425592 26593 425634 26829
rect 425314 26509 425634 26593
rect 425314 26273 425356 26509
rect 425592 26273 425634 26509
rect 425314 26241 425634 26273
rect 426262 26829 426582 26861
rect 426262 26593 426304 26829
rect 426540 26593 426582 26829
rect 426262 26509 426582 26593
rect 426262 26273 426304 26509
rect 426540 26273 426582 26509
rect 426262 26241 426582 26273
rect 405092 23454 405412 23486
rect 405092 23218 405134 23454
rect 405370 23218 405412 23454
rect 405092 23134 405412 23218
rect 405092 22898 405134 23134
rect 405370 22898 405412 23134
rect 405092 22866 405412 22898
rect 409040 23454 409360 23486
rect 409040 23218 409082 23454
rect 409318 23218 409360 23454
rect 409040 23134 409360 23218
rect 409040 22898 409082 23134
rect 409318 22898 409360 23134
rect 409040 22866 409360 22898
rect 412988 23454 413308 23486
rect 412988 23218 413030 23454
rect 413266 23218 413308 23454
rect 412988 23134 413308 23218
rect 412988 22898 413030 23134
rect 413266 22898 413308 23134
rect 412988 22866 413308 22898
rect 423892 23454 424212 23486
rect 423892 23218 423934 23454
rect 424170 23218 424212 23454
rect 423892 23134 424212 23218
rect 423892 22898 423934 23134
rect 424170 22898 424212 23134
rect 423892 22866 424212 22898
rect 424840 23454 425160 23486
rect 424840 23218 424882 23454
rect 425118 23218 425160 23454
rect 424840 23134 425160 23218
rect 424840 22898 424882 23134
rect 425118 22898 425160 23134
rect 424840 22866 425160 22898
rect 425788 23454 426108 23486
rect 425788 23218 425830 23454
rect 426066 23218 426108 23454
rect 425788 23134 426108 23218
rect 425788 22898 425830 23134
rect 426066 22898 426108 23134
rect 425788 22866 426108 22898
rect 429334 13429 429394 699755
rect 429994 698454 430614 705242
rect 429994 698218 430026 698454
rect 430262 698218 430346 698454
rect 430582 698218 430614 698454
rect 429994 698134 430614 698218
rect 429994 697898 430026 698134
rect 430262 697898 430346 698134
rect 430582 697898 430614 698134
rect 429994 671454 430614 697898
rect 429994 671218 430026 671454
rect 430262 671218 430346 671454
rect 430582 671218 430614 671454
rect 429994 671134 430614 671218
rect 429994 670898 430026 671134
rect 430262 670898 430346 671134
rect 430582 670898 430614 671134
rect 429994 644454 430614 670898
rect 429994 644218 430026 644454
rect 430262 644218 430346 644454
rect 430582 644218 430614 644454
rect 429994 644134 430614 644218
rect 429994 643898 430026 644134
rect 430262 643898 430346 644134
rect 430582 643898 430614 644134
rect 429994 617454 430614 643898
rect 429994 617218 430026 617454
rect 430262 617218 430346 617454
rect 430582 617218 430614 617454
rect 429994 617134 430614 617218
rect 429994 616898 430026 617134
rect 430262 616898 430346 617134
rect 430582 616898 430614 617134
rect 429994 590454 430614 616898
rect 429994 590218 430026 590454
rect 430262 590218 430346 590454
rect 430582 590218 430614 590454
rect 429994 590134 430614 590218
rect 429994 589898 430026 590134
rect 430262 589898 430346 590134
rect 430582 589898 430614 590134
rect 429994 563454 430614 589898
rect 429994 563218 430026 563454
rect 430262 563218 430346 563454
rect 430582 563218 430614 563454
rect 429994 563134 430614 563218
rect 429994 562898 430026 563134
rect 430262 562898 430346 563134
rect 430582 562898 430614 563134
rect 429994 536454 430614 562898
rect 429994 536218 430026 536454
rect 430262 536218 430346 536454
rect 430582 536218 430614 536454
rect 429994 536134 430614 536218
rect 429994 535898 430026 536134
rect 430262 535898 430346 536134
rect 430582 535898 430614 536134
rect 429994 509454 430614 535898
rect 429994 509218 430026 509454
rect 430262 509218 430346 509454
rect 430582 509218 430614 509454
rect 429994 509134 430614 509218
rect 429994 508898 430026 509134
rect 430262 508898 430346 509134
rect 430582 508898 430614 509134
rect 429994 482454 430614 508898
rect 429994 482218 430026 482454
rect 430262 482218 430346 482454
rect 430582 482218 430614 482454
rect 429994 482134 430614 482218
rect 429994 481898 430026 482134
rect 430262 481898 430346 482134
rect 430582 481898 430614 482134
rect 429994 455454 430614 481898
rect 429994 455218 430026 455454
rect 430262 455218 430346 455454
rect 430582 455218 430614 455454
rect 429994 455134 430614 455218
rect 429994 454898 430026 455134
rect 430262 454898 430346 455134
rect 430582 454898 430614 455134
rect 429994 428454 430614 454898
rect 429994 428218 430026 428454
rect 430262 428218 430346 428454
rect 430582 428218 430614 428454
rect 429994 428134 430614 428218
rect 429994 427898 430026 428134
rect 430262 427898 430346 428134
rect 430582 427898 430614 428134
rect 429994 401454 430614 427898
rect 429994 401218 430026 401454
rect 430262 401218 430346 401454
rect 430582 401218 430614 401454
rect 429994 401134 430614 401218
rect 429994 400898 430026 401134
rect 430262 400898 430346 401134
rect 430582 400898 430614 401134
rect 429994 374454 430614 400898
rect 429994 374218 430026 374454
rect 430262 374218 430346 374454
rect 430582 374218 430614 374454
rect 429994 374134 430614 374218
rect 429994 373898 430026 374134
rect 430262 373898 430346 374134
rect 430582 373898 430614 374134
rect 429994 347454 430614 373898
rect 429994 347218 430026 347454
rect 430262 347218 430346 347454
rect 430582 347218 430614 347454
rect 429994 347134 430614 347218
rect 429994 346898 430026 347134
rect 430262 346898 430346 347134
rect 430582 346898 430614 347134
rect 429994 320454 430614 346898
rect 429994 320218 430026 320454
rect 430262 320218 430346 320454
rect 430582 320218 430614 320454
rect 429994 320134 430614 320218
rect 429994 319898 430026 320134
rect 430262 319898 430346 320134
rect 430582 319898 430614 320134
rect 429994 293454 430614 319898
rect 429994 293218 430026 293454
rect 430262 293218 430346 293454
rect 430582 293218 430614 293454
rect 429994 293134 430614 293218
rect 429994 292898 430026 293134
rect 430262 292898 430346 293134
rect 430582 292898 430614 293134
rect 429994 266454 430614 292898
rect 429994 266218 430026 266454
rect 430262 266218 430346 266454
rect 430582 266218 430614 266454
rect 429994 266134 430614 266218
rect 429994 265898 430026 266134
rect 430262 265898 430346 266134
rect 430582 265898 430614 266134
rect 429994 239454 430614 265898
rect 429994 239218 430026 239454
rect 430262 239218 430346 239454
rect 430582 239218 430614 239454
rect 429994 239134 430614 239218
rect 429994 238898 430026 239134
rect 430262 238898 430346 239134
rect 430582 238898 430614 239134
rect 429994 212454 430614 238898
rect 429994 212218 430026 212454
rect 430262 212218 430346 212454
rect 430582 212218 430614 212454
rect 429994 212134 430614 212218
rect 429994 211898 430026 212134
rect 430262 211898 430346 212134
rect 430582 211898 430614 212134
rect 429994 185454 430614 211898
rect 429994 185218 430026 185454
rect 430262 185218 430346 185454
rect 430582 185218 430614 185454
rect 429994 185134 430614 185218
rect 429994 184898 430026 185134
rect 430262 184898 430346 185134
rect 430582 184898 430614 185134
rect 429994 158454 430614 184898
rect 429994 158218 430026 158454
rect 430262 158218 430346 158454
rect 430582 158218 430614 158454
rect 429994 158134 430614 158218
rect 429994 157898 430026 158134
rect 430262 157898 430346 158134
rect 430582 157898 430614 158134
rect 429994 131454 430614 157898
rect 429994 131218 430026 131454
rect 430262 131218 430346 131454
rect 430582 131218 430614 131454
rect 429994 131134 430614 131218
rect 429994 130898 430026 131134
rect 430262 130898 430346 131134
rect 430582 130898 430614 131134
rect 429994 104454 430614 130898
rect 429994 104218 430026 104454
rect 430262 104218 430346 104454
rect 430582 104218 430614 104454
rect 429994 104134 430614 104218
rect 429994 103898 430026 104134
rect 430262 103898 430346 104134
rect 430582 103898 430614 104134
rect 429994 77454 430614 103898
rect 429994 77218 430026 77454
rect 430262 77218 430346 77454
rect 430582 77218 430614 77454
rect 429994 77134 430614 77218
rect 429994 76898 430026 77134
rect 430262 76898 430346 77134
rect 430582 76898 430614 77134
rect 429994 69000 430614 76898
rect 433494 704838 434114 711590
rect 433494 704602 433526 704838
rect 433762 704602 433846 704838
rect 434082 704602 434114 704838
rect 433494 704518 434114 704602
rect 433494 704282 433526 704518
rect 433762 704282 433846 704518
rect 434082 704282 434114 704518
rect 433494 701829 434114 704282
rect 433494 701593 433526 701829
rect 433762 701593 433846 701829
rect 434082 701593 434114 701829
rect 433494 701509 434114 701593
rect 433494 701273 433526 701509
rect 433762 701273 433846 701509
rect 434082 701273 434114 701509
rect 433494 674829 434114 701273
rect 433494 674593 433526 674829
rect 433762 674593 433846 674829
rect 434082 674593 434114 674829
rect 433494 674509 434114 674593
rect 433494 674273 433526 674509
rect 433762 674273 433846 674509
rect 434082 674273 434114 674509
rect 433494 647829 434114 674273
rect 433494 647593 433526 647829
rect 433762 647593 433846 647829
rect 434082 647593 434114 647829
rect 433494 647509 434114 647593
rect 433494 647273 433526 647509
rect 433762 647273 433846 647509
rect 434082 647273 434114 647509
rect 433494 620829 434114 647273
rect 433494 620593 433526 620829
rect 433762 620593 433846 620829
rect 434082 620593 434114 620829
rect 433494 620509 434114 620593
rect 433494 620273 433526 620509
rect 433762 620273 433846 620509
rect 434082 620273 434114 620509
rect 433494 593829 434114 620273
rect 433494 593593 433526 593829
rect 433762 593593 433846 593829
rect 434082 593593 434114 593829
rect 433494 593509 434114 593593
rect 433494 593273 433526 593509
rect 433762 593273 433846 593509
rect 434082 593273 434114 593509
rect 433494 566829 434114 593273
rect 433494 566593 433526 566829
rect 433762 566593 433846 566829
rect 434082 566593 434114 566829
rect 433494 566509 434114 566593
rect 433494 566273 433526 566509
rect 433762 566273 433846 566509
rect 434082 566273 434114 566509
rect 433494 539829 434114 566273
rect 433494 539593 433526 539829
rect 433762 539593 433846 539829
rect 434082 539593 434114 539829
rect 433494 539509 434114 539593
rect 433494 539273 433526 539509
rect 433762 539273 433846 539509
rect 434082 539273 434114 539509
rect 433494 512829 434114 539273
rect 433494 512593 433526 512829
rect 433762 512593 433846 512829
rect 434082 512593 434114 512829
rect 433494 512509 434114 512593
rect 433494 512273 433526 512509
rect 433762 512273 433846 512509
rect 434082 512273 434114 512509
rect 433494 485829 434114 512273
rect 433494 485593 433526 485829
rect 433762 485593 433846 485829
rect 434082 485593 434114 485829
rect 433494 485509 434114 485593
rect 433494 485273 433526 485509
rect 433762 485273 433846 485509
rect 434082 485273 434114 485509
rect 433494 458829 434114 485273
rect 433494 458593 433526 458829
rect 433762 458593 433846 458829
rect 434082 458593 434114 458829
rect 433494 458509 434114 458593
rect 433494 458273 433526 458509
rect 433762 458273 433846 458509
rect 434082 458273 434114 458509
rect 433494 431829 434114 458273
rect 433494 431593 433526 431829
rect 433762 431593 433846 431829
rect 434082 431593 434114 431829
rect 433494 431509 434114 431593
rect 433494 431273 433526 431509
rect 433762 431273 433846 431509
rect 434082 431273 434114 431509
rect 433494 404829 434114 431273
rect 433494 404593 433526 404829
rect 433762 404593 433846 404829
rect 434082 404593 434114 404829
rect 433494 404509 434114 404593
rect 433494 404273 433526 404509
rect 433762 404273 433846 404509
rect 434082 404273 434114 404509
rect 433494 377829 434114 404273
rect 433494 377593 433526 377829
rect 433762 377593 433846 377829
rect 434082 377593 434114 377829
rect 433494 377509 434114 377593
rect 433494 377273 433526 377509
rect 433762 377273 433846 377509
rect 434082 377273 434114 377509
rect 433494 350829 434114 377273
rect 433494 350593 433526 350829
rect 433762 350593 433846 350829
rect 434082 350593 434114 350829
rect 433494 350509 434114 350593
rect 433494 350273 433526 350509
rect 433762 350273 433846 350509
rect 434082 350273 434114 350509
rect 433494 323829 434114 350273
rect 433494 323593 433526 323829
rect 433762 323593 433846 323829
rect 434082 323593 434114 323829
rect 433494 323509 434114 323593
rect 433494 323273 433526 323509
rect 433762 323273 433846 323509
rect 434082 323273 434114 323509
rect 433494 296829 434114 323273
rect 433494 296593 433526 296829
rect 433762 296593 433846 296829
rect 434082 296593 434114 296829
rect 433494 296509 434114 296593
rect 433494 296273 433526 296509
rect 433762 296273 433846 296509
rect 434082 296273 434114 296509
rect 433494 269829 434114 296273
rect 433494 269593 433526 269829
rect 433762 269593 433846 269829
rect 434082 269593 434114 269829
rect 433494 269509 434114 269593
rect 433494 269273 433526 269509
rect 433762 269273 433846 269509
rect 434082 269273 434114 269509
rect 433494 242829 434114 269273
rect 433494 242593 433526 242829
rect 433762 242593 433846 242829
rect 434082 242593 434114 242829
rect 433494 242509 434114 242593
rect 433494 242273 433526 242509
rect 433762 242273 433846 242509
rect 434082 242273 434114 242509
rect 433494 215829 434114 242273
rect 433494 215593 433526 215829
rect 433762 215593 433846 215829
rect 434082 215593 434114 215829
rect 433494 215509 434114 215593
rect 433494 215273 433526 215509
rect 433762 215273 433846 215509
rect 434082 215273 434114 215509
rect 433494 188829 434114 215273
rect 433494 188593 433526 188829
rect 433762 188593 433846 188829
rect 434082 188593 434114 188829
rect 433494 188509 434114 188593
rect 433494 188273 433526 188509
rect 433762 188273 433846 188509
rect 434082 188273 434114 188509
rect 433494 161829 434114 188273
rect 433494 161593 433526 161829
rect 433762 161593 433846 161829
rect 434082 161593 434114 161829
rect 433494 161509 434114 161593
rect 433494 161273 433526 161509
rect 433762 161273 433846 161509
rect 434082 161273 434114 161509
rect 433494 134829 434114 161273
rect 433494 134593 433526 134829
rect 433762 134593 433846 134829
rect 434082 134593 434114 134829
rect 433494 134509 434114 134593
rect 433494 134273 433526 134509
rect 433762 134273 433846 134509
rect 434082 134273 434114 134509
rect 433494 107829 434114 134273
rect 433494 107593 433526 107829
rect 433762 107593 433846 107829
rect 434082 107593 434114 107829
rect 433494 107509 434114 107593
rect 433494 107273 433526 107509
rect 433762 107273 433846 107509
rect 434082 107273 434114 107509
rect 433494 80829 434114 107273
rect 433494 80593 433526 80829
rect 433762 80593 433846 80829
rect 434082 80593 434114 80829
rect 433494 80509 434114 80593
rect 433494 80273 433526 80509
rect 433762 80273 433846 80509
rect 434082 80273 434114 80509
rect 433494 69000 434114 80273
rect 457994 705798 458614 711590
rect 457994 705562 458026 705798
rect 458262 705562 458346 705798
rect 458582 705562 458614 705798
rect 457994 705478 458614 705562
rect 457994 705242 458026 705478
rect 458262 705242 458346 705478
rect 458582 705242 458614 705478
rect 457994 698454 458614 705242
rect 457994 698218 458026 698454
rect 458262 698218 458346 698454
rect 458582 698218 458614 698454
rect 457994 698134 458614 698218
rect 457994 697898 458026 698134
rect 458262 697898 458346 698134
rect 458582 697898 458614 698134
rect 457994 671454 458614 697898
rect 457994 671218 458026 671454
rect 458262 671218 458346 671454
rect 458582 671218 458614 671454
rect 457994 671134 458614 671218
rect 457994 670898 458026 671134
rect 458262 670898 458346 671134
rect 458582 670898 458614 671134
rect 457994 644454 458614 670898
rect 457994 644218 458026 644454
rect 458262 644218 458346 644454
rect 458582 644218 458614 644454
rect 457994 644134 458614 644218
rect 457994 643898 458026 644134
rect 458262 643898 458346 644134
rect 458582 643898 458614 644134
rect 457994 617454 458614 643898
rect 457994 617218 458026 617454
rect 458262 617218 458346 617454
rect 458582 617218 458614 617454
rect 457994 617134 458614 617218
rect 457994 616898 458026 617134
rect 458262 616898 458346 617134
rect 458582 616898 458614 617134
rect 457994 590454 458614 616898
rect 457994 590218 458026 590454
rect 458262 590218 458346 590454
rect 458582 590218 458614 590454
rect 457994 590134 458614 590218
rect 457994 589898 458026 590134
rect 458262 589898 458346 590134
rect 458582 589898 458614 590134
rect 457994 563454 458614 589898
rect 457994 563218 458026 563454
rect 458262 563218 458346 563454
rect 458582 563218 458614 563454
rect 457994 563134 458614 563218
rect 457994 562898 458026 563134
rect 458262 562898 458346 563134
rect 458582 562898 458614 563134
rect 457994 536454 458614 562898
rect 457994 536218 458026 536454
rect 458262 536218 458346 536454
rect 458582 536218 458614 536454
rect 457994 536134 458614 536218
rect 457994 535898 458026 536134
rect 458262 535898 458346 536134
rect 458582 535898 458614 536134
rect 457994 509454 458614 535898
rect 457994 509218 458026 509454
rect 458262 509218 458346 509454
rect 458582 509218 458614 509454
rect 457994 509134 458614 509218
rect 457994 508898 458026 509134
rect 458262 508898 458346 509134
rect 458582 508898 458614 509134
rect 457994 482454 458614 508898
rect 457994 482218 458026 482454
rect 458262 482218 458346 482454
rect 458582 482218 458614 482454
rect 457994 482134 458614 482218
rect 457994 481898 458026 482134
rect 458262 481898 458346 482134
rect 458582 481898 458614 482134
rect 457994 455454 458614 481898
rect 457994 455218 458026 455454
rect 458262 455218 458346 455454
rect 458582 455218 458614 455454
rect 457994 455134 458614 455218
rect 457994 454898 458026 455134
rect 458262 454898 458346 455134
rect 458582 454898 458614 455134
rect 457994 428454 458614 454898
rect 457994 428218 458026 428454
rect 458262 428218 458346 428454
rect 458582 428218 458614 428454
rect 457994 428134 458614 428218
rect 457994 427898 458026 428134
rect 458262 427898 458346 428134
rect 458582 427898 458614 428134
rect 457994 401454 458614 427898
rect 457994 401218 458026 401454
rect 458262 401218 458346 401454
rect 458582 401218 458614 401454
rect 457994 401134 458614 401218
rect 457994 400898 458026 401134
rect 458262 400898 458346 401134
rect 458582 400898 458614 401134
rect 457994 374454 458614 400898
rect 457994 374218 458026 374454
rect 458262 374218 458346 374454
rect 458582 374218 458614 374454
rect 457994 374134 458614 374218
rect 457994 373898 458026 374134
rect 458262 373898 458346 374134
rect 458582 373898 458614 374134
rect 457994 347454 458614 373898
rect 457994 347218 458026 347454
rect 458262 347218 458346 347454
rect 458582 347218 458614 347454
rect 457994 347134 458614 347218
rect 457994 346898 458026 347134
rect 458262 346898 458346 347134
rect 458582 346898 458614 347134
rect 457994 320454 458614 346898
rect 457994 320218 458026 320454
rect 458262 320218 458346 320454
rect 458582 320218 458614 320454
rect 457994 320134 458614 320218
rect 457994 319898 458026 320134
rect 458262 319898 458346 320134
rect 458582 319898 458614 320134
rect 457994 293454 458614 319898
rect 457994 293218 458026 293454
rect 458262 293218 458346 293454
rect 458582 293218 458614 293454
rect 457994 293134 458614 293218
rect 457994 292898 458026 293134
rect 458262 292898 458346 293134
rect 458582 292898 458614 293134
rect 457994 266454 458614 292898
rect 457994 266218 458026 266454
rect 458262 266218 458346 266454
rect 458582 266218 458614 266454
rect 457994 266134 458614 266218
rect 457994 265898 458026 266134
rect 458262 265898 458346 266134
rect 458582 265898 458614 266134
rect 457994 239454 458614 265898
rect 457994 239218 458026 239454
rect 458262 239218 458346 239454
rect 458582 239218 458614 239454
rect 457994 239134 458614 239218
rect 457994 238898 458026 239134
rect 458262 238898 458346 239134
rect 458582 238898 458614 239134
rect 457994 212454 458614 238898
rect 457994 212218 458026 212454
rect 458262 212218 458346 212454
rect 458582 212218 458614 212454
rect 457994 212134 458614 212218
rect 457994 211898 458026 212134
rect 458262 211898 458346 212134
rect 458582 211898 458614 212134
rect 457994 185454 458614 211898
rect 457994 185218 458026 185454
rect 458262 185218 458346 185454
rect 458582 185218 458614 185454
rect 457994 185134 458614 185218
rect 457994 184898 458026 185134
rect 458262 184898 458346 185134
rect 458582 184898 458614 185134
rect 457994 158454 458614 184898
rect 457994 158218 458026 158454
rect 458262 158218 458346 158454
rect 458582 158218 458614 158454
rect 457994 158134 458614 158218
rect 457994 157898 458026 158134
rect 458262 157898 458346 158134
rect 458582 157898 458614 158134
rect 457994 131454 458614 157898
rect 457994 131218 458026 131454
rect 458262 131218 458346 131454
rect 458582 131218 458614 131454
rect 457994 131134 458614 131218
rect 457994 130898 458026 131134
rect 458262 130898 458346 131134
rect 458582 130898 458614 131134
rect 457994 104454 458614 130898
rect 457994 104218 458026 104454
rect 458262 104218 458346 104454
rect 458582 104218 458614 104454
rect 457994 104134 458614 104218
rect 457994 103898 458026 104134
rect 458262 103898 458346 104134
rect 458582 103898 458614 104134
rect 457994 77454 458614 103898
rect 457994 77218 458026 77454
rect 458262 77218 458346 77454
rect 458582 77218 458614 77454
rect 457994 77134 458614 77218
rect 457994 76898 458026 77134
rect 458262 76898 458346 77134
rect 458582 76898 458614 77134
rect 457994 69000 458614 76898
rect 461494 704838 462114 711590
rect 461494 704602 461526 704838
rect 461762 704602 461846 704838
rect 462082 704602 462114 704838
rect 461494 704518 462114 704602
rect 461494 704282 461526 704518
rect 461762 704282 461846 704518
rect 462082 704282 462114 704518
rect 461494 701829 462114 704282
rect 461494 701593 461526 701829
rect 461762 701593 461846 701829
rect 462082 701593 462114 701829
rect 461494 701509 462114 701593
rect 461494 701273 461526 701509
rect 461762 701273 461846 701509
rect 462082 701273 462114 701509
rect 461494 674829 462114 701273
rect 461494 674593 461526 674829
rect 461762 674593 461846 674829
rect 462082 674593 462114 674829
rect 461494 674509 462114 674593
rect 461494 674273 461526 674509
rect 461762 674273 461846 674509
rect 462082 674273 462114 674509
rect 461494 647829 462114 674273
rect 461494 647593 461526 647829
rect 461762 647593 461846 647829
rect 462082 647593 462114 647829
rect 461494 647509 462114 647593
rect 461494 647273 461526 647509
rect 461762 647273 461846 647509
rect 462082 647273 462114 647509
rect 461494 620829 462114 647273
rect 461494 620593 461526 620829
rect 461762 620593 461846 620829
rect 462082 620593 462114 620829
rect 461494 620509 462114 620593
rect 461494 620273 461526 620509
rect 461762 620273 461846 620509
rect 462082 620273 462114 620509
rect 461494 593829 462114 620273
rect 461494 593593 461526 593829
rect 461762 593593 461846 593829
rect 462082 593593 462114 593829
rect 461494 593509 462114 593593
rect 461494 593273 461526 593509
rect 461762 593273 461846 593509
rect 462082 593273 462114 593509
rect 461494 566829 462114 593273
rect 461494 566593 461526 566829
rect 461762 566593 461846 566829
rect 462082 566593 462114 566829
rect 461494 566509 462114 566593
rect 461494 566273 461526 566509
rect 461762 566273 461846 566509
rect 462082 566273 462114 566509
rect 461494 539829 462114 566273
rect 461494 539593 461526 539829
rect 461762 539593 461846 539829
rect 462082 539593 462114 539829
rect 461494 539509 462114 539593
rect 461494 539273 461526 539509
rect 461762 539273 461846 539509
rect 462082 539273 462114 539509
rect 461494 512829 462114 539273
rect 461494 512593 461526 512829
rect 461762 512593 461846 512829
rect 462082 512593 462114 512829
rect 461494 512509 462114 512593
rect 461494 512273 461526 512509
rect 461762 512273 461846 512509
rect 462082 512273 462114 512509
rect 461494 485829 462114 512273
rect 461494 485593 461526 485829
rect 461762 485593 461846 485829
rect 462082 485593 462114 485829
rect 461494 485509 462114 485593
rect 461494 485273 461526 485509
rect 461762 485273 461846 485509
rect 462082 485273 462114 485509
rect 461494 458829 462114 485273
rect 461494 458593 461526 458829
rect 461762 458593 461846 458829
rect 462082 458593 462114 458829
rect 461494 458509 462114 458593
rect 461494 458273 461526 458509
rect 461762 458273 461846 458509
rect 462082 458273 462114 458509
rect 461494 431829 462114 458273
rect 461494 431593 461526 431829
rect 461762 431593 461846 431829
rect 462082 431593 462114 431829
rect 461494 431509 462114 431593
rect 461494 431273 461526 431509
rect 461762 431273 461846 431509
rect 462082 431273 462114 431509
rect 461494 404829 462114 431273
rect 461494 404593 461526 404829
rect 461762 404593 461846 404829
rect 462082 404593 462114 404829
rect 461494 404509 462114 404593
rect 461494 404273 461526 404509
rect 461762 404273 461846 404509
rect 462082 404273 462114 404509
rect 461494 377829 462114 404273
rect 461494 377593 461526 377829
rect 461762 377593 461846 377829
rect 462082 377593 462114 377829
rect 461494 377509 462114 377593
rect 461494 377273 461526 377509
rect 461762 377273 461846 377509
rect 462082 377273 462114 377509
rect 461494 350829 462114 377273
rect 461494 350593 461526 350829
rect 461762 350593 461846 350829
rect 462082 350593 462114 350829
rect 461494 350509 462114 350593
rect 461494 350273 461526 350509
rect 461762 350273 461846 350509
rect 462082 350273 462114 350509
rect 461494 323829 462114 350273
rect 461494 323593 461526 323829
rect 461762 323593 461846 323829
rect 462082 323593 462114 323829
rect 461494 323509 462114 323593
rect 461494 323273 461526 323509
rect 461762 323273 461846 323509
rect 462082 323273 462114 323509
rect 461494 296829 462114 323273
rect 461494 296593 461526 296829
rect 461762 296593 461846 296829
rect 462082 296593 462114 296829
rect 461494 296509 462114 296593
rect 461494 296273 461526 296509
rect 461762 296273 461846 296509
rect 462082 296273 462114 296509
rect 461494 269829 462114 296273
rect 461494 269593 461526 269829
rect 461762 269593 461846 269829
rect 462082 269593 462114 269829
rect 461494 269509 462114 269593
rect 461494 269273 461526 269509
rect 461762 269273 461846 269509
rect 462082 269273 462114 269509
rect 461494 242829 462114 269273
rect 461494 242593 461526 242829
rect 461762 242593 461846 242829
rect 462082 242593 462114 242829
rect 461494 242509 462114 242593
rect 461494 242273 461526 242509
rect 461762 242273 461846 242509
rect 462082 242273 462114 242509
rect 461494 215829 462114 242273
rect 461494 215593 461526 215829
rect 461762 215593 461846 215829
rect 462082 215593 462114 215829
rect 461494 215509 462114 215593
rect 461494 215273 461526 215509
rect 461762 215273 461846 215509
rect 462082 215273 462114 215509
rect 461494 188829 462114 215273
rect 461494 188593 461526 188829
rect 461762 188593 461846 188829
rect 462082 188593 462114 188829
rect 461494 188509 462114 188593
rect 461494 188273 461526 188509
rect 461762 188273 461846 188509
rect 462082 188273 462114 188509
rect 461494 161829 462114 188273
rect 461494 161593 461526 161829
rect 461762 161593 461846 161829
rect 462082 161593 462114 161829
rect 461494 161509 462114 161593
rect 461494 161273 461526 161509
rect 461762 161273 461846 161509
rect 462082 161273 462114 161509
rect 461494 134829 462114 161273
rect 461494 134593 461526 134829
rect 461762 134593 461846 134829
rect 462082 134593 462114 134829
rect 461494 134509 462114 134593
rect 461494 134273 461526 134509
rect 461762 134273 461846 134509
rect 462082 134273 462114 134509
rect 461494 107829 462114 134273
rect 461494 107593 461526 107829
rect 461762 107593 461846 107829
rect 462082 107593 462114 107829
rect 461494 107509 462114 107593
rect 461494 107273 461526 107509
rect 461762 107273 461846 107509
rect 462082 107273 462114 107509
rect 461494 80829 462114 107273
rect 461494 80593 461526 80829
rect 461762 80593 461846 80829
rect 462082 80593 462114 80829
rect 461494 80509 462114 80593
rect 461494 80273 461526 80509
rect 461762 80273 461846 80509
rect 462082 80273 462114 80509
rect 461494 69000 462114 80273
rect 485994 705798 486614 711590
rect 485994 705562 486026 705798
rect 486262 705562 486346 705798
rect 486582 705562 486614 705798
rect 485994 705478 486614 705562
rect 485994 705242 486026 705478
rect 486262 705242 486346 705478
rect 486582 705242 486614 705478
rect 485994 698454 486614 705242
rect 485994 698218 486026 698454
rect 486262 698218 486346 698454
rect 486582 698218 486614 698454
rect 485994 698134 486614 698218
rect 485994 697898 486026 698134
rect 486262 697898 486346 698134
rect 486582 697898 486614 698134
rect 485994 671454 486614 697898
rect 485994 671218 486026 671454
rect 486262 671218 486346 671454
rect 486582 671218 486614 671454
rect 485994 671134 486614 671218
rect 485994 670898 486026 671134
rect 486262 670898 486346 671134
rect 486582 670898 486614 671134
rect 485994 644454 486614 670898
rect 485994 644218 486026 644454
rect 486262 644218 486346 644454
rect 486582 644218 486614 644454
rect 485994 644134 486614 644218
rect 485994 643898 486026 644134
rect 486262 643898 486346 644134
rect 486582 643898 486614 644134
rect 485994 617454 486614 643898
rect 485994 617218 486026 617454
rect 486262 617218 486346 617454
rect 486582 617218 486614 617454
rect 485994 617134 486614 617218
rect 485994 616898 486026 617134
rect 486262 616898 486346 617134
rect 486582 616898 486614 617134
rect 485994 590454 486614 616898
rect 485994 590218 486026 590454
rect 486262 590218 486346 590454
rect 486582 590218 486614 590454
rect 485994 590134 486614 590218
rect 485994 589898 486026 590134
rect 486262 589898 486346 590134
rect 486582 589898 486614 590134
rect 485994 563454 486614 589898
rect 485994 563218 486026 563454
rect 486262 563218 486346 563454
rect 486582 563218 486614 563454
rect 485994 563134 486614 563218
rect 485994 562898 486026 563134
rect 486262 562898 486346 563134
rect 486582 562898 486614 563134
rect 485994 536454 486614 562898
rect 485994 536218 486026 536454
rect 486262 536218 486346 536454
rect 486582 536218 486614 536454
rect 485994 536134 486614 536218
rect 485994 535898 486026 536134
rect 486262 535898 486346 536134
rect 486582 535898 486614 536134
rect 485994 509454 486614 535898
rect 485994 509218 486026 509454
rect 486262 509218 486346 509454
rect 486582 509218 486614 509454
rect 485994 509134 486614 509218
rect 485994 508898 486026 509134
rect 486262 508898 486346 509134
rect 486582 508898 486614 509134
rect 485994 482454 486614 508898
rect 485994 482218 486026 482454
rect 486262 482218 486346 482454
rect 486582 482218 486614 482454
rect 485994 482134 486614 482218
rect 485994 481898 486026 482134
rect 486262 481898 486346 482134
rect 486582 481898 486614 482134
rect 485994 455454 486614 481898
rect 485994 455218 486026 455454
rect 486262 455218 486346 455454
rect 486582 455218 486614 455454
rect 485994 455134 486614 455218
rect 485994 454898 486026 455134
rect 486262 454898 486346 455134
rect 486582 454898 486614 455134
rect 485994 428454 486614 454898
rect 485994 428218 486026 428454
rect 486262 428218 486346 428454
rect 486582 428218 486614 428454
rect 485994 428134 486614 428218
rect 485994 427898 486026 428134
rect 486262 427898 486346 428134
rect 486582 427898 486614 428134
rect 485994 401454 486614 427898
rect 485994 401218 486026 401454
rect 486262 401218 486346 401454
rect 486582 401218 486614 401454
rect 485994 401134 486614 401218
rect 485994 400898 486026 401134
rect 486262 400898 486346 401134
rect 486582 400898 486614 401134
rect 485994 374454 486614 400898
rect 485994 374218 486026 374454
rect 486262 374218 486346 374454
rect 486582 374218 486614 374454
rect 485994 374134 486614 374218
rect 485994 373898 486026 374134
rect 486262 373898 486346 374134
rect 486582 373898 486614 374134
rect 485994 347454 486614 373898
rect 485994 347218 486026 347454
rect 486262 347218 486346 347454
rect 486582 347218 486614 347454
rect 485994 347134 486614 347218
rect 485994 346898 486026 347134
rect 486262 346898 486346 347134
rect 486582 346898 486614 347134
rect 485994 320454 486614 346898
rect 485994 320218 486026 320454
rect 486262 320218 486346 320454
rect 486582 320218 486614 320454
rect 485994 320134 486614 320218
rect 485994 319898 486026 320134
rect 486262 319898 486346 320134
rect 486582 319898 486614 320134
rect 485994 293454 486614 319898
rect 485994 293218 486026 293454
rect 486262 293218 486346 293454
rect 486582 293218 486614 293454
rect 485994 293134 486614 293218
rect 485994 292898 486026 293134
rect 486262 292898 486346 293134
rect 486582 292898 486614 293134
rect 485994 266454 486614 292898
rect 485994 266218 486026 266454
rect 486262 266218 486346 266454
rect 486582 266218 486614 266454
rect 485994 266134 486614 266218
rect 485994 265898 486026 266134
rect 486262 265898 486346 266134
rect 486582 265898 486614 266134
rect 485994 239454 486614 265898
rect 485994 239218 486026 239454
rect 486262 239218 486346 239454
rect 486582 239218 486614 239454
rect 485994 239134 486614 239218
rect 485994 238898 486026 239134
rect 486262 238898 486346 239134
rect 486582 238898 486614 239134
rect 485994 212454 486614 238898
rect 485994 212218 486026 212454
rect 486262 212218 486346 212454
rect 486582 212218 486614 212454
rect 485994 212134 486614 212218
rect 485994 211898 486026 212134
rect 486262 211898 486346 212134
rect 486582 211898 486614 212134
rect 485994 185454 486614 211898
rect 485994 185218 486026 185454
rect 486262 185218 486346 185454
rect 486582 185218 486614 185454
rect 485994 185134 486614 185218
rect 485994 184898 486026 185134
rect 486262 184898 486346 185134
rect 486582 184898 486614 185134
rect 485994 158454 486614 184898
rect 485994 158218 486026 158454
rect 486262 158218 486346 158454
rect 486582 158218 486614 158454
rect 485994 158134 486614 158218
rect 485994 157898 486026 158134
rect 486262 157898 486346 158134
rect 486582 157898 486614 158134
rect 485994 131454 486614 157898
rect 485994 131218 486026 131454
rect 486262 131218 486346 131454
rect 486582 131218 486614 131454
rect 485994 131134 486614 131218
rect 485994 130898 486026 131134
rect 486262 130898 486346 131134
rect 486582 130898 486614 131134
rect 485994 104454 486614 130898
rect 485994 104218 486026 104454
rect 486262 104218 486346 104454
rect 486582 104218 486614 104454
rect 485994 104134 486614 104218
rect 485994 103898 486026 104134
rect 486262 103898 486346 104134
rect 486582 103898 486614 104134
rect 485994 77454 486614 103898
rect 485994 77218 486026 77454
rect 486262 77218 486346 77454
rect 486582 77218 486614 77454
rect 485994 77134 486614 77218
rect 485994 76898 486026 77134
rect 486262 76898 486346 77134
rect 486582 76898 486614 77134
rect 485994 69000 486614 76898
rect 489494 704838 490114 711590
rect 489494 704602 489526 704838
rect 489762 704602 489846 704838
rect 490082 704602 490114 704838
rect 489494 704518 490114 704602
rect 489494 704282 489526 704518
rect 489762 704282 489846 704518
rect 490082 704282 490114 704518
rect 489494 701829 490114 704282
rect 489494 701593 489526 701829
rect 489762 701593 489846 701829
rect 490082 701593 490114 701829
rect 489494 701509 490114 701593
rect 489494 701273 489526 701509
rect 489762 701273 489846 701509
rect 490082 701273 490114 701509
rect 489494 674829 490114 701273
rect 489494 674593 489526 674829
rect 489762 674593 489846 674829
rect 490082 674593 490114 674829
rect 489494 674509 490114 674593
rect 489494 674273 489526 674509
rect 489762 674273 489846 674509
rect 490082 674273 490114 674509
rect 489494 647829 490114 674273
rect 489494 647593 489526 647829
rect 489762 647593 489846 647829
rect 490082 647593 490114 647829
rect 489494 647509 490114 647593
rect 489494 647273 489526 647509
rect 489762 647273 489846 647509
rect 490082 647273 490114 647509
rect 489494 620829 490114 647273
rect 489494 620593 489526 620829
rect 489762 620593 489846 620829
rect 490082 620593 490114 620829
rect 489494 620509 490114 620593
rect 489494 620273 489526 620509
rect 489762 620273 489846 620509
rect 490082 620273 490114 620509
rect 489494 593829 490114 620273
rect 489494 593593 489526 593829
rect 489762 593593 489846 593829
rect 490082 593593 490114 593829
rect 489494 593509 490114 593593
rect 489494 593273 489526 593509
rect 489762 593273 489846 593509
rect 490082 593273 490114 593509
rect 489494 566829 490114 593273
rect 489494 566593 489526 566829
rect 489762 566593 489846 566829
rect 490082 566593 490114 566829
rect 489494 566509 490114 566593
rect 489494 566273 489526 566509
rect 489762 566273 489846 566509
rect 490082 566273 490114 566509
rect 489494 539829 490114 566273
rect 489494 539593 489526 539829
rect 489762 539593 489846 539829
rect 490082 539593 490114 539829
rect 489494 539509 490114 539593
rect 489494 539273 489526 539509
rect 489762 539273 489846 539509
rect 490082 539273 490114 539509
rect 489494 512829 490114 539273
rect 489494 512593 489526 512829
rect 489762 512593 489846 512829
rect 490082 512593 490114 512829
rect 489494 512509 490114 512593
rect 489494 512273 489526 512509
rect 489762 512273 489846 512509
rect 490082 512273 490114 512509
rect 489494 485829 490114 512273
rect 489494 485593 489526 485829
rect 489762 485593 489846 485829
rect 490082 485593 490114 485829
rect 489494 485509 490114 485593
rect 489494 485273 489526 485509
rect 489762 485273 489846 485509
rect 490082 485273 490114 485509
rect 489494 458829 490114 485273
rect 489494 458593 489526 458829
rect 489762 458593 489846 458829
rect 490082 458593 490114 458829
rect 489494 458509 490114 458593
rect 489494 458273 489526 458509
rect 489762 458273 489846 458509
rect 490082 458273 490114 458509
rect 489494 431829 490114 458273
rect 489494 431593 489526 431829
rect 489762 431593 489846 431829
rect 490082 431593 490114 431829
rect 489494 431509 490114 431593
rect 489494 431273 489526 431509
rect 489762 431273 489846 431509
rect 490082 431273 490114 431509
rect 489494 404829 490114 431273
rect 489494 404593 489526 404829
rect 489762 404593 489846 404829
rect 490082 404593 490114 404829
rect 489494 404509 490114 404593
rect 489494 404273 489526 404509
rect 489762 404273 489846 404509
rect 490082 404273 490114 404509
rect 489494 377829 490114 404273
rect 489494 377593 489526 377829
rect 489762 377593 489846 377829
rect 490082 377593 490114 377829
rect 489494 377509 490114 377593
rect 489494 377273 489526 377509
rect 489762 377273 489846 377509
rect 490082 377273 490114 377509
rect 489494 350829 490114 377273
rect 489494 350593 489526 350829
rect 489762 350593 489846 350829
rect 490082 350593 490114 350829
rect 489494 350509 490114 350593
rect 489494 350273 489526 350509
rect 489762 350273 489846 350509
rect 490082 350273 490114 350509
rect 489494 323829 490114 350273
rect 489494 323593 489526 323829
rect 489762 323593 489846 323829
rect 490082 323593 490114 323829
rect 489494 323509 490114 323593
rect 489494 323273 489526 323509
rect 489762 323273 489846 323509
rect 490082 323273 490114 323509
rect 489494 296829 490114 323273
rect 489494 296593 489526 296829
rect 489762 296593 489846 296829
rect 490082 296593 490114 296829
rect 489494 296509 490114 296593
rect 489494 296273 489526 296509
rect 489762 296273 489846 296509
rect 490082 296273 490114 296509
rect 489494 269829 490114 296273
rect 489494 269593 489526 269829
rect 489762 269593 489846 269829
rect 490082 269593 490114 269829
rect 489494 269509 490114 269593
rect 489494 269273 489526 269509
rect 489762 269273 489846 269509
rect 490082 269273 490114 269509
rect 489494 242829 490114 269273
rect 489494 242593 489526 242829
rect 489762 242593 489846 242829
rect 490082 242593 490114 242829
rect 489494 242509 490114 242593
rect 489494 242273 489526 242509
rect 489762 242273 489846 242509
rect 490082 242273 490114 242509
rect 489494 215829 490114 242273
rect 489494 215593 489526 215829
rect 489762 215593 489846 215829
rect 490082 215593 490114 215829
rect 489494 215509 490114 215593
rect 489494 215273 489526 215509
rect 489762 215273 489846 215509
rect 490082 215273 490114 215509
rect 489494 188829 490114 215273
rect 489494 188593 489526 188829
rect 489762 188593 489846 188829
rect 490082 188593 490114 188829
rect 489494 188509 490114 188593
rect 489494 188273 489526 188509
rect 489762 188273 489846 188509
rect 490082 188273 490114 188509
rect 489494 161829 490114 188273
rect 489494 161593 489526 161829
rect 489762 161593 489846 161829
rect 490082 161593 490114 161829
rect 489494 161509 490114 161593
rect 489494 161273 489526 161509
rect 489762 161273 489846 161509
rect 490082 161273 490114 161509
rect 489494 134829 490114 161273
rect 489494 134593 489526 134829
rect 489762 134593 489846 134829
rect 490082 134593 490114 134829
rect 489494 134509 490114 134593
rect 489494 134273 489526 134509
rect 489762 134273 489846 134509
rect 490082 134273 490114 134509
rect 489494 107829 490114 134273
rect 489494 107593 489526 107829
rect 489762 107593 489846 107829
rect 490082 107593 490114 107829
rect 489494 107509 490114 107593
rect 489494 107273 489526 107509
rect 489762 107273 489846 107509
rect 490082 107273 490114 107509
rect 489494 80829 490114 107273
rect 489494 80593 489526 80829
rect 489762 80593 489846 80829
rect 490082 80593 490114 80829
rect 489494 80509 490114 80593
rect 489494 80273 489526 80509
rect 489762 80273 489846 80509
rect 490082 80273 490114 80509
rect 489494 69000 490114 80273
rect 513994 705798 514614 711590
rect 513994 705562 514026 705798
rect 514262 705562 514346 705798
rect 514582 705562 514614 705798
rect 513994 705478 514614 705562
rect 513994 705242 514026 705478
rect 514262 705242 514346 705478
rect 514582 705242 514614 705478
rect 513994 698454 514614 705242
rect 513994 698218 514026 698454
rect 514262 698218 514346 698454
rect 514582 698218 514614 698454
rect 513994 698134 514614 698218
rect 513994 697898 514026 698134
rect 514262 697898 514346 698134
rect 514582 697898 514614 698134
rect 513994 671454 514614 697898
rect 513994 671218 514026 671454
rect 514262 671218 514346 671454
rect 514582 671218 514614 671454
rect 513994 671134 514614 671218
rect 513994 670898 514026 671134
rect 514262 670898 514346 671134
rect 514582 670898 514614 671134
rect 513994 644454 514614 670898
rect 513994 644218 514026 644454
rect 514262 644218 514346 644454
rect 514582 644218 514614 644454
rect 513994 644134 514614 644218
rect 513994 643898 514026 644134
rect 514262 643898 514346 644134
rect 514582 643898 514614 644134
rect 513994 617454 514614 643898
rect 513994 617218 514026 617454
rect 514262 617218 514346 617454
rect 514582 617218 514614 617454
rect 513994 617134 514614 617218
rect 513994 616898 514026 617134
rect 514262 616898 514346 617134
rect 514582 616898 514614 617134
rect 513994 590454 514614 616898
rect 513994 590218 514026 590454
rect 514262 590218 514346 590454
rect 514582 590218 514614 590454
rect 513994 590134 514614 590218
rect 513994 589898 514026 590134
rect 514262 589898 514346 590134
rect 514582 589898 514614 590134
rect 513994 563454 514614 589898
rect 513994 563218 514026 563454
rect 514262 563218 514346 563454
rect 514582 563218 514614 563454
rect 513994 563134 514614 563218
rect 513994 562898 514026 563134
rect 514262 562898 514346 563134
rect 514582 562898 514614 563134
rect 513994 536454 514614 562898
rect 513994 536218 514026 536454
rect 514262 536218 514346 536454
rect 514582 536218 514614 536454
rect 513994 536134 514614 536218
rect 513994 535898 514026 536134
rect 514262 535898 514346 536134
rect 514582 535898 514614 536134
rect 513994 509454 514614 535898
rect 513994 509218 514026 509454
rect 514262 509218 514346 509454
rect 514582 509218 514614 509454
rect 513994 509134 514614 509218
rect 513994 508898 514026 509134
rect 514262 508898 514346 509134
rect 514582 508898 514614 509134
rect 513994 482454 514614 508898
rect 513994 482218 514026 482454
rect 514262 482218 514346 482454
rect 514582 482218 514614 482454
rect 513994 482134 514614 482218
rect 513994 481898 514026 482134
rect 514262 481898 514346 482134
rect 514582 481898 514614 482134
rect 513994 455454 514614 481898
rect 513994 455218 514026 455454
rect 514262 455218 514346 455454
rect 514582 455218 514614 455454
rect 513994 455134 514614 455218
rect 513994 454898 514026 455134
rect 514262 454898 514346 455134
rect 514582 454898 514614 455134
rect 513994 428454 514614 454898
rect 513994 428218 514026 428454
rect 514262 428218 514346 428454
rect 514582 428218 514614 428454
rect 513994 428134 514614 428218
rect 513994 427898 514026 428134
rect 514262 427898 514346 428134
rect 514582 427898 514614 428134
rect 513994 401454 514614 427898
rect 513994 401218 514026 401454
rect 514262 401218 514346 401454
rect 514582 401218 514614 401454
rect 513994 401134 514614 401218
rect 513994 400898 514026 401134
rect 514262 400898 514346 401134
rect 514582 400898 514614 401134
rect 513994 374454 514614 400898
rect 513994 374218 514026 374454
rect 514262 374218 514346 374454
rect 514582 374218 514614 374454
rect 513994 374134 514614 374218
rect 513994 373898 514026 374134
rect 514262 373898 514346 374134
rect 514582 373898 514614 374134
rect 513994 347454 514614 373898
rect 513994 347218 514026 347454
rect 514262 347218 514346 347454
rect 514582 347218 514614 347454
rect 513994 347134 514614 347218
rect 513994 346898 514026 347134
rect 514262 346898 514346 347134
rect 514582 346898 514614 347134
rect 513994 320454 514614 346898
rect 513994 320218 514026 320454
rect 514262 320218 514346 320454
rect 514582 320218 514614 320454
rect 513994 320134 514614 320218
rect 513994 319898 514026 320134
rect 514262 319898 514346 320134
rect 514582 319898 514614 320134
rect 513994 293454 514614 319898
rect 513994 293218 514026 293454
rect 514262 293218 514346 293454
rect 514582 293218 514614 293454
rect 513994 293134 514614 293218
rect 513994 292898 514026 293134
rect 514262 292898 514346 293134
rect 514582 292898 514614 293134
rect 513994 266454 514614 292898
rect 513994 266218 514026 266454
rect 514262 266218 514346 266454
rect 514582 266218 514614 266454
rect 513994 266134 514614 266218
rect 513994 265898 514026 266134
rect 514262 265898 514346 266134
rect 514582 265898 514614 266134
rect 513994 239454 514614 265898
rect 513994 239218 514026 239454
rect 514262 239218 514346 239454
rect 514582 239218 514614 239454
rect 513994 239134 514614 239218
rect 513994 238898 514026 239134
rect 514262 238898 514346 239134
rect 514582 238898 514614 239134
rect 513994 212454 514614 238898
rect 513994 212218 514026 212454
rect 514262 212218 514346 212454
rect 514582 212218 514614 212454
rect 513994 212134 514614 212218
rect 513994 211898 514026 212134
rect 514262 211898 514346 212134
rect 514582 211898 514614 212134
rect 513994 185454 514614 211898
rect 513994 185218 514026 185454
rect 514262 185218 514346 185454
rect 514582 185218 514614 185454
rect 513994 185134 514614 185218
rect 513994 184898 514026 185134
rect 514262 184898 514346 185134
rect 514582 184898 514614 185134
rect 513994 158454 514614 184898
rect 513994 158218 514026 158454
rect 514262 158218 514346 158454
rect 514582 158218 514614 158454
rect 513994 158134 514614 158218
rect 513994 157898 514026 158134
rect 514262 157898 514346 158134
rect 514582 157898 514614 158134
rect 513994 131454 514614 157898
rect 513994 131218 514026 131454
rect 514262 131218 514346 131454
rect 514582 131218 514614 131454
rect 513994 131134 514614 131218
rect 513994 130898 514026 131134
rect 514262 130898 514346 131134
rect 514582 130898 514614 131134
rect 513994 104454 514614 130898
rect 513994 104218 514026 104454
rect 514262 104218 514346 104454
rect 514582 104218 514614 104454
rect 513994 104134 514614 104218
rect 513994 103898 514026 104134
rect 514262 103898 514346 104134
rect 514582 103898 514614 104134
rect 513994 77454 514614 103898
rect 513994 77218 514026 77454
rect 514262 77218 514346 77454
rect 514582 77218 514614 77454
rect 513994 77134 514614 77218
rect 513994 76898 514026 77134
rect 514262 76898 514346 77134
rect 514582 76898 514614 77134
rect 513994 69000 514614 76898
rect 517494 704838 518114 711590
rect 517494 704602 517526 704838
rect 517762 704602 517846 704838
rect 518082 704602 518114 704838
rect 517494 704518 518114 704602
rect 517494 704282 517526 704518
rect 517762 704282 517846 704518
rect 518082 704282 518114 704518
rect 517494 701829 518114 704282
rect 517494 701593 517526 701829
rect 517762 701593 517846 701829
rect 518082 701593 518114 701829
rect 517494 701509 518114 701593
rect 517494 701273 517526 701509
rect 517762 701273 517846 701509
rect 518082 701273 518114 701509
rect 517494 674829 518114 701273
rect 541994 705798 542614 711590
rect 541994 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 542614 705798
rect 541994 705478 542614 705562
rect 541994 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 542614 705478
rect 527403 699820 527469 699821
rect 527403 699756 527404 699820
rect 527468 699756 527469 699820
rect 527403 699755 527469 699756
rect 517494 674593 517526 674829
rect 517762 674593 517846 674829
rect 518082 674593 518114 674829
rect 517494 674509 518114 674593
rect 517494 674273 517526 674509
rect 517762 674273 517846 674509
rect 518082 674273 518114 674509
rect 517494 647829 518114 674273
rect 517494 647593 517526 647829
rect 517762 647593 517846 647829
rect 518082 647593 518114 647829
rect 517494 647509 518114 647593
rect 517494 647273 517526 647509
rect 517762 647273 517846 647509
rect 518082 647273 518114 647509
rect 517494 620829 518114 647273
rect 517494 620593 517526 620829
rect 517762 620593 517846 620829
rect 518082 620593 518114 620829
rect 517494 620509 518114 620593
rect 517494 620273 517526 620509
rect 517762 620273 517846 620509
rect 518082 620273 518114 620509
rect 517494 593829 518114 620273
rect 517494 593593 517526 593829
rect 517762 593593 517846 593829
rect 518082 593593 518114 593829
rect 517494 593509 518114 593593
rect 517494 593273 517526 593509
rect 517762 593273 517846 593509
rect 518082 593273 518114 593509
rect 517494 566829 518114 593273
rect 517494 566593 517526 566829
rect 517762 566593 517846 566829
rect 518082 566593 518114 566829
rect 517494 566509 518114 566593
rect 517494 566273 517526 566509
rect 517762 566273 517846 566509
rect 518082 566273 518114 566509
rect 517494 539829 518114 566273
rect 517494 539593 517526 539829
rect 517762 539593 517846 539829
rect 518082 539593 518114 539829
rect 517494 539509 518114 539593
rect 517494 539273 517526 539509
rect 517762 539273 517846 539509
rect 518082 539273 518114 539509
rect 517494 512829 518114 539273
rect 517494 512593 517526 512829
rect 517762 512593 517846 512829
rect 518082 512593 518114 512829
rect 517494 512509 518114 512593
rect 517494 512273 517526 512509
rect 517762 512273 517846 512509
rect 518082 512273 518114 512509
rect 517494 485829 518114 512273
rect 517494 485593 517526 485829
rect 517762 485593 517846 485829
rect 518082 485593 518114 485829
rect 517494 485509 518114 485593
rect 517494 485273 517526 485509
rect 517762 485273 517846 485509
rect 518082 485273 518114 485509
rect 517494 458829 518114 485273
rect 517494 458593 517526 458829
rect 517762 458593 517846 458829
rect 518082 458593 518114 458829
rect 517494 458509 518114 458593
rect 517494 458273 517526 458509
rect 517762 458273 517846 458509
rect 518082 458273 518114 458509
rect 517494 431829 518114 458273
rect 517494 431593 517526 431829
rect 517762 431593 517846 431829
rect 518082 431593 518114 431829
rect 517494 431509 518114 431593
rect 517494 431273 517526 431509
rect 517762 431273 517846 431509
rect 518082 431273 518114 431509
rect 517494 404829 518114 431273
rect 517494 404593 517526 404829
rect 517762 404593 517846 404829
rect 518082 404593 518114 404829
rect 517494 404509 518114 404593
rect 517494 404273 517526 404509
rect 517762 404273 517846 404509
rect 518082 404273 518114 404509
rect 517494 377829 518114 404273
rect 517494 377593 517526 377829
rect 517762 377593 517846 377829
rect 518082 377593 518114 377829
rect 517494 377509 518114 377593
rect 517494 377273 517526 377509
rect 517762 377273 517846 377509
rect 518082 377273 518114 377509
rect 517494 350829 518114 377273
rect 517494 350593 517526 350829
rect 517762 350593 517846 350829
rect 518082 350593 518114 350829
rect 517494 350509 518114 350593
rect 517494 350273 517526 350509
rect 517762 350273 517846 350509
rect 518082 350273 518114 350509
rect 517494 323829 518114 350273
rect 517494 323593 517526 323829
rect 517762 323593 517846 323829
rect 518082 323593 518114 323829
rect 517494 323509 518114 323593
rect 517494 323273 517526 323509
rect 517762 323273 517846 323509
rect 518082 323273 518114 323509
rect 517494 296829 518114 323273
rect 517494 296593 517526 296829
rect 517762 296593 517846 296829
rect 518082 296593 518114 296829
rect 517494 296509 518114 296593
rect 517494 296273 517526 296509
rect 517762 296273 517846 296509
rect 518082 296273 518114 296509
rect 517494 269829 518114 296273
rect 517494 269593 517526 269829
rect 517762 269593 517846 269829
rect 518082 269593 518114 269829
rect 517494 269509 518114 269593
rect 517494 269273 517526 269509
rect 517762 269273 517846 269509
rect 518082 269273 518114 269509
rect 517494 242829 518114 269273
rect 517494 242593 517526 242829
rect 517762 242593 517846 242829
rect 518082 242593 518114 242829
rect 517494 242509 518114 242593
rect 517494 242273 517526 242509
rect 517762 242273 517846 242509
rect 518082 242273 518114 242509
rect 517494 215829 518114 242273
rect 517494 215593 517526 215829
rect 517762 215593 517846 215829
rect 518082 215593 518114 215829
rect 517494 215509 518114 215593
rect 517494 215273 517526 215509
rect 517762 215273 517846 215509
rect 518082 215273 518114 215509
rect 517494 188829 518114 215273
rect 517494 188593 517526 188829
rect 517762 188593 517846 188829
rect 518082 188593 518114 188829
rect 517494 188509 518114 188593
rect 517494 188273 517526 188509
rect 517762 188273 517846 188509
rect 518082 188273 518114 188509
rect 517494 161829 518114 188273
rect 517494 161593 517526 161829
rect 517762 161593 517846 161829
rect 518082 161593 518114 161829
rect 517494 161509 518114 161593
rect 517494 161273 517526 161509
rect 517762 161273 517846 161509
rect 518082 161273 518114 161509
rect 517494 134829 518114 161273
rect 517494 134593 517526 134829
rect 517762 134593 517846 134829
rect 518082 134593 518114 134829
rect 517494 134509 518114 134593
rect 517494 134273 517526 134509
rect 517762 134273 517846 134509
rect 518082 134273 518114 134509
rect 517494 107829 518114 134273
rect 517494 107593 517526 107829
rect 517762 107593 517846 107829
rect 518082 107593 518114 107829
rect 517494 107509 518114 107593
rect 517494 107273 517526 107509
rect 517762 107273 517846 107509
rect 518082 107273 518114 107509
rect 517494 80829 518114 107273
rect 517494 80593 517526 80829
rect 517762 80593 517846 80829
rect 518082 80593 518114 80829
rect 517494 80509 518114 80593
rect 517494 80273 517526 80509
rect 517762 80273 517846 80509
rect 518082 80273 518114 80509
rect 517494 69000 518114 80273
rect 432814 53829 433134 53861
rect 432814 53593 432856 53829
rect 433092 53593 433134 53829
rect 432814 53509 433134 53593
rect 432814 53273 432856 53509
rect 433092 53273 433134 53509
rect 432814 53241 433134 53273
rect 436762 53829 437082 53861
rect 436762 53593 436804 53829
rect 437040 53593 437082 53829
rect 436762 53509 437082 53593
rect 436762 53273 436804 53509
rect 437040 53273 437082 53509
rect 436762 53241 437082 53273
rect 445218 53829 445538 53861
rect 445218 53593 445260 53829
rect 445496 53593 445538 53829
rect 445218 53509 445538 53593
rect 445218 53273 445260 53509
rect 445496 53273 445538 53509
rect 445218 53241 445538 53273
rect 446166 53829 446486 53861
rect 446166 53593 446208 53829
rect 446444 53593 446486 53829
rect 446166 53509 446486 53593
rect 446166 53273 446208 53509
rect 446444 53273 446486 53509
rect 446166 53241 446486 53273
rect 447114 53829 447434 53861
rect 447114 53593 447156 53829
rect 447392 53593 447434 53829
rect 447114 53509 447434 53593
rect 447114 53273 447156 53509
rect 447392 53273 447434 53509
rect 447114 53241 447434 53273
rect 448062 53829 448382 53861
rect 448062 53593 448104 53829
rect 448340 53593 448382 53829
rect 448062 53509 448382 53593
rect 448062 53273 448104 53509
rect 448340 53273 448382 53509
rect 448062 53241 448382 53273
rect 453918 53829 454238 53861
rect 453918 53593 453960 53829
rect 454196 53593 454238 53829
rect 453918 53509 454238 53593
rect 453918 53273 453960 53509
rect 454196 53273 454238 53509
rect 453918 53241 454238 53273
rect 457866 53829 458186 53861
rect 457866 53593 457908 53829
rect 458144 53593 458186 53829
rect 457866 53509 458186 53593
rect 457866 53273 457908 53509
rect 458144 53273 458186 53509
rect 457866 53241 458186 53273
rect 461814 53829 462134 53861
rect 461814 53593 461856 53829
rect 462092 53593 462134 53829
rect 461814 53509 462134 53593
rect 461814 53273 461856 53509
rect 462092 53273 462134 53509
rect 461814 53241 462134 53273
rect 465762 53829 466082 53861
rect 465762 53593 465804 53829
rect 466040 53593 466082 53829
rect 465762 53509 466082 53593
rect 465762 53273 465804 53509
rect 466040 53273 466082 53509
rect 465762 53241 466082 53273
rect 474218 53829 474538 53861
rect 474218 53593 474260 53829
rect 474496 53593 474538 53829
rect 474218 53509 474538 53593
rect 474218 53273 474260 53509
rect 474496 53273 474538 53509
rect 474218 53241 474538 53273
rect 475166 53829 475486 53861
rect 475166 53593 475208 53829
rect 475444 53593 475486 53829
rect 475166 53509 475486 53593
rect 475166 53273 475208 53509
rect 475444 53273 475486 53509
rect 475166 53241 475486 53273
rect 476114 53829 476434 53861
rect 476114 53593 476156 53829
rect 476392 53593 476434 53829
rect 476114 53509 476434 53593
rect 476114 53273 476156 53509
rect 476392 53273 476434 53509
rect 476114 53241 476434 53273
rect 477062 53829 477382 53861
rect 477062 53593 477104 53829
rect 477340 53593 477382 53829
rect 477062 53509 477382 53593
rect 477062 53273 477104 53509
rect 477340 53273 477382 53509
rect 477062 53241 477382 53273
rect 482918 53829 483238 53861
rect 482918 53593 482960 53829
rect 483196 53593 483238 53829
rect 482918 53509 483238 53593
rect 482918 53273 482960 53509
rect 483196 53273 483238 53509
rect 482918 53241 483238 53273
rect 486866 53829 487186 53861
rect 486866 53593 486908 53829
rect 487144 53593 487186 53829
rect 486866 53509 487186 53593
rect 486866 53273 486908 53509
rect 487144 53273 487186 53509
rect 486866 53241 487186 53273
rect 490814 53829 491134 53861
rect 490814 53593 490856 53829
rect 491092 53593 491134 53829
rect 490814 53509 491134 53593
rect 490814 53273 490856 53509
rect 491092 53273 491134 53509
rect 490814 53241 491134 53273
rect 494762 53829 495082 53861
rect 494762 53593 494804 53829
rect 495040 53593 495082 53829
rect 494762 53509 495082 53593
rect 494762 53273 494804 53509
rect 495040 53273 495082 53509
rect 494762 53241 495082 53273
rect 503218 53829 503538 53861
rect 503218 53593 503260 53829
rect 503496 53593 503538 53829
rect 503218 53509 503538 53593
rect 503218 53273 503260 53509
rect 503496 53273 503538 53509
rect 503218 53241 503538 53273
rect 504166 53829 504486 53861
rect 504166 53593 504208 53829
rect 504444 53593 504486 53829
rect 504166 53509 504486 53593
rect 504166 53273 504208 53509
rect 504444 53273 504486 53509
rect 504166 53241 504486 53273
rect 505114 53829 505434 53861
rect 505114 53593 505156 53829
rect 505392 53593 505434 53829
rect 505114 53509 505434 53593
rect 505114 53273 505156 53509
rect 505392 53273 505434 53509
rect 505114 53241 505434 53273
rect 506062 53829 506382 53861
rect 506062 53593 506104 53829
rect 506340 53593 506382 53829
rect 506062 53509 506382 53593
rect 506062 53273 506104 53509
rect 506340 53273 506382 53509
rect 506062 53241 506382 53273
rect 511918 53829 512238 53861
rect 511918 53593 511960 53829
rect 512196 53593 512238 53829
rect 511918 53509 512238 53593
rect 511918 53273 511960 53509
rect 512196 53273 512238 53509
rect 511918 53241 512238 53273
rect 515866 53829 516186 53861
rect 515866 53593 515908 53829
rect 516144 53593 516186 53829
rect 515866 53509 516186 53593
rect 515866 53273 515908 53509
rect 516144 53273 516186 53509
rect 515866 53241 516186 53273
rect 519814 53829 520134 53861
rect 519814 53593 519856 53829
rect 520092 53593 520134 53829
rect 519814 53509 520134 53593
rect 519814 53273 519856 53509
rect 520092 53273 520134 53509
rect 519814 53241 520134 53273
rect 523762 53829 524082 53861
rect 523762 53593 523804 53829
rect 524040 53593 524082 53829
rect 523762 53509 524082 53593
rect 523762 53273 523804 53509
rect 524040 53273 524082 53509
rect 523762 53241 524082 53273
rect 430840 50454 431160 50486
rect 430840 50218 430882 50454
rect 431118 50218 431160 50454
rect 430840 50134 431160 50218
rect 430840 49898 430882 50134
rect 431118 49898 431160 50134
rect 430840 49866 431160 49898
rect 434788 50454 435108 50486
rect 434788 50218 434830 50454
rect 435066 50218 435108 50454
rect 434788 50134 435108 50218
rect 434788 49898 434830 50134
rect 435066 49898 435108 50134
rect 434788 49866 435108 49898
rect 445692 50454 446012 50486
rect 445692 50218 445734 50454
rect 445970 50218 446012 50454
rect 445692 50134 446012 50218
rect 445692 49898 445734 50134
rect 445970 49898 446012 50134
rect 445692 49866 446012 49898
rect 446640 50454 446960 50486
rect 446640 50218 446682 50454
rect 446918 50218 446960 50454
rect 446640 50134 446960 50218
rect 446640 49898 446682 50134
rect 446918 49898 446960 50134
rect 446640 49866 446960 49898
rect 447588 50454 447908 50486
rect 447588 50218 447630 50454
rect 447866 50218 447908 50454
rect 447588 50134 447908 50218
rect 447588 49898 447630 50134
rect 447866 49898 447908 50134
rect 447588 49866 447908 49898
rect 455892 50454 456212 50486
rect 455892 50218 455934 50454
rect 456170 50218 456212 50454
rect 455892 50134 456212 50218
rect 455892 49898 455934 50134
rect 456170 49898 456212 50134
rect 455892 49866 456212 49898
rect 459840 50454 460160 50486
rect 459840 50218 459882 50454
rect 460118 50218 460160 50454
rect 459840 50134 460160 50218
rect 459840 49898 459882 50134
rect 460118 49898 460160 50134
rect 459840 49866 460160 49898
rect 463788 50454 464108 50486
rect 463788 50218 463830 50454
rect 464066 50218 464108 50454
rect 463788 50134 464108 50218
rect 463788 49898 463830 50134
rect 464066 49898 464108 50134
rect 463788 49866 464108 49898
rect 474692 50454 475012 50486
rect 474692 50218 474734 50454
rect 474970 50218 475012 50454
rect 474692 50134 475012 50218
rect 474692 49898 474734 50134
rect 474970 49898 475012 50134
rect 474692 49866 475012 49898
rect 475640 50454 475960 50486
rect 475640 50218 475682 50454
rect 475918 50218 475960 50454
rect 475640 50134 475960 50218
rect 475640 49898 475682 50134
rect 475918 49898 475960 50134
rect 475640 49866 475960 49898
rect 476588 50454 476908 50486
rect 476588 50218 476630 50454
rect 476866 50218 476908 50454
rect 476588 50134 476908 50218
rect 476588 49898 476630 50134
rect 476866 49898 476908 50134
rect 476588 49866 476908 49898
rect 484892 50454 485212 50486
rect 484892 50218 484934 50454
rect 485170 50218 485212 50454
rect 484892 50134 485212 50218
rect 484892 49898 484934 50134
rect 485170 49898 485212 50134
rect 484892 49866 485212 49898
rect 488840 50454 489160 50486
rect 488840 50218 488882 50454
rect 489118 50218 489160 50454
rect 488840 50134 489160 50218
rect 488840 49898 488882 50134
rect 489118 49898 489160 50134
rect 488840 49866 489160 49898
rect 492788 50454 493108 50486
rect 492788 50218 492830 50454
rect 493066 50218 493108 50454
rect 492788 50134 493108 50218
rect 492788 49898 492830 50134
rect 493066 49898 493108 50134
rect 492788 49866 493108 49898
rect 503692 50454 504012 50486
rect 503692 50218 503734 50454
rect 503970 50218 504012 50454
rect 503692 50134 504012 50218
rect 503692 49898 503734 50134
rect 503970 49898 504012 50134
rect 503692 49866 504012 49898
rect 504640 50454 504960 50486
rect 504640 50218 504682 50454
rect 504918 50218 504960 50454
rect 504640 50134 504960 50218
rect 504640 49898 504682 50134
rect 504918 49898 504960 50134
rect 504640 49866 504960 49898
rect 505588 50454 505908 50486
rect 505588 50218 505630 50454
rect 505866 50218 505908 50454
rect 505588 50134 505908 50218
rect 505588 49898 505630 50134
rect 505866 49898 505908 50134
rect 505588 49866 505908 49898
rect 513892 50454 514212 50486
rect 513892 50218 513934 50454
rect 514170 50218 514212 50454
rect 513892 50134 514212 50218
rect 513892 49898 513934 50134
rect 514170 49898 514212 50134
rect 513892 49866 514212 49898
rect 517840 50454 518160 50486
rect 517840 50218 517882 50454
rect 518118 50218 518160 50454
rect 517840 50134 518160 50218
rect 517840 49898 517882 50134
rect 518118 49898 518160 50134
rect 517840 49866 518160 49898
rect 521788 50454 522108 50486
rect 521788 50218 521830 50454
rect 522066 50218 522108 50454
rect 521788 50134 522108 50218
rect 521788 49898 521830 50134
rect 522066 49898 522108 50134
rect 521788 49866 522108 49898
rect 432118 26829 432438 26861
rect 432118 26593 432160 26829
rect 432396 26593 432438 26829
rect 432118 26509 432438 26593
rect 432118 26273 432160 26509
rect 432396 26273 432438 26509
rect 432118 26241 432438 26273
rect 436066 26829 436386 26861
rect 436066 26593 436108 26829
rect 436344 26593 436386 26829
rect 436066 26509 436386 26593
rect 436066 26273 436108 26509
rect 436344 26273 436386 26509
rect 436066 26241 436386 26273
rect 440014 26829 440334 26861
rect 440014 26593 440056 26829
rect 440292 26593 440334 26829
rect 440014 26509 440334 26593
rect 440014 26273 440056 26509
rect 440292 26273 440334 26509
rect 440014 26241 440334 26273
rect 443962 26829 444282 26861
rect 443962 26593 444004 26829
rect 444240 26593 444282 26829
rect 443962 26509 444282 26593
rect 443962 26273 444004 26509
rect 444240 26273 444282 26509
rect 443962 26241 444282 26273
rect 452418 26829 452738 26861
rect 452418 26593 452460 26829
rect 452696 26593 452738 26829
rect 452418 26509 452738 26593
rect 452418 26273 452460 26509
rect 452696 26273 452738 26509
rect 452418 26241 452738 26273
rect 453366 26829 453686 26861
rect 453366 26593 453408 26829
rect 453644 26593 453686 26829
rect 453366 26509 453686 26593
rect 453366 26273 453408 26509
rect 453644 26273 453686 26509
rect 453366 26241 453686 26273
rect 454314 26829 454634 26861
rect 454314 26593 454356 26829
rect 454592 26593 454634 26829
rect 454314 26509 454634 26593
rect 454314 26273 454356 26509
rect 454592 26273 454634 26509
rect 454314 26241 454634 26273
rect 455262 26829 455582 26861
rect 455262 26593 455304 26829
rect 455540 26593 455582 26829
rect 455262 26509 455582 26593
rect 455262 26273 455304 26509
rect 455540 26273 455582 26509
rect 455262 26241 455582 26273
rect 461118 26829 461438 26861
rect 461118 26593 461160 26829
rect 461396 26593 461438 26829
rect 461118 26509 461438 26593
rect 461118 26273 461160 26509
rect 461396 26273 461438 26509
rect 461118 26241 461438 26273
rect 465066 26829 465386 26861
rect 465066 26593 465108 26829
rect 465344 26593 465386 26829
rect 465066 26509 465386 26593
rect 465066 26273 465108 26509
rect 465344 26273 465386 26509
rect 465066 26241 465386 26273
rect 469014 26829 469334 26861
rect 469014 26593 469056 26829
rect 469292 26593 469334 26829
rect 469014 26509 469334 26593
rect 469014 26273 469056 26509
rect 469292 26273 469334 26509
rect 469014 26241 469334 26273
rect 472962 26829 473282 26861
rect 472962 26593 473004 26829
rect 473240 26593 473282 26829
rect 472962 26509 473282 26593
rect 472962 26273 473004 26509
rect 473240 26273 473282 26509
rect 472962 26241 473282 26273
rect 481418 26829 481738 26861
rect 481418 26593 481460 26829
rect 481696 26593 481738 26829
rect 481418 26509 481738 26593
rect 481418 26273 481460 26509
rect 481696 26273 481738 26509
rect 481418 26241 481738 26273
rect 482366 26829 482686 26861
rect 482366 26593 482408 26829
rect 482644 26593 482686 26829
rect 482366 26509 482686 26593
rect 482366 26273 482408 26509
rect 482644 26273 482686 26509
rect 482366 26241 482686 26273
rect 483314 26829 483634 26861
rect 483314 26593 483356 26829
rect 483592 26593 483634 26829
rect 483314 26509 483634 26593
rect 483314 26273 483356 26509
rect 483592 26273 483634 26509
rect 483314 26241 483634 26273
rect 484262 26829 484582 26861
rect 484262 26593 484304 26829
rect 484540 26593 484582 26829
rect 484262 26509 484582 26593
rect 484262 26273 484304 26509
rect 484540 26273 484582 26509
rect 484262 26241 484582 26273
rect 490118 26829 490438 26861
rect 490118 26593 490160 26829
rect 490396 26593 490438 26829
rect 490118 26509 490438 26593
rect 490118 26273 490160 26509
rect 490396 26273 490438 26509
rect 490118 26241 490438 26273
rect 494066 26829 494386 26861
rect 494066 26593 494108 26829
rect 494344 26593 494386 26829
rect 494066 26509 494386 26593
rect 494066 26273 494108 26509
rect 494344 26273 494386 26509
rect 494066 26241 494386 26273
rect 498014 26829 498334 26861
rect 498014 26593 498056 26829
rect 498292 26593 498334 26829
rect 498014 26509 498334 26593
rect 498014 26273 498056 26509
rect 498292 26273 498334 26509
rect 498014 26241 498334 26273
rect 501962 26829 502282 26861
rect 501962 26593 502004 26829
rect 502240 26593 502282 26829
rect 501962 26509 502282 26593
rect 501962 26273 502004 26509
rect 502240 26273 502282 26509
rect 501962 26241 502282 26273
rect 510418 26829 510738 26861
rect 510418 26593 510460 26829
rect 510696 26593 510738 26829
rect 510418 26509 510738 26593
rect 510418 26273 510460 26509
rect 510696 26273 510738 26509
rect 510418 26241 510738 26273
rect 511366 26829 511686 26861
rect 511366 26593 511408 26829
rect 511644 26593 511686 26829
rect 511366 26509 511686 26593
rect 511366 26273 511408 26509
rect 511644 26273 511686 26509
rect 511366 26241 511686 26273
rect 512314 26829 512634 26861
rect 512314 26593 512356 26829
rect 512592 26593 512634 26829
rect 512314 26509 512634 26593
rect 512314 26273 512356 26509
rect 512592 26273 512634 26509
rect 512314 26241 512634 26273
rect 513262 26829 513582 26861
rect 513262 26593 513304 26829
rect 513540 26593 513582 26829
rect 513262 26509 513582 26593
rect 513262 26273 513304 26509
rect 513540 26273 513582 26509
rect 513262 26241 513582 26273
rect 519118 26829 519438 26861
rect 519118 26593 519160 26829
rect 519396 26593 519438 26829
rect 519118 26509 519438 26593
rect 519118 26273 519160 26509
rect 519396 26273 519438 26509
rect 519118 26241 519438 26273
rect 523066 26829 523386 26861
rect 523066 26593 523108 26829
rect 523344 26593 523386 26829
rect 523066 26509 523386 26593
rect 523066 26273 523108 26509
rect 523344 26273 523386 26509
rect 523066 26241 523386 26273
rect 527014 26829 527334 26861
rect 527014 26593 527056 26829
rect 527292 26593 527334 26829
rect 527014 26509 527334 26593
rect 527014 26273 527056 26509
rect 527292 26273 527334 26509
rect 527014 26241 527334 26273
rect 434092 23454 434412 23486
rect 434092 23218 434134 23454
rect 434370 23218 434412 23454
rect 434092 23134 434412 23218
rect 434092 22898 434134 23134
rect 434370 22898 434412 23134
rect 434092 22866 434412 22898
rect 438040 23454 438360 23486
rect 438040 23218 438082 23454
rect 438318 23218 438360 23454
rect 438040 23134 438360 23218
rect 438040 22898 438082 23134
rect 438318 22898 438360 23134
rect 438040 22866 438360 22898
rect 441988 23454 442308 23486
rect 441988 23218 442030 23454
rect 442266 23218 442308 23454
rect 441988 23134 442308 23218
rect 441988 22898 442030 23134
rect 442266 22898 442308 23134
rect 441988 22866 442308 22898
rect 452892 23454 453212 23486
rect 452892 23218 452934 23454
rect 453170 23218 453212 23454
rect 452892 23134 453212 23218
rect 452892 22898 452934 23134
rect 453170 22898 453212 23134
rect 452892 22866 453212 22898
rect 453840 23454 454160 23486
rect 453840 23218 453882 23454
rect 454118 23218 454160 23454
rect 453840 23134 454160 23218
rect 453840 22898 453882 23134
rect 454118 22898 454160 23134
rect 453840 22866 454160 22898
rect 454788 23454 455108 23486
rect 454788 23218 454830 23454
rect 455066 23218 455108 23454
rect 454788 23134 455108 23218
rect 454788 22898 454830 23134
rect 455066 22898 455108 23134
rect 454788 22866 455108 22898
rect 463092 23454 463412 23486
rect 463092 23218 463134 23454
rect 463370 23218 463412 23454
rect 463092 23134 463412 23218
rect 463092 22898 463134 23134
rect 463370 22898 463412 23134
rect 463092 22866 463412 22898
rect 467040 23454 467360 23486
rect 467040 23218 467082 23454
rect 467318 23218 467360 23454
rect 467040 23134 467360 23218
rect 467040 22898 467082 23134
rect 467318 22898 467360 23134
rect 467040 22866 467360 22898
rect 470988 23454 471308 23486
rect 470988 23218 471030 23454
rect 471266 23218 471308 23454
rect 470988 23134 471308 23218
rect 470988 22898 471030 23134
rect 471266 22898 471308 23134
rect 470988 22866 471308 22898
rect 481892 23454 482212 23486
rect 481892 23218 481934 23454
rect 482170 23218 482212 23454
rect 481892 23134 482212 23218
rect 481892 22898 481934 23134
rect 482170 22898 482212 23134
rect 481892 22866 482212 22898
rect 482840 23454 483160 23486
rect 482840 23218 482882 23454
rect 483118 23218 483160 23454
rect 482840 23134 483160 23218
rect 482840 22898 482882 23134
rect 483118 22898 483160 23134
rect 482840 22866 483160 22898
rect 483788 23454 484108 23486
rect 483788 23218 483830 23454
rect 484066 23218 484108 23454
rect 483788 23134 484108 23218
rect 483788 22898 483830 23134
rect 484066 22898 484108 23134
rect 483788 22866 484108 22898
rect 492092 23454 492412 23486
rect 492092 23218 492134 23454
rect 492370 23218 492412 23454
rect 492092 23134 492412 23218
rect 492092 22898 492134 23134
rect 492370 22898 492412 23134
rect 492092 22866 492412 22898
rect 496040 23454 496360 23486
rect 496040 23218 496082 23454
rect 496318 23218 496360 23454
rect 496040 23134 496360 23218
rect 496040 22898 496082 23134
rect 496318 22898 496360 23134
rect 496040 22866 496360 22898
rect 499988 23454 500308 23486
rect 499988 23218 500030 23454
rect 500266 23218 500308 23454
rect 499988 23134 500308 23218
rect 499988 22898 500030 23134
rect 500266 22898 500308 23134
rect 499988 22866 500308 22898
rect 510892 23454 511212 23486
rect 510892 23218 510934 23454
rect 511170 23218 511212 23454
rect 510892 23134 511212 23218
rect 510892 22898 510934 23134
rect 511170 22898 511212 23134
rect 510892 22866 511212 22898
rect 511840 23454 512160 23486
rect 511840 23218 511882 23454
rect 512118 23218 512160 23454
rect 511840 23134 512160 23218
rect 511840 22898 511882 23134
rect 512118 22898 512160 23134
rect 511840 22866 512160 22898
rect 512788 23454 513108 23486
rect 512788 23218 512830 23454
rect 513066 23218 513108 23454
rect 512788 23134 513108 23218
rect 512788 22898 512830 23134
rect 513066 22898 513108 23134
rect 512788 22866 513108 22898
rect 521092 23454 521412 23486
rect 521092 23218 521134 23454
rect 521370 23218 521412 23454
rect 521092 23134 521412 23218
rect 521092 22898 521134 23134
rect 521370 22898 521412 23134
rect 521092 22866 521412 22898
rect 525040 23454 525360 23486
rect 525040 23218 525082 23454
rect 525318 23218 525360 23454
rect 525040 23134 525360 23218
rect 525040 22898 525082 23134
rect 525318 22898 525360 23134
rect 525040 22866 525360 22898
rect 429331 13428 429397 13429
rect 429331 13364 429332 13428
rect 429396 13364 429397 13428
rect 429331 13363 429397 13364
rect 397683 13292 397749 13293
rect 397683 13228 397684 13292
rect 397748 13228 397749 13292
rect 397683 13227 397749 13228
rect 169707 13156 169773 13157
rect 169707 13092 169708 13156
rect 169772 13092 169773 13156
rect 169707 13091 169773 13092
rect 527406 13021 527466 699755
rect 541994 698454 542614 705242
rect 541994 698218 542026 698454
rect 542262 698218 542346 698454
rect 542582 698218 542614 698454
rect 541994 698134 542614 698218
rect 541994 697898 542026 698134
rect 542262 697898 542346 698134
rect 542582 697898 542614 698134
rect 541994 671454 542614 697898
rect 541994 671218 542026 671454
rect 542262 671218 542346 671454
rect 542582 671218 542614 671454
rect 541994 671134 542614 671218
rect 541994 670898 542026 671134
rect 542262 670898 542346 671134
rect 542582 670898 542614 671134
rect 541994 644454 542614 670898
rect 541994 644218 542026 644454
rect 542262 644218 542346 644454
rect 542582 644218 542614 644454
rect 541994 644134 542614 644218
rect 541994 643898 542026 644134
rect 542262 643898 542346 644134
rect 542582 643898 542614 644134
rect 541994 617454 542614 643898
rect 541994 617218 542026 617454
rect 542262 617218 542346 617454
rect 542582 617218 542614 617454
rect 541994 617134 542614 617218
rect 541994 616898 542026 617134
rect 542262 616898 542346 617134
rect 542582 616898 542614 617134
rect 541994 590454 542614 616898
rect 541994 590218 542026 590454
rect 542262 590218 542346 590454
rect 542582 590218 542614 590454
rect 541994 590134 542614 590218
rect 541994 589898 542026 590134
rect 542262 589898 542346 590134
rect 542582 589898 542614 590134
rect 541994 563454 542614 589898
rect 541994 563218 542026 563454
rect 542262 563218 542346 563454
rect 542582 563218 542614 563454
rect 541994 563134 542614 563218
rect 541994 562898 542026 563134
rect 542262 562898 542346 563134
rect 542582 562898 542614 563134
rect 541994 536454 542614 562898
rect 541994 536218 542026 536454
rect 542262 536218 542346 536454
rect 542582 536218 542614 536454
rect 541994 536134 542614 536218
rect 541994 535898 542026 536134
rect 542262 535898 542346 536134
rect 542582 535898 542614 536134
rect 541994 509454 542614 535898
rect 541994 509218 542026 509454
rect 542262 509218 542346 509454
rect 542582 509218 542614 509454
rect 541994 509134 542614 509218
rect 541994 508898 542026 509134
rect 542262 508898 542346 509134
rect 542582 508898 542614 509134
rect 541994 482454 542614 508898
rect 541994 482218 542026 482454
rect 542262 482218 542346 482454
rect 542582 482218 542614 482454
rect 541994 482134 542614 482218
rect 541994 481898 542026 482134
rect 542262 481898 542346 482134
rect 542582 481898 542614 482134
rect 541994 455454 542614 481898
rect 541994 455218 542026 455454
rect 542262 455218 542346 455454
rect 542582 455218 542614 455454
rect 541994 455134 542614 455218
rect 541994 454898 542026 455134
rect 542262 454898 542346 455134
rect 542582 454898 542614 455134
rect 541994 428454 542614 454898
rect 541994 428218 542026 428454
rect 542262 428218 542346 428454
rect 542582 428218 542614 428454
rect 541994 428134 542614 428218
rect 541994 427898 542026 428134
rect 542262 427898 542346 428134
rect 542582 427898 542614 428134
rect 541994 401454 542614 427898
rect 541994 401218 542026 401454
rect 542262 401218 542346 401454
rect 542582 401218 542614 401454
rect 541994 401134 542614 401218
rect 541994 400898 542026 401134
rect 542262 400898 542346 401134
rect 542582 400898 542614 401134
rect 541994 374454 542614 400898
rect 541994 374218 542026 374454
rect 542262 374218 542346 374454
rect 542582 374218 542614 374454
rect 541994 374134 542614 374218
rect 541994 373898 542026 374134
rect 542262 373898 542346 374134
rect 542582 373898 542614 374134
rect 541994 347454 542614 373898
rect 541994 347218 542026 347454
rect 542262 347218 542346 347454
rect 542582 347218 542614 347454
rect 541994 347134 542614 347218
rect 541994 346898 542026 347134
rect 542262 346898 542346 347134
rect 542582 346898 542614 347134
rect 541994 320454 542614 346898
rect 541994 320218 542026 320454
rect 542262 320218 542346 320454
rect 542582 320218 542614 320454
rect 541994 320134 542614 320218
rect 541994 319898 542026 320134
rect 542262 319898 542346 320134
rect 542582 319898 542614 320134
rect 541994 293454 542614 319898
rect 541994 293218 542026 293454
rect 542262 293218 542346 293454
rect 542582 293218 542614 293454
rect 541994 293134 542614 293218
rect 541994 292898 542026 293134
rect 542262 292898 542346 293134
rect 542582 292898 542614 293134
rect 541994 266454 542614 292898
rect 541994 266218 542026 266454
rect 542262 266218 542346 266454
rect 542582 266218 542614 266454
rect 541994 266134 542614 266218
rect 541994 265898 542026 266134
rect 542262 265898 542346 266134
rect 542582 265898 542614 266134
rect 541994 239454 542614 265898
rect 541994 239218 542026 239454
rect 542262 239218 542346 239454
rect 542582 239218 542614 239454
rect 541994 239134 542614 239218
rect 541994 238898 542026 239134
rect 542262 238898 542346 239134
rect 542582 238898 542614 239134
rect 541994 212454 542614 238898
rect 541994 212218 542026 212454
rect 542262 212218 542346 212454
rect 542582 212218 542614 212454
rect 541994 212134 542614 212218
rect 541994 211898 542026 212134
rect 542262 211898 542346 212134
rect 542582 211898 542614 212134
rect 541994 185454 542614 211898
rect 541994 185218 542026 185454
rect 542262 185218 542346 185454
rect 542582 185218 542614 185454
rect 541994 185134 542614 185218
rect 541994 184898 542026 185134
rect 542262 184898 542346 185134
rect 542582 184898 542614 185134
rect 541994 158454 542614 184898
rect 541994 158218 542026 158454
rect 542262 158218 542346 158454
rect 542582 158218 542614 158454
rect 541994 158134 542614 158218
rect 541994 157898 542026 158134
rect 542262 157898 542346 158134
rect 542582 157898 542614 158134
rect 541994 131454 542614 157898
rect 541994 131218 542026 131454
rect 542262 131218 542346 131454
rect 542582 131218 542614 131454
rect 541994 131134 542614 131218
rect 541994 130898 542026 131134
rect 542262 130898 542346 131134
rect 542582 130898 542614 131134
rect 541994 104454 542614 130898
rect 541994 104218 542026 104454
rect 542262 104218 542346 104454
rect 542582 104218 542614 104454
rect 541994 104134 542614 104218
rect 541994 103898 542026 104134
rect 542262 103898 542346 104134
rect 542582 103898 542614 104134
rect 541994 77454 542614 103898
rect 541994 77218 542026 77454
rect 542262 77218 542346 77454
rect 542582 77218 542614 77454
rect 541994 77134 542614 77218
rect 541994 76898 542026 77134
rect 542262 76898 542346 77134
rect 542582 76898 542614 77134
rect 541994 69000 542614 76898
rect 545494 704838 546114 711590
rect 545494 704602 545526 704838
rect 545762 704602 545846 704838
rect 546082 704602 546114 704838
rect 545494 704518 546114 704602
rect 545494 704282 545526 704518
rect 545762 704282 545846 704518
rect 546082 704282 546114 704518
rect 545494 701829 546114 704282
rect 545494 701593 545526 701829
rect 545762 701593 545846 701829
rect 546082 701593 546114 701829
rect 545494 701509 546114 701593
rect 545494 701273 545526 701509
rect 545762 701273 545846 701509
rect 546082 701273 546114 701509
rect 545494 674829 546114 701273
rect 569994 705798 570614 711590
rect 569994 705562 570026 705798
rect 570262 705562 570346 705798
rect 570582 705562 570614 705798
rect 569994 705478 570614 705562
rect 569994 705242 570026 705478
rect 570262 705242 570346 705478
rect 570582 705242 570614 705478
rect 558867 699820 558933 699821
rect 558867 699756 558868 699820
rect 558932 699756 558933 699820
rect 558867 699755 558933 699756
rect 545494 674593 545526 674829
rect 545762 674593 545846 674829
rect 546082 674593 546114 674829
rect 545494 674509 546114 674593
rect 545494 674273 545526 674509
rect 545762 674273 545846 674509
rect 546082 674273 546114 674509
rect 545494 647829 546114 674273
rect 545494 647593 545526 647829
rect 545762 647593 545846 647829
rect 546082 647593 546114 647829
rect 545494 647509 546114 647593
rect 545494 647273 545526 647509
rect 545762 647273 545846 647509
rect 546082 647273 546114 647509
rect 545494 620829 546114 647273
rect 545494 620593 545526 620829
rect 545762 620593 545846 620829
rect 546082 620593 546114 620829
rect 545494 620509 546114 620593
rect 545494 620273 545526 620509
rect 545762 620273 545846 620509
rect 546082 620273 546114 620509
rect 545494 593829 546114 620273
rect 545494 593593 545526 593829
rect 545762 593593 545846 593829
rect 546082 593593 546114 593829
rect 545494 593509 546114 593593
rect 545494 593273 545526 593509
rect 545762 593273 545846 593509
rect 546082 593273 546114 593509
rect 545494 566829 546114 593273
rect 545494 566593 545526 566829
rect 545762 566593 545846 566829
rect 546082 566593 546114 566829
rect 545494 566509 546114 566593
rect 545494 566273 545526 566509
rect 545762 566273 545846 566509
rect 546082 566273 546114 566509
rect 545494 539829 546114 566273
rect 545494 539593 545526 539829
rect 545762 539593 545846 539829
rect 546082 539593 546114 539829
rect 545494 539509 546114 539593
rect 545494 539273 545526 539509
rect 545762 539273 545846 539509
rect 546082 539273 546114 539509
rect 545494 512829 546114 539273
rect 545494 512593 545526 512829
rect 545762 512593 545846 512829
rect 546082 512593 546114 512829
rect 545494 512509 546114 512593
rect 545494 512273 545526 512509
rect 545762 512273 545846 512509
rect 546082 512273 546114 512509
rect 545494 485829 546114 512273
rect 545494 485593 545526 485829
rect 545762 485593 545846 485829
rect 546082 485593 546114 485829
rect 545494 485509 546114 485593
rect 545494 485273 545526 485509
rect 545762 485273 545846 485509
rect 546082 485273 546114 485509
rect 545494 458829 546114 485273
rect 545494 458593 545526 458829
rect 545762 458593 545846 458829
rect 546082 458593 546114 458829
rect 545494 458509 546114 458593
rect 545494 458273 545526 458509
rect 545762 458273 545846 458509
rect 546082 458273 546114 458509
rect 545494 431829 546114 458273
rect 545494 431593 545526 431829
rect 545762 431593 545846 431829
rect 546082 431593 546114 431829
rect 545494 431509 546114 431593
rect 545494 431273 545526 431509
rect 545762 431273 545846 431509
rect 546082 431273 546114 431509
rect 545494 404829 546114 431273
rect 545494 404593 545526 404829
rect 545762 404593 545846 404829
rect 546082 404593 546114 404829
rect 545494 404509 546114 404593
rect 545494 404273 545526 404509
rect 545762 404273 545846 404509
rect 546082 404273 546114 404509
rect 545494 377829 546114 404273
rect 545494 377593 545526 377829
rect 545762 377593 545846 377829
rect 546082 377593 546114 377829
rect 545494 377509 546114 377593
rect 545494 377273 545526 377509
rect 545762 377273 545846 377509
rect 546082 377273 546114 377509
rect 545494 350829 546114 377273
rect 545494 350593 545526 350829
rect 545762 350593 545846 350829
rect 546082 350593 546114 350829
rect 545494 350509 546114 350593
rect 545494 350273 545526 350509
rect 545762 350273 545846 350509
rect 546082 350273 546114 350509
rect 545494 323829 546114 350273
rect 545494 323593 545526 323829
rect 545762 323593 545846 323829
rect 546082 323593 546114 323829
rect 545494 323509 546114 323593
rect 545494 323273 545526 323509
rect 545762 323273 545846 323509
rect 546082 323273 546114 323509
rect 545494 296829 546114 323273
rect 545494 296593 545526 296829
rect 545762 296593 545846 296829
rect 546082 296593 546114 296829
rect 545494 296509 546114 296593
rect 545494 296273 545526 296509
rect 545762 296273 545846 296509
rect 546082 296273 546114 296509
rect 545494 269829 546114 296273
rect 545494 269593 545526 269829
rect 545762 269593 545846 269829
rect 546082 269593 546114 269829
rect 545494 269509 546114 269593
rect 545494 269273 545526 269509
rect 545762 269273 545846 269509
rect 546082 269273 546114 269509
rect 545494 242829 546114 269273
rect 545494 242593 545526 242829
rect 545762 242593 545846 242829
rect 546082 242593 546114 242829
rect 545494 242509 546114 242593
rect 545494 242273 545526 242509
rect 545762 242273 545846 242509
rect 546082 242273 546114 242509
rect 545494 215829 546114 242273
rect 545494 215593 545526 215829
rect 545762 215593 545846 215829
rect 546082 215593 546114 215829
rect 545494 215509 546114 215593
rect 545494 215273 545526 215509
rect 545762 215273 545846 215509
rect 546082 215273 546114 215509
rect 545494 188829 546114 215273
rect 545494 188593 545526 188829
rect 545762 188593 545846 188829
rect 546082 188593 546114 188829
rect 545494 188509 546114 188593
rect 545494 188273 545526 188509
rect 545762 188273 545846 188509
rect 546082 188273 546114 188509
rect 545494 161829 546114 188273
rect 545494 161593 545526 161829
rect 545762 161593 545846 161829
rect 546082 161593 546114 161829
rect 545494 161509 546114 161593
rect 545494 161273 545526 161509
rect 545762 161273 545846 161509
rect 546082 161273 546114 161509
rect 545494 134829 546114 161273
rect 545494 134593 545526 134829
rect 545762 134593 545846 134829
rect 546082 134593 546114 134829
rect 545494 134509 546114 134593
rect 545494 134273 545526 134509
rect 545762 134273 545846 134509
rect 546082 134273 546114 134509
rect 545494 107829 546114 134273
rect 545494 107593 545526 107829
rect 545762 107593 545846 107829
rect 546082 107593 546114 107829
rect 545494 107509 546114 107593
rect 545494 107273 545526 107509
rect 545762 107273 545846 107509
rect 546082 107273 546114 107509
rect 545494 80829 546114 107273
rect 545494 80593 545526 80829
rect 545762 80593 545846 80829
rect 546082 80593 546114 80829
rect 545494 80509 546114 80593
rect 545494 80273 545526 80509
rect 545762 80273 545846 80509
rect 546082 80273 546114 80509
rect 545494 69000 546114 80273
rect 532218 53829 532538 53861
rect 532218 53593 532260 53829
rect 532496 53593 532538 53829
rect 532218 53509 532538 53593
rect 532218 53273 532260 53509
rect 532496 53273 532538 53509
rect 532218 53241 532538 53273
rect 533166 53829 533486 53861
rect 533166 53593 533208 53829
rect 533444 53593 533486 53829
rect 533166 53509 533486 53593
rect 533166 53273 533208 53509
rect 533444 53273 533486 53509
rect 533166 53241 533486 53273
rect 534114 53829 534434 53861
rect 534114 53593 534156 53829
rect 534392 53593 534434 53829
rect 534114 53509 534434 53593
rect 534114 53273 534156 53509
rect 534392 53273 534434 53509
rect 534114 53241 534434 53273
rect 535062 53829 535382 53861
rect 535062 53593 535104 53829
rect 535340 53593 535382 53829
rect 535062 53509 535382 53593
rect 535062 53273 535104 53509
rect 535340 53273 535382 53509
rect 535062 53241 535382 53273
rect 540918 53829 541238 53861
rect 540918 53593 540960 53829
rect 541196 53593 541238 53829
rect 540918 53509 541238 53593
rect 540918 53273 540960 53509
rect 541196 53273 541238 53509
rect 540918 53241 541238 53273
rect 544866 53829 545186 53861
rect 544866 53593 544908 53829
rect 545144 53593 545186 53829
rect 544866 53509 545186 53593
rect 544866 53273 544908 53509
rect 545144 53273 545186 53509
rect 544866 53241 545186 53273
rect 548814 53829 549134 53861
rect 548814 53593 548856 53829
rect 549092 53593 549134 53829
rect 548814 53509 549134 53593
rect 548814 53273 548856 53509
rect 549092 53273 549134 53509
rect 548814 53241 549134 53273
rect 552762 53829 553082 53861
rect 552762 53593 552804 53829
rect 553040 53593 553082 53829
rect 552762 53509 553082 53593
rect 552762 53273 552804 53509
rect 553040 53273 553082 53509
rect 552762 53241 553082 53273
rect 532692 50454 533012 50486
rect 532692 50218 532734 50454
rect 532970 50218 533012 50454
rect 532692 50134 533012 50218
rect 532692 49898 532734 50134
rect 532970 49898 533012 50134
rect 532692 49866 533012 49898
rect 533640 50454 533960 50486
rect 533640 50218 533682 50454
rect 533918 50218 533960 50454
rect 533640 50134 533960 50218
rect 533640 49898 533682 50134
rect 533918 49898 533960 50134
rect 533640 49866 533960 49898
rect 534588 50454 534908 50486
rect 534588 50218 534630 50454
rect 534866 50218 534908 50454
rect 534588 50134 534908 50218
rect 534588 49898 534630 50134
rect 534866 49898 534908 50134
rect 534588 49866 534908 49898
rect 542892 50454 543212 50486
rect 542892 50218 542934 50454
rect 543170 50218 543212 50454
rect 542892 50134 543212 50218
rect 542892 49898 542934 50134
rect 543170 49898 543212 50134
rect 542892 49866 543212 49898
rect 546840 50454 547160 50486
rect 546840 50218 546882 50454
rect 547118 50218 547160 50454
rect 546840 50134 547160 50218
rect 546840 49898 546882 50134
rect 547118 49898 547160 50134
rect 546840 49866 547160 49898
rect 550788 50454 551108 50486
rect 550788 50218 550830 50454
rect 551066 50218 551108 50454
rect 550788 50134 551108 50218
rect 550788 49898 550830 50134
rect 551066 49898 551108 50134
rect 550788 49866 551108 49898
rect 530962 26829 531282 26861
rect 530962 26593 531004 26829
rect 531240 26593 531282 26829
rect 530962 26509 531282 26593
rect 530962 26273 531004 26509
rect 531240 26273 531282 26509
rect 530962 26241 531282 26273
rect 539418 26829 539738 26861
rect 539418 26593 539460 26829
rect 539696 26593 539738 26829
rect 539418 26509 539738 26593
rect 539418 26273 539460 26509
rect 539696 26273 539738 26509
rect 539418 26241 539738 26273
rect 540366 26829 540686 26861
rect 540366 26593 540408 26829
rect 540644 26593 540686 26829
rect 540366 26509 540686 26593
rect 540366 26273 540408 26509
rect 540644 26273 540686 26509
rect 540366 26241 540686 26273
rect 541314 26829 541634 26861
rect 541314 26593 541356 26829
rect 541592 26593 541634 26829
rect 541314 26509 541634 26593
rect 541314 26273 541356 26509
rect 541592 26273 541634 26509
rect 541314 26241 541634 26273
rect 542262 26829 542582 26861
rect 542262 26593 542304 26829
rect 542540 26593 542582 26829
rect 542262 26509 542582 26593
rect 542262 26273 542304 26509
rect 542540 26273 542582 26509
rect 542262 26241 542582 26273
rect 548118 26829 548438 26861
rect 548118 26593 548160 26829
rect 548396 26593 548438 26829
rect 548118 26509 548438 26593
rect 548118 26273 548160 26509
rect 548396 26273 548438 26509
rect 548118 26241 548438 26273
rect 552066 26829 552386 26861
rect 552066 26593 552108 26829
rect 552344 26593 552386 26829
rect 552066 26509 552386 26593
rect 552066 26273 552108 26509
rect 552344 26273 552386 26509
rect 552066 26241 552386 26273
rect 556014 26829 556334 26861
rect 556014 26593 556056 26829
rect 556292 26593 556334 26829
rect 556014 26509 556334 26593
rect 556014 26273 556056 26509
rect 556292 26273 556334 26509
rect 556014 26241 556334 26273
rect 528988 23454 529308 23486
rect 528988 23218 529030 23454
rect 529266 23218 529308 23454
rect 528988 23134 529308 23218
rect 528988 22898 529030 23134
rect 529266 22898 529308 23134
rect 528988 22866 529308 22898
rect 539892 23454 540212 23486
rect 539892 23218 539934 23454
rect 540170 23218 540212 23454
rect 539892 23134 540212 23218
rect 539892 22898 539934 23134
rect 540170 22898 540212 23134
rect 539892 22866 540212 22898
rect 540840 23454 541160 23486
rect 540840 23218 540882 23454
rect 541118 23218 541160 23454
rect 540840 23134 541160 23218
rect 540840 22898 540882 23134
rect 541118 22898 541160 23134
rect 540840 22866 541160 22898
rect 541788 23454 542108 23486
rect 541788 23218 541830 23454
rect 542066 23218 542108 23454
rect 541788 23134 542108 23218
rect 541788 22898 541830 23134
rect 542066 22898 542108 23134
rect 541788 22866 542108 22898
rect 550092 23454 550412 23486
rect 550092 23218 550134 23454
rect 550370 23218 550412 23454
rect 550092 23134 550412 23218
rect 550092 22898 550134 23134
rect 550370 22898 550412 23134
rect 550092 22866 550412 22898
rect 554040 23454 554360 23486
rect 554040 23218 554082 23454
rect 554318 23218 554360 23454
rect 554040 23134 554360 23218
rect 554040 22898 554082 23134
rect 554318 22898 554360 23134
rect 554040 22866 554360 22898
rect 557988 23454 558308 23486
rect 557988 23218 558030 23454
rect 558266 23218 558308 23454
rect 557988 23134 558308 23218
rect 557988 22898 558030 23134
rect 558266 22898 558308 23134
rect 557988 22866 558308 22898
rect 558870 13565 558930 699755
rect 569994 698454 570614 705242
rect 569994 698218 570026 698454
rect 570262 698218 570346 698454
rect 570582 698218 570614 698454
rect 569994 698134 570614 698218
rect 569994 697898 570026 698134
rect 570262 697898 570346 698134
rect 570582 697898 570614 698134
rect 569994 671454 570614 697898
rect 569994 671218 570026 671454
rect 570262 671218 570346 671454
rect 570582 671218 570614 671454
rect 569994 671134 570614 671218
rect 569994 670898 570026 671134
rect 570262 670898 570346 671134
rect 570582 670898 570614 671134
rect 569994 644454 570614 670898
rect 569994 644218 570026 644454
rect 570262 644218 570346 644454
rect 570582 644218 570614 644454
rect 569994 644134 570614 644218
rect 569994 643898 570026 644134
rect 570262 643898 570346 644134
rect 570582 643898 570614 644134
rect 569994 617454 570614 643898
rect 569994 617218 570026 617454
rect 570262 617218 570346 617454
rect 570582 617218 570614 617454
rect 569994 617134 570614 617218
rect 569994 616898 570026 617134
rect 570262 616898 570346 617134
rect 570582 616898 570614 617134
rect 569994 590454 570614 616898
rect 569994 590218 570026 590454
rect 570262 590218 570346 590454
rect 570582 590218 570614 590454
rect 569994 590134 570614 590218
rect 569994 589898 570026 590134
rect 570262 589898 570346 590134
rect 570582 589898 570614 590134
rect 569994 563454 570614 589898
rect 569994 563218 570026 563454
rect 570262 563218 570346 563454
rect 570582 563218 570614 563454
rect 569994 563134 570614 563218
rect 569994 562898 570026 563134
rect 570262 562898 570346 563134
rect 570582 562898 570614 563134
rect 569994 536454 570614 562898
rect 569994 536218 570026 536454
rect 570262 536218 570346 536454
rect 570582 536218 570614 536454
rect 569994 536134 570614 536218
rect 569994 535898 570026 536134
rect 570262 535898 570346 536134
rect 570582 535898 570614 536134
rect 569994 509454 570614 535898
rect 569994 509218 570026 509454
rect 570262 509218 570346 509454
rect 570582 509218 570614 509454
rect 569994 509134 570614 509218
rect 569994 508898 570026 509134
rect 570262 508898 570346 509134
rect 570582 508898 570614 509134
rect 569994 482454 570614 508898
rect 569994 482218 570026 482454
rect 570262 482218 570346 482454
rect 570582 482218 570614 482454
rect 569994 482134 570614 482218
rect 569994 481898 570026 482134
rect 570262 481898 570346 482134
rect 570582 481898 570614 482134
rect 569994 455454 570614 481898
rect 569994 455218 570026 455454
rect 570262 455218 570346 455454
rect 570582 455218 570614 455454
rect 569994 455134 570614 455218
rect 569994 454898 570026 455134
rect 570262 454898 570346 455134
rect 570582 454898 570614 455134
rect 569994 428454 570614 454898
rect 569994 428218 570026 428454
rect 570262 428218 570346 428454
rect 570582 428218 570614 428454
rect 569994 428134 570614 428218
rect 569994 427898 570026 428134
rect 570262 427898 570346 428134
rect 570582 427898 570614 428134
rect 569994 401454 570614 427898
rect 569994 401218 570026 401454
rect 570262 401218 570346 401454
rect 570582 401218 570614 401454
rect 569994 401134 570614 401218
rect 569994 400898 570026 401134
rect 570262 400898 570346 401134
rect 570582 400898 570614 401134
rect 569994 374454 570614 400898
rect 569994 374218 570026 374454
rect 570262 374218 570346 374454
rect 570582 374218 570614 374454
rect 569994 374134 570614 374218
rect 569994 373898 570026 374134
rect 570262 373898 570346 374134
rect 570582 373898 570614 374134
rect 569994 347454 570614 373898
rect 569994 347218 570026 347454
rect 570262 347218 570346 347454
rect 570582 347218 570614 347454
rect 569994 347134 570614 347218
rect 569994 346898 570026 347134
rect 570262 346898 570346 347134
rect 570582 346898 570614 347134
rect 569994 320454 570614 346898
rect 569994 320218 570026 320454
rect 570262 320218 570346 320454
rect 570582 320218 570614 320454
rect 569994 320134 570614 320218
rect 569994 319898 570026 320134
rect 570262 319898 570346 320134
rect 570582 319898 570614 320134
rect 569994 293454 570614 319898
rect 569994 293218 570026 293454
rect 570262 293218 570346 293454
rect 570582 293218 570614 293454
rect 569994 293134 570614 293218
rect 569994 292898 570026 293134
rect 570262 292898 570346 293134
rect 570582 292898 570614 293134
rect 569994 266454 570614 292898
rect 569994 266218 570026 266454
rect 570262 266218 570346 266454
rect 570582 266218 570614 266454
rect 569994 266134 570614 266218
rect 569994 265898 570026 266134
rect 570262 265898 570346 266134
rect 570582 265898 570614 266134
rect 569994 239454 570614 265898
rect 569994 239218 570026 239454
rect 570262 239218 570346 239454
rect 570582 239218 570614 239454
rect 569994 239134 570614 239218
rect 569994 238898 570026 239134
rect 570262 238898 570346 239134
rect 570582 238898 570614 239134
rect 569994 212454 570614 238898
rect 569994 212218 570026 212454
rect 570262 212218 570346 212454
rect 570582 212218 570614 212454
rect 569994 212134 570614 212218
rect 569994 211898 570026 212134
rect 570262 211898 570346 212134
rect 570582 211898 570614 212134
rect 569994 185454 570614 211898
rect 569994 185218 570026 185454
rect 570262 185218 570346 185454
rect 570582 185218 570614 185454
rect 569994 185134 570614 185218
rect 569994 184898 570026 185134
rect 570262 184898 570346 185134
rect 570582 184898 570614 185134
rect 569994 158454 570614 184898
rect 569994 158218 570026 158454
rect 570262 158218 570346 158454
rect 570582 158218 570614 158454
rect 569994 158134 570614 158218
rect 569994 157898 570026 158134
rect 570262 157898 570346 158134
rect 570582 157898 570614 158134
rect 569994 131454 570614 157898
rect 569994 131218 570026 131454
rect 570262 131218 570346 131454
rect 570582 131218 570614 131454
rect 569994 131134 570614 131218
rect 569994 130898 570026 131134
rect 570262 130898 570346 131134
rect 570582 130898 570614 131134
rect 569994 104454 570614 130898
rect 569994 104218 570026 104454
rect 570262 104218 570346 104454
rect 570582 104218 570614 104454
rect 569994 104134 570614 104218
rect 569994 103898 570026 104134
rect 570262 103898 570346 104134
rect 570582 103898 570614 104134
rect 569994 77454 570614 103898
rect 569994 77218 570026 77454
rect 570262 77218 570346 77454
rect 570582 77218 570614 77454
rect 569994 77134 570614 77218
rect 569994 76898 570026 77134
rect 570262 76898 570346 77134
rect 570582 76898 570614 77134
rect 561218 53829 561538 53861
rect 561218 53593 561260 53829
rect 561496 53593 561538 53829
rect 561218 53509 561538 53593
rect 561218 53273 561260 53509
rect 561496 53273 561538 53509
rect 561218 53241 561538 53273
rect 562166 53829 562486 53861
rect 562166 53593 562208 53829
rect 562444 53593 562486 53829
rect 562166 53509 562486 53593
rect 562166 53273 562208 53509
rect 562444 53273 562486 53509
rect 562166 53241 562486 53273
rect 563114 53829 563434 53861
rect 563114 53593 563156 53829
rect 563392 53593 563434 53829
rect 563114 53509 563434 53593
rect 563114 53273 563156 53509
rect 563392 53273 563434 53509
rect 563114 53241 563434 53273
rect 564062 53829 564382 53861
rect 564062 53593 564104 53829
rect 564340 53593 564382 53829
rect 564062 53509 564382 53593
rect 564062 53273 564104 53509
rect 564340 53273 564382 53509
rect 564062 53241 564382 53273
rect 561692 50454 562012 50486
rect 561692 50218 561734 50454
rect 561970 50218 562012 50454
rect 561692 50134 562012 50218
rect 561692 49898 561734 50134
rect 561970 49898 562012 50134
rect 561692 49866 562012 49898
rect 562640 50454 562960 50486
rect 562640 50218 562682 50454
rect 562918 50218 562960 50454
rect 562640 50134 562960 50218
rect 562640 49898 562682 50134
rect 562918 49898 562960 50134
rect 562640 49866 562960 49898
rect 563588 50454 563908 50486
rect 563588 50218 563630 50454
rect 563866 50218 563908 50454
rect 563588 50134 563908 50218
rect 563588 49898 563630 50134
rect 563866 49898 563908 50134
rect 563588 49866 563908 49898
rect 569994 50454 570614 76898
rect 569994 50218 570026 50454
rect 570262 50218 570346 50454
rect 570582 50218 570614 50454
rect 569994 50134 570614 50218
rect 569994 49898 570026 50134
rect 570262 49898 570346 50134
rect 570582 49898 570614 50134
rect 559962 26829 560282 26861
rect 559962 26593 560004 26829
rect 560240 26593 560282 26829
rect 559962 26509 560282 26593
rect 559962 26273 560004 26509
rect 560240 26273 560282 26509
rect 559962 26241 560282 26273
rect 569994 23454 570614 49898
rect 569994 23218 570026 23454
rect 570262 23218 570346 23454
rect 570582 23218 570614 23454
rect 569994 23134 570614 23218
rect 569994 22898 570026 23134
rect 570262 22898 570346 23134
rect 570582 22898 570614 23134
rect 558867 13564 558933 13565
rect 558867 13500 558868 13564
rect 558932 13500 558933 13564
rect 558867 13499 558933 13500
rect 527403 13020 527469 13021
rect 527403 12956 527404 13020
rect 527468 12956 527469 13020
rect 527403 12955 527469 12956
rect 69494 -582 69526 -346
rect 69762 -582 69846 -346
rect 70082 -582 70114 -346
rect 69494 -666 70114 -582
rect 69494 -902 69526 -666
rect 69762 -902 69846 -666
rect 70082 -902 70114 -666
rect 69494 -7654 70114 -902
rect 569994 -1306 570614 22898
rect 569994 -1542 570026 -1306
rect 570262 -1542 570346 -1306
rect 570582 -1542 570614 -1306
rect 569994 -1626 570614 -1542
rect 569994 -1862 570026 -1626
rect 570262 -1862 570346 -1626
rect 570582 -1862 570614 -1626
rect 569994 -7654 570614 -1862
rect 573494 704838 574114 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 573494 704602 573526 704838
rect 573762 704602 573846 704838
rect 574082 704602 574114 704838
rect 573494 704518 574114 704602
rect 573494 704282 573526 704518
rect 573762 704282 573846 704518
rect 574082 704282 574114 704518
rect 573494 701829 574114 704282
rect 573494 701593 573526 701829
rect 573762 701593 573846 701829
rect 574082 701593 574114 701829
rect 573494 701509 574114 701593
rect 573494 701273 573526 701509
rect 573762 701273 573846 701509
rect 574082 701273 574114 701509
rect 573494 674829 574114 701273
rect 573494 674593 573526 674829
rect 573762 674593 573846 674829
rect 574082 674593 574114 674829
rect 573494 674509 574114 674593
rect 573494 674273 573526 674509
rect 573762 674273 573846 674509
rect 574082 674273 574114 674509
rect 573494 647829 574114 674273
rect 573494 647593 573526 647829
rect 573762 647593 573846 647829
rect 574082 647593 574114 647829
rect 573494 647509 574114 647593
rect 573494 647273 573526 647509
rect 573762 647273 573846 647509
rect 574082 647273 574114 647509
rect 573494 620829 574114 647273
rect 573494 620593 573526 620829
rect 573762 620593 573846 620829
rect 574082 620593 574114 620829
rect 573494 620509 574114 620593
rect 573494 620273 573526 620509
rect 573762 620273 573846 620509
rect 574082 620273 574114 620509
rect 573494 593829 574114 620273
rect 573494 593593 573526 593829
rect 573762 593593 573846 593829
rect 574082 593593 574114 593829
rect 573494 593509 574114 593593
rect 573494 593273 573526 593509
rect 573762 593273 573846 593509
rect 574082 593273 574114 593509
rect 573494 566829 574114 593273
rect 573494 566593 573526 566829
rect 573762 566593 573846 566829
rect 574082 566593 574114 566829
rect 573494 566509 574114 566593
rect 573494 566273 573526 566509
rect 573762 566273 573846 566509
rect 574082 566273 574114 566509
rect 573494 539829 574114 566273
rect 573494 539593 573526 539829
rect 573762 539593 573846 539829
rect 574082 539593 574114 539829
rect 573494 539509 574114 539593
rect 573494 539273 573526 539509
rect 573762 539273 573846 539509
rect 574082 539273 574114 539509
rect 573494 512829 574114 539273
rect 573494 512593 573526 512829
rect 573762 512593 573846 512829
rect 574082 512593 574114 512829
rect 573494 512509 574114 512593
rect 573494 512273 573526 512509
rect 573762 512273 573846 512509
rect 574082 512273 574114 512509
rect 573494 485829 574114 512273
rect 573494 485593 573526 485829
rect 573762 485593 573846 485829
rect 574082 485593 574114 485829
rect 573494 485509 574114 485593
rect 573494 485273 573526 485509
rect 573762 485273 573846 485509
rect 574082 485273 574114 485509
rect 573494 458829 574114 485273
rect 573494 458593 573526 458829
rect 573762 458593 573846 458829
rect 574082 458593 574114 458829
rect 573494 458509 574114 458593
rect 573494 458273 573526 458509
rect 573762 458273 573846 458509
rect 574082 458273 574114 458509
rect 573494 431829 574114 458273
rect 573494 431593 573526 431829
rect 573762 431593 573846 431829
rect 574082 431593 574114 431829
rect 573494 431509 574114 431593
rect 573494 431273 573526 431509
rect 573762 431273 573846 431509
rect 574082 431273 574114 431509
rect 573494 404829 574114 431273
rect 573494 404593 573526 404829
rect 573762 404593 573846 404829
rect 574082 404593 574114 404829
rect 573494 404509 574114 404593
rect 573494 404273 573526 404509
rect 573762 404273 573846 404509
rect 574082 404273 574114 404509
rect 573494 377829 574114 404273
rect 573494 377593 573526 377829
rect 573762 377593 573846 377829
rect 574082 377593 574114 377829
rect 573494 377509 574114 377593
rect 573494 377273 573526 377509
rect 573762 377273 573846 377509
rect 574082 377273 574114 377509
rect 573494 350829 574114 377273
rect 573494 350593 573526 350829
rect 573762 350593 573846 350829
rect 574082 350593 574114 350829
rect 573494 350509 574114 350593
rect 573494 350273 573526 350509
rect 573762 350273 573846 350509
rect 574082 350273 574114 350509
rect 573494 323829 574114 350273
rect 573494 323593 573526 323829
rect 573762 323593 573846 323829
rect 574082 323593 574114 323829
rect 573494 323509 574114 323593
rect 573494 323273 573526 323509
rect 573762 323273 573846 323509
rect 574082 323273 574114 323509
rect 573494 296829 574114 323273
rect 573494 296593 573526 296829
rect 573762 296593 573846 296829
rect 574082 296593 574114 296829
rect 573494 296509 574114 296593
rect 573494 296273 573526 296509
rect 573762 296273 573846 296509
rect 574082 296273 574114 296509
rect 573494 269829 574114 296273
rect 573494 269593 573526 269829
rect 573762 269593 573846 269829
rect 574082 269593 574114 269829
rect 573494 269509 574114 269593
rect 573494 269273 573526 269509
rect 573762 269273 573846 269509
rect 574082 269273 574114 269509
rect 573494 242829 574114 269273
rect 573494 242593 573526 242829
rect 573762 242593 573846 242829
rect 574082 242593 574114 242829
rect 573494 242509 574114 242593
rect 573494 242273 573526 242509
rect 573762 242273 573846 242509
rect 574082 242273 574114 242509
rect 573494 215829 574114 242273
rect 573494 215593 573526 215829
rect 573762 215593 573846 215829
rect 574082 215593 574114 215829
rect 573494 215509 574114 215593
rect 573494 215273 573526 215509
rect 573762 215273 573846 215509
rect 574082 215273 574114 215509
rect 573494 188829 574114 215273
rect 573494 188593 573526 188829
rect 573762 188593 573846 188829
rect 574082 188593 574114 188829
rect 573494 188509 574114 188593
rect 573494 188273 573526 188509
rect 573762 188273 573846 188509
rect 574082 188273 574114 188509
rect 573494 161829 574114 188273
rect 573494 161593 573526 161829
rect 573762 161593 573846 161829
rect 574082 161593 574114 161829
rect 573494 161509 574114 161593
rect 573494 161273 573526 161509
rect 573762 161273 573846 161509
rect 574082 161273 574114 161509
rect 573494 134829 574114 161273
rect 573494 134593 573526 134829
rect 573762 134593 573846 134829
rect 574082 134593 574114 134829
rect 573494 134509 574114 134593
rect 573494 134273 573526 134509
rect 573762 134273 573846 134509
rect 574082 134273 574114 134509
rect 573494 107829 574114 134273
rect 573494 107593 573526 107829
rect 573762 107593 573846 107829
rect 574082 107593 574114 107829
rect 573494 107509 574114 107593
rect 573494 107273 573526 107509
rect 573762 107273 573846 107509
rect 574082 107273 574114 107509
rect 573494 80829 574114 107273
rect 573494 80593 573526 80829
rect 573762 80593 573846 80829
rect 574082 80593 574114 80829
rect 573494 80509 574114 80593
rect 573494 80273 573526 80509
rect 573762 80273 573846 80509
rect 574082 80273 574114 80509
rect 573494 53829 574114 80273
rect 573494 53593 573526 53829
rect 573762 53593 573846 53829
rect 574082 53593 574114 53829
rect 573494 53509 574114 53593
rect 573494 53273 573526 53509
rect 573762 53273 573846 53509
rect 574082 53273 574114 53509
rect 573494 26829 574114 53273
rect 573494 26593 573526 26829
rect 573762 26593 573846 26829
rect 574082 26593 574114 26829
rect 573494 26509 574114 26593
rect 573494 26273 573526 26509
rect 573762 26273 573846 26509
rect 574082 26273 574114 26509
rect 573494 -346 574114 26273
rect 573494 -582 573526 -346
rect 573762 -582 573846 -346
rect 574082 -582 574114 -346
rect 573494 -666 574114 -582
rect 573494 -902 573526 -666
rect 573762 -902 573846 -666
rect 574082 -902 574114 -666
rect 573494 -7654 574114 -902
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 701829 585930 704282
rect 585310 701593 585342 701829
rect 585578 701593 585662 701829
rect 585898 701593 585930 701829
rect 585310 701509 585930 701593
rect 585310 701273 585342 701509
rect 585578 701273 585662 701509
rect 585898 701273 585930 701509
rect 585310 674829 585930 701273
rect 585310 674593 585342 674829
rect 585578 674593 585662 674829
rect 585898 674593 585930 674829
rect 585310 674509 585930 674593
rect 585310 674273 585342 674509
rect 585578 674273 585662 674509
rect 585898 674273 585930 674509
rect 585310 647829 585930 674273
rect 585310 647593 585342 647829
rect 585578 647593 585662 647829
rect 585898 647593 585930 647829
rect 585310 647509 585930 647593
rect 585310 647273 585342 647509
rect 585578 647273 585662 647509
rect 585898 647273 585930 647509
rect 585310 620829 585930 647273
rect 585310 620593 585342 620829
rect 585578 620593 585662 620829
rect 585898 620593 585930 620829
rect 585310 620509 585930 620593
rect 585310 620273 585342 620509
rect 585578 620273 585662 620509
rect 585898 620273 585930 620509
rect 585310 593829 585930 620273
rect 585310 593593 585342 593829
rect 585578 593593 585662 593829
rect 585898 593593 585930 593829
rect 585310 593509 585930 593593
rect 585310 593273 585342 593509
rect 585578 593273 585662 593509
rect 585898 593273 585930 593509
rect 585310 566829 585930 593273
rect 585310 566593 585342 566829
rect 585578 566593 585662 566829
rect 585898 566593 585930 566829
rect 585310 566509 585930 566593
rect 585310 566273 585342 566509
rect 585578 566273 585662 566509
rect 585898 566273 585930 566509
rect 585310 539829 585930 566273
rect 585310 539593 585342 539829
rect 585578 539593 585662 539829
rect 585898 539593 585930 539829
rect 585310 539509 585930 539593
rect 585310 539273 585342 539509
rect 585578 539273 585662 539509
rect 585898 539273 585930 539509
rect 585310 512829 585930 539273
rect 585310 512593 585342 512829
rect 585578 512593 585662 512829
rect 585898 512593 585930 512829
rect 585310 512509 585930 512593
rect 585310 512273 585342 512509
rect 585578 512273 585662 512509
rect 585898 512273 585930 512509
rect 585310 485829 585930 512273
rect 585310 485593 585342 485829
rect 585578 485593 585662 485829
rect 585898 485593 585930 485829
rect 585310 485509 585930 485593
rect 585310 485273 585342 485509
rect 585578 485273 585662 485509
rect 585898 485273 585930 485509
rect 585310 458829 585930 485273
rect 585310 458593 585342 458829
rect 585578 458593 585662 458829
rect 585898 458593 585930 458829
rect 585310 458509 585930 458593
rect 585310 458273 585342 458509
rect 585578 458273 585662 458509
rect 585898 458273 585930 458509
rect 585310 431829 585930 458273
rect 585310 431593 585342 431829
rect 585578 431593 585662 431829
rect 585898 431593 585930 431829
rect 585310 431509 585930 431593
rect 585310 431273 585342 431509
rect 585578 431273 585662 431509
rect 585898 431273 585930 431509
rect 585310 404829 585930 431273
rect 585310 404593 585342 404829
rect 585578 404593 585662 404829
rect 585898 404593 585930 404829
rect 585310 404509 585930 404593
rect 585310 404273 585342 404509
rect 585578 404273 585662 404509
rect 585898 404273 585930 404509
rect 585310 377829 585930 404273
rect 585310 377593 585342 377829
rect 585578 377593 585662 377829
rect 585898 377593 585930 377829
rect 585310 377509 585930 377593
rect 585310 377273 585342 377509
rect 585578 377273 585662 377509
rect 585898 377273 585930 377509
rect 585310 350829 585930 377273
rect 585310 350593 585342 350829
rect 585578 350593 585662 350829
rect 585898 350593 585930 350829
rect 585310 350509 585930 350593
rect 585310 350273 585342 350509
rect 585578 350273 585662 350509
rect 585898 350273 585930 350509
rect 585310 323829 585930 350273
rect 585310 323593 585342 323829
rect 585578 323593 585662 323829
rect 585898 323593 585930 323829
rect 585310 323509 585930 323593
rect 585310 323273 585342 323509
rect 585578 323273 585662 323509
rect 585898 323273 585930 323509
rect 585310 296829 585930 323273
rect 585310 296593 585342 296829
rect 585578 296593 585662 296829
rect 585898 296593 585930 296829
rect 585310 296509 585930 296593
rect 585310 296273 585342 296509
rect 585578 296273 585662 296509
rect 585898 296273 585930 296509
rect 585310 269829 585930 296273
rect 585310 269593 585342 269829
rect 585578 269593 585662 269829
rect 585898 269593 585930 269829
rect 585310 269509 585930 269593
rect 585310 269273 585342 269509
rect 585578 269273 585662 269509
rect 585898 269273 585930 269509
rect 585310 242829 585930 269273
rect 585310 242593 585342 242829
rect 585578 242593 585662 242829
rect 585898 242593 585930 242829
rect 585310 242509 585930 242593
rect 585310 242273 585342 242509
rect 585578 242273 585662 242509
rect 585898 242273 585930 242509
rect 585310 215829 585930 242273
rect 585310 215593 585342 215829
rect 585578 215593 585662 215829
rect 585898 215593 585930 215829
rect 585310 215509 585930 215593
rect 585310 215273 585342 215509
rect 585578 215273 585662 215509
rect 585898 215273 585930 215509
rect 585310 188829 585930 215273
rect 585310 188593 585342 188829
rect 585578 188593 585662 188829
rect 585898 188593 585930 188829
rect 585310 188509 585930 188593
rect 585310 188273 585342 188509
rect 585578 188273 585662 188509
rect 585898 188273 585930 188509
rect 585310 161829 585930 188273
rect 585310 161593 585342 161829
rect 585578 161593 585662 161829
rect 585898 161593 585930 161829
rect 585310 161509 585930 161593
rect 585310 161273 585342 161509
rect 585578 161273 585662 161509
rect 585898 161273 585930 161509
rect 585310 134829 585930 161273
rect 585310 134593 585342 134829
rect 585578 134593 585662 134829
rect 585898 134593 585930 134829
rect 585310 134509 585930 134593
rect 585310 134273 585342 134509
rect 585578 134273 585662 134509
rect 585898 134273 585930 134509
rect 585310 107829 585930 134273
rect 585310 107593 585342 107829
rect 585578 107593 585662 107829
rect 585898 107593 585930 107829
rect 585310 107509 585930 107593
rect 585310 107273 585342 107509
rect 585578 107273 585662 107509
rect 585898 107273 585930 107509
rect 585310 80829 585930 107273
rect 585310 80593 585342 80829
rect 585578 80593 585662 80829
rect 585898 80593 585930 80829
rect 585310 80509 585930 80593
rect 585310 80273 585342 80509
rect 585578 80273 585662 80509
rect 585898 80273 585930 80509
rect 585310 53829 585930 80273
rect 585310 53593 585342 53829
rect 585578 53593 585662 53829
rect 585898 53593 585930 53829
rect 585310 53509 585930 53593
rect 585310 53273 585342 53509
rect 585578 53273 585662 53509
rect 585898 53273 585930 53509
rect 585310 26829 585930 53273
rect 585310 26593 585342 26829
rect 585578 26593 585662 26829
rect 585898 26593 585930 26829
rect 585310 26509 585930 26593
rect 585310 26273 585342 26509
rect 585578 26273 585662 26509
rect 585898 26273 585930 26509
rect 585310 -346 585930 26273
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 698454 586890 705242
rect 586270 698218 586302 698454
rect 586538 698218 586622 698454
rect 586858 698218 586890 698454
rect 586270 698134 586890 698218
rect 586270 697898 586302 698134
rect 586538 697898 586622 698134
rect 586858 697898 586890 698134
rect 586270 671454 586890 697898
rect 586270 671218 586302 671454
rect 586538 671218 586622 671454
rect 586858 671218 586890 671454
rect 586270 671134 586890 671218
rect 586270 670898 586302 671134
rect 586538 670898 586622 671134
rect 586858 670898 586890 671134
rect 586270 644454 586890 670898
rect 586270 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 586890 644454
rect 586270 644134 586890 644218
rect 586270 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 586890 644134
rect 586270 617454 586890 643898
rect 586270 617218 586302 617454
rect 586538 617218 586622 617454
rect 586858 617218 586890 617454
rect 586270 617134 586890 617218
rect 586270 616898 586302 617134
rect 586538 616898 586622 617134
rect 586858 616898 586890 617134
rect 586270 590454 586890 616898
rect 586270 590218 586302 590454
rect 586538 590218 586622 590454
rect 586858 590218 586890 590454
rect 586270 590134 586890 590218
rect 586270 589898 586302 590134
rect 586538 589898 586622 590134
rect 586858 589898 586890 590134
rect 586270 563454 586890 589898
rect 586270 563218 586302 563454
rect 586538 563218 586622 563454
rect 586858 563218 586890 563454
rect 586270 563134 586890 563218
rect 586270 562898 586302 563134
rect 586538 562898 586622 563134
rect 586858 562898 586890 563134
rect 586270 536454 586890 562898
rect 586270 536218 586302 536454
rect 586538 536218 586622 536454
rect 586858 536218 586890 536454
rect 586270 536134 586890 536218
rect 586270 535898 586302 536134
rect 586538 535898 586622 536134
rect 586858 535898 586890 536134
rect 586270 509454 586890 535898
rect 586270 509218 586302 509454
rect 586538 509218 586622 509454
rect 586858 509218 586890 509454
rect 586270 509134 586890 509218
rect 586270 508898 586302 509134
rect 586538 508898 586622 509134
rect 586858 508898 586890 509134
rect 586270 482454 586890 508898
rect 586270 482218 586302 482454
rect 586538 482218 586622 482454
rect 586858 482218 586890 482454
rect 586270 482134 586890 482218
rect 586270 481898 586302 482134
rect 586538 481898 586622 482134
rect 586858 481898 586890 482134
rect 586270 455454 586890 481898
rect 586270 455218 586302 455454
rect 586538 455218 586622 455454
rect 586858 455218 586890 455454
rect 586270 455134 586890 455218
rect 586270 454898 586302 455134
rect 586538 454898 586622 455134
rect 586858 454898 586890 455134
rect 586270 428454 586890 454898
rect 586270 428218 586302 428454
rect 586538 428218 586622 428454
rect 586858 428218 586890 428454
rect 586270 428134 586890 428218
rect 586270 427898 586302 428134
rect 586538 427898 586622 428134
rect 586858 427898 586890 428134
rect 586270 401454 586890 427898
rect 586270 401218 586302 401454
rect 586538 401218 586622 401454
rect 586858 401218 586890 401454
rect 586270 401134 586890 401218
rect 586270 400898 586302 401134
rect 586538 400898 586622 401134
rect 586858 400898 586890 401134
rect 586270 374454 586890 400898
rect 586270 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 586890 374454
rect 586270 374134 586890 374218
rect 586270 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 586890 374134
rect 586270 347454 586890 373898
rect 586270 347218 586302 347454
rect 586538 347218 586622 347454
rect 586858 347218 586890 347454
rect 586270 347134 586890 347218
rect 586270 346898 586302 347134
rect 586538 346898 586622 347134
rect 586858 346898 586890 347134
rect 586270 320454 586890 346898
rect 586270 320218 586302 320454
rect 586538 320218 586622 320454
rect 586858 320218 586890 320454
rect 586270 320134 586890 320218
rect 586270 319898 586302 320134
rect 586538 319898 586622 320134
rect 586858 319898 586890 320134
rect 586270 293454 586890 319898
rect 586270 293218 586302 293454
rect 586538 293218 586622 293454
rect 586858 293218 586890 293454
rect 586270 293134 586890 293218
rect 586270 292898 586302 293134
rect 586538 292898 586622 293134
rect 586858 292898 586890 293134
rect 586270 266454 586890 292898
rect 586270 266218 586302 266454
rect 586538 266218 586622 266454
rect 586858 266218 586890 266454
rect 586270 266134 586890 266218
rect 586270 265898 586302 266134
rect 586538 265898 586622 266134
rect 586858 265898 586890 266134
rect 586270 239454 586890 265898
rect 586270 239218 586302 239454
rect 586538 239218 586622 239454
rect 586858 239218 586890 239454
rect 586270 239134 586890 239218
rect 586270 238898 586302 239134
rect 586538 238898 586622 239134
rect 586858 238898 586890 239134
rect 586270 212454 586890 238898
rect 586270 212218 586302 212454
rect 586538 212218 586622 212454
rect 586858 212218 586890 212454
rect 586270 212134 586890 212218
rect 586270 211898 586302 212134
rect 586538 211898 586622 212134
rect 586858 211898 586890 212134
rect 586270 185454 586890 211898
rect 586270 185218 586302 185454
rect 586538 185218 586622 185454
rect 586858 185218 586890 185454
rect 586270 185134 586890 185218
rect 586270 184898 586302 185134
rect 586538 184898 586622 185134
rect 586858 184898 586890 185134
rect 586270 158454 586890 184898
rect 586270 158218 586302 158454
rect 586538 158218 586622 158454
rect 586858 158218 586890 158454
rect 586270 158134 586890 158218
rect 586270 157898 586302 158134
rect 586538 157898 586622 158134
rect 586858 157898 586890 158134
rect 586270 131454 586890 157898
rect 586270 131218 586302 131454
rect 586538 131218 586622 131454
rect 586858 131218 586890 131454
rect 586270 131134 586890 131218
rect 586270 130898 586302 131134
rect 586538 130898 586622 131134
rect 586858 130898 586890 131134
rect 586270 104454 586890 130898
rect 586270 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 586890 104454
rect 586270 104134 586890 104218
rect 586270 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 586890 104134
rect 586270 77454 586890 103898
rect 586270 77218 586302 77454
rect 586538 77218 586622 77454
rect 586858 77218 586890 77454
rect 586270 77134 586890 77218
rect 586270 76898 586302 77134
rect 586538 76898 586622 77134
rect 586858 76898 586890 77134
rect 586270 50454 586890 76898
rect 586270 50218 586302 50454
rect 586538 50218 586622 50454
rect 586858 50218 586890 50454
rect 586270 50134 586890 50218
rect 586270 49898 586302 50134
rect 586538 49898 586622 50134
rect 586858 49898 586890 50134
rect 586270 23454 586890 49898
rect 586270 23218 586302 23454
rect 586538 23218 586622 23454
rect 586858 23218 586890 23454
rect 586270 23134 586890 23218
rect 586270 22898 586302 23134
rect 586538 22898 586622 23134
rect 586858 22898 586890 23134
rect 586270 -1306 586890 22898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 -2266 587850 706202
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 -3226 588810 707162
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 -4186 589770 708122
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 -5146 590730 709082
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 -6106 591690 710042
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 -7066 592650 711002
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect 38026 705562 38262 705798
rect 38346 705562 38582 705798
rect 38026 705242 38262 705478
rect 38346 705242 38582 705478
rect -2934 698218 -2698 698454
rect -2614 698218 -2378 698454
rect -2934 697898 -2698 698134
rect -2614 697898 -2378 698134
rect -2934 671218 -2698 671454
rect -2614 671218 -2378 671454
rect -2934 670898 -2698 671134
rect -2614 670898 -2378 671134
rect -2934 644218 -2698 644454
rect -2614 644218 -2378 644454
rect -2934 643898 -2698 644134
rect -2614 643898 -2378 644134
rect -2934 617218 -2698 617454
rect -2614 617218 -2378 617454
rect -2934 616898 -2698 617134
rect -2614 616898 -2378 617134
rect -2934 590218 -2698 590454
rect -2614 590218 -2378 590454
rect -2934 589898 -2698 590134
rect -2614 589898 -2378 590134
rect -2934 563218 -2698 563454
rect -2614 563218 -2378 563454
rect -2934 562898 -2698 563134
rect -2614 562898 -2378 563134
rect -2934 536218 -2698 536454
rect -2614 536218 -2378 536454
rect -2934 535898 -2698 536134
rect -2614 535898 -2378 536134
rect -2934 509218 -2698 509454
rect -2614 509218 -2378 509454
rect -2934 508898 -2698 509134
rect -2614 508898 -2378 509134
rect -2934 482218 -2698 482454
rect -2614 482218 -2378 482454
rect -2934 481898 -2698 482134
rect -2614 481898 -2378 482134
rect -2934 455218 -2698 455454
rect -2614 455218 -2378 455454
rect -2934 454898 -2698 455134
rect -2614 454898 -2378 455134
rect -2934 428218 -2698 428454
rect -2614 428218 -2378 428454
rect -2934 427898 -2698 428134
rect -2614 427898 -2378 428134
rect -2934 401218 -2698 401454
rect -2614 401218 -2378 401454
rect -2934 400898 -2698 401134
rect -2614 400898 -2378 401134
rect -2934 374218 -2698 374454
rect -2614 374218 -2378 374454
rect -2934 373898 -2698 374134
rect -2614 373898 -2378 374134
rect -2934 347218 -2698 347454
rect -2614 347218 -2378 347454
rect -2934 346898 -2698 347134
rect -2614 346898 -2378 347134
rect -2934 320218 -2698 320454
rect -2614 320218 -2378 320454
rect -2934 319898 -2698 320134
rect -2614 319898 -2378 320134
rect -2934 293218 -2698 293454
rect -2614 293218 -2378 293454
rect -2934 292898 -2698 293134
rect -2614 292898 -2378 293134
rect -2934 266218 -2698 266454
rect -2614 266218 -2378 266454
rect -2934 265898 -2698 266134
rect -2614 265898 -2378 266134
rect -2934 239218 -2698 239454
rect -2614 239218 -2378 239454
rect -2934 238898 -2698 239134
rect -2614 238898 -2378 239134
rect -2934 212218 -2698 212454
rect -2614 212218 -2378 212454
rect -2934 211898 -2698 212134
rect -2614 211898 -2378 212134
rect -2934 185218 -2698 185454
rect -2614 185218 -2378 185454
rect -2934 184898 -2698 185134
rect -2614 184898 -2378 185134
rect -2934 158218 -2698 158454
rect -2614 158218 -2378 158454
rect -2934 157898 -2698 158134
rect -2614 157898 -2378 158134
rect -2934 131218 -2698 131454
rect -2614 131218 -2378 131454
rect -2934 130898 -2698 131134
rect -2614 130898 -2378 131134
rect -2934 104218 -2698 104454
rect -2614 104218 -2378 104454
rect -2934 103898 -2698 104134
rect -2614 103898 -2378 104134
rect -2934 77218 -2698 77454
rect -2614 77218 -2378 77454
rect -2934 76898 -2698 77134
rect -2614 76898 -2378 77134
rect -2934 50218 -2698 50454
rect -2614 50218 -2378 50454
rect -2934 49898 -2698 50134
rect -2614 49898 -2378 50134
rect -2934 23218 -2698 23454
rect -2614 23218 -2378 23454
rect -2934 22898 -2698 23134
rect -2614 22898 -2378 23134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 701593 -1738 701829
rect -1654 701593 -1418 701829
rect -1974 701273 -1738 701509
rect -1654 701273 -1418 701509
rect 38026 698218 38262 698454
rect 38346 698218 38582 698454
rect 38026 697898 38262 698134
rect 38346 697898 38582 698134
rect -1974 674593 -1738 674829
rect -1654 674593 -1418 674829
rect -1974 674273 -1738 674509
rect -1654 674273 -1418 674509
rect -1974 647593 -1738 647829
rect -1654 647593 -1418 647829
rect -1974 647273 -1738 647509
rect -1654 647273 -1418 647509
rect -1974 620593 -1738 620829
rect -1654 620593 -1418 620829
rect -1974 620273 -1738 620509
rect -1654 620273 -1418 620509
rect -1974 593593 -1738 593829
rect -1654 593593 -1418 593829
rect -1974 593273 -1738 593509
rect -1654 593273 -1418 593509
rect -1974 566593 -1738 566829
rect -1654 566593 -1418 566829
rect -1974 566273 -1738 566509
rect -1654 566273 -1418 566509
rect -1974 539593 -1738 539829
rect -1654 539593 -1418 539829
rect -1974 539273 -1738 539509
rect -1654 539273 -1418 539509
rect -1974 512593 -1738 512829
rect -1654 512593 -1418 512829
rect -1974 512273 -1738 512509
rect -1654 512273 -1418 512509
rect -1974 485593 -1738 485829
rect -1654 485593 -1418 485829
rect -1974 485273 -1738 485509
rect -1654 485273 -1418 485509
rect -1974 458593 -1738 458829
rect -1654 458593 -1418 458829
rect -1974 458273 -1738 458509
rect -1654 458273 -1418 458509
rect -1974 431593 -1738 431829
rect -1654 431593 -1418 431829
rect -1974 431273 -1738 431509
rect -1654 431273 -1418 431509
rect -1974 404593 -1738 404829
rect -1654 404593 -1418 404829
rect -1974 404273 -1738 404509
rect -1654 404273 -1418 404509
rect -1974 377593 -1738 377829
rect -1654 377593 -1418 377829
rect -1974 377273 -1738 377509
rect -1654 377273 -1418 377509
rect -1974 350593 -1738 350829
rect -1654 350593 -1418 350829
rect -1974 350273 -1738 350509
rect -1654 350273 -1418 350509
rect -1974 323593 -1738 323829
rect -1654 323593 -1418 323829
rect -1974 323273 -1738 323509
rect -1654 323273 -1418 323509
rect -1974 296593 -1738 296829
rect -1654 296593 -1418 296829
rect -1974 296273 -1738 296509
rect -1654 296273 -1418 296509
rect -1974 269593 -1738 269829
rect -1654 269593 -1418 269829
rect -1974 269273 -1738 269509
rect -1654 269273 -1418 269509
rect -1974 242593 -1738 242829
rect -1654 242593 -1418 242829
rect -1974 242273 -1738 242509
rect -1654 242273 -1418 242509
rect -1974 215593 -1738 215829
rect -1654 215593 -1418 215829
rect -1974 215273 -1738 215509
rect -1654 215273 -1418 215509
rect -1974 188593 -1738 188829
rect -1654 188593 -1418 188829
rect -1974 188273 -1738 188509
rect -1654 188273 -1418 188509
rect -1974 161593 -1738 161829
rect -1654 161593 -1418 161829
rect -1974 161273 -1738 161509
rect -1654 161273 -1418 161509
rect -1974 134593 -1738 134829
rect -1654 134593 -1418 134829
rect -1974 134273 -1738 134509
rect -1654 134273 -1418 134509
rect -1974 107593 -1738 107829
rect -1654 107593 -1418 107829
rect -1974 107273 -1738 107509
rect -1654 107273 -1418 107509
rect -1974 80593 -1738 80829
rect -1654 80593 -1418 80829
rect -1974 80273 -1738 80509
rect -1654 80273 -1418 80509
rect -1974 53593 -1738 53829
rect -1654 53593 -1418 53829
rect -1974 53273 -1738 53509
rect -1654 53273 -1418 53509
rect 38026 671218 38262 671454
rect 38346 671218 38582 671454
rect 38026 670898 38262 671134
rect 38346 670898 38582 671134
rect 38026 644218 38262 644454
rect 38346 644218 38582 644454
rect 38026 643898 38262 644134
rect 38346 643898 38582 644134
rect 38026 617218 38262 617454
rect 38346 617218 38582 617454
rect 38026 616898 38262 617134
rect 38346 616898 38582 617134
rect -1974 26593 -1738 26829
rect -1654 26593 -1418 26829
rect -1974 26273 -1738 26509
rect -1654 26273 -1418 26509
rect 38026 590218 38262 590454
rect 38346 590218 38582 590454
rect 38026 589898 38262 590134
rect 38346 589898 38582 590134
rect 38026 563218 38262 563454
rect 38346 563218 38582 563454
rect 38026 562898 38262 563134
rect 38346 562898 38582 563134
rect 38026 536218 38262 536454
rect 38346 536218 38582 536454
rect 38026 535898 38262 536134
rect 38346 535898 38582 536134
rect 38026 509218 38262 509454
rect 38346 509218 38582 509454
rect 38026 508898 38262 509134
rect 38346 508898 38582 509134
rect 38026 482218 38262 482454
rect 38346 482218 38582 482454
rect 38026 481898 38262 482134
rect 38346 481898 38582 482134
rect 38026 455218 38262 455454
rect 38346 455218 38582 455454
rect 38026 454898 38262 455134
rect 38346 454898 38582 455134
rect 38026 428218 38262 428454
rect 38346 428218 38582 428454
rect 38026 427898 38262 428134
rect 38346 427898 38582 428134
rect 38026 401218 38262 401454
rect 38346 401218 38582 401454
rect 38026 400898 38262 401134
rect 38346 400898 38582 401134
rect 38026 374218 38262 374454
rect 38346 374218 38582 374454
rect 38026 373898 38262 374134
rect 38346 373898 38582 374134
rect 38026 347218 38262 347454
rect 38346 347218 38582 347454
rect 38026 346898 38262 347134
rect 38346 346898 38582 347134
rect 38026 320218 38262 320454
rect 38346 320218 38582 320454
rect 38026 319898 38262 320134
rect 38346 319898 38582 320134
rect 38026 293218 38262 293454
rect 38346 293218 38582 293454
rect 38026 292898 38262 293134
rect 38346 292898 38582 293134
rect 38026 266218 38262 266454
rect 38346 266218 38582 266454
rect 38026 265898 38262 266134
rect 38346 265898 38582 266134
rect 38026 239218 38262 239454
rect 38346 239218 38582 239454
rect 38026 238898 38262 239134
rect 38346 238898 38582 239134
rect 38026 212218 38262 212454
rect 38346 212218 38582 212454
rect 38026 211898 38262 212134
rect 38346 211898 38582 212134
rect 38026 185218 38262 185454
rect 38346 185218 38582 185454
rect 38026 184898 38262 185134
rect 38346 184898 38582 185134
rect 38026 158218 38262 158454
rect 38346 158218 38582 158454
rect 38026 157898 38262 158134
rect 38346 157898 38582 158134
rect 38026 131218 38262 131454
rect 38346 131218 38582 131454
rect 38026 130898 38262 131134
rect 38346 130898 38582 131134
rect 38026 104218 38262 104454
rect 38346 104218 38582 104454
rect 38026 103898 38262 104134
rect 38346 103898 38582 104134
rect 38026 77218 38262 77454
rect 38346 77218 38582 77454
rect 38026 76898 38262 77134
rect 38346 76898 38582 77134
rect 38026 50218 38262 50454
rect 38346 50218 38582 50454
rect 38026 49898 38262 50134
rect 38346 49898 38582 50134
rect 41526 704602 41762 704838
rect 41846 704602 42082 704838
rect 41526 704282 41762 704518
rect 41846 704282 42082 704518
rect 41526 701593 41762 701829
rect 41846 701593 42082 701829
rect 41526 701273 41762 701509
rect 41846 701273 42082 701509
rect 41526 674593 41762 674829
rect 41846 674593 42082 674829
rect 41526 674273 41762 674509
rect 41846 674273 42082 674509
rect 41526 647593 41762 647829
rect 41846 647593 42082 647829
rect 41526 647273 41762 647509
rect 41846 647273 42082 647509
rect 41526 620593 41762 620829
rect 41846 620593 42082 620829
rect 41526 620273 41762 620509
rect 41846 620273 42082 620509
rect 41526 593593 41762 593829
rect 41846 593593 42082 593829
rect 41526 593273 41762 593509
rect 41846 593273 42082 593509
rect 41526 566593 41762 566829
rect 41846 566593 42082 566829
rect 41526 566273 41762 566509
rect 41846 566273 42082 566509
rect 41526 539593 41762 539829
rect 41846 539593 42082 539829
rect 41526 539273 41762 539509
rect 41846 539273 42082 539509
rect 41526 512593 41762 512829
rect 41846 512593 42082 512829
rect 41526 512273 41762 512509
rect 41846 512273 42082 512509
rect 66026 705562 66262 705798
rect 66346 705562 66582 705798
rect 66026 705242 66262 705478
rect 66346 705242 66582 705478
rect 66026 698218 66262 698454
rect 66346 698218 66582 698454
rect 66026 697898 66262 698134
rect 66346 697898 66582 698134
rect 66026 671218 66262 671454
rect 66346 671218 66582 671454
rect 66026 670898 66262 671134
rect 66346 670898 66582 671134
rect 66026 644218 66262 644454
rect 66346 644218 66582 644454
rect 66026 643898 66262 644134
rect 66346 643898 66582 644134
rect 66026 617218 66262 617454
rect 66346 617218 66582 617454
rect 66026 616898 66262 617134
rect 66346 616898 66582 617134
rect 66026 590218 66262 590454
rect 66346 590218 66582 590454
rect 66026 589898 66262 590134
rect 66346 589898 66582 590134
rect 66026 563218 66262 563454
rect 66346 563218 66582 563454
rect 66026 562898 66262 563134
rect 66346 562898 66582 563134
rect 66026 536218 66262 536454
rect 66346 536218 66582 536454
rect 66026 535898 66262 536134
rect 66346 535898 66582 536134
rect 66026 509218 66262 509454
rect 66346 509218 66582 509454
rect 66026 508898 66262 509134
rect 66346 508898 66582 509134
rect 41526 485593 41762 485829
rect 41846 485593 42082 485829
rect 41526 485273 41762 485509
rect 41846 485273 42082 485509
rect 41526 458593 41762 458829
rect 41846 458593 42082 458829
rect 41526 458273 41762 458509
rect 41846 458273 42082 458509
rect 41526 431593 41762 431829
rect 41846 431593 42082 431829
rect 41526 431273 41762 431509
rect 41846 431273 42082 431509
rect 41526 404593 41762 404829
rect 41846 404593 42082 404829
rect 41526 404273 41762 404509
rect 41846 404273 42082 404509
rect 41526 377593 41762 377829
rect 41846 377593 42082 377829
rect 41526 377273 41762 377509
rect 41846 377273 42082 377509
rect 41526 350593 41762 350829
rect 41846 350593 42082 350829
rect 41526 350273 41762 350509
rect 41846 350273 42082 350509
rect 41526 323593 41762 323829
rect 41846 323593 42082 323829
rect 41526 323273 41762 323509
rect 41846 323273 42082 323509
rect 41526 296593 41762 296829
rect 41846 296593 42082 296829
rect 41526 296273 41762 296509
rect 41846 296273 42082 296509
rect 41526 269593 41762 269829
rect 41846 269593 42082 269829
rect 41526 269273 41762 269509
rect 41846 269273 42082 269509
rect 41526 242593 41762 242829
rect 41846 242593 42082 242829
rect 41526 242273 41762 242509
rect 41846 242273 42082 242509
rect 41526 215593 41762 215829
rect 41846 215593 42082 215829
rect 41526 215273 41762 215509
rect 41846 215273 42082 215509
rect 41526 188593 41762 188829
rect 41846 188593 42082 188829
rect 41526 188273 41762 188509
rect 41846 188273 42082 188509
rect 41526 161593 41762 161829
rect 41846 161593 42082 161829
rect 41526 161273 41762 161509
rect 41846 161273 42082 161509
rect 41526 134593 41762 134829
rect 41846 134593 42082 134829
rect 41526 134273 41762 134509
rect 41846 134273 42082 134509
rect 41526 107593 41762 107829
rect 41846 107593 42082 107829
rect 41526 107273 41762 107509
rect 41846 107273 42082 107509
rect 41526 80593 41762 80829
rect 41846 80593 42082 80829
rect 41526 80273 41762 80509
rect 41846 80273 42082 80509
rect 41526 53593 41762 53829
rect 41846 53593 42082 53829
rect 41526 53273 41762 53509
rect 41846 53273 42082 53509
rect 22460 26593 22696 26829
rect 22460 26273 22696 26509
rect 33408 26593 33644 26829
rect 33408 26273 33644 26509
rect 27934 23218 28170 23454
rect 27934 22898 28170 23134
rect 38882 23218 39118 23454
rect 38882 22898 39118 23134
rect 44356 26593 44592 26829
rect 44356 26273 44592 26509
rect 66026 482218 66262 482454
rect 66346 482218 66582 482454
rect 66026 481898 66262 482134
rect 66346 481898 66582 482134
rect 49830 23218 50066 23454
rect 49830 22898 50066 23134
rect 66026 455218 66262 455454
rect 66346 455218 66582 455454
rect 66026 454898 66262 455134
rect 66346 454898 66582 455134
rect 66026 428218 66262 428454
rect 66346 428218 66582 428454
rect 66026 427898 66262 428134
rect 66346 427898 66582 428134
rect 66026 401218 66262 401454
rect 66346 401218 66582 401454
rect 66026 400898 66262 401134
rect 66346 400898 66582 401134
rect 66026 374218 66262 374454
rect 66346 374218 66582 374454
rect 66026 373898 66262 374134
rect 66346 373898 66582 374134
rect 66026 347218 66262 347454
rect 66346 347218 66582 347454
rect 66026 346898 66262 347134
rect 66346 346898 66582 347134
rect 66026 320218 66262 320454
rect 66346 320218 66582 320454
rect 66026 319898 66262 320134
rect 66346 319898 66582 320134
rect 66026 293218 66262 293454
rect 66346 293218 66582 293454
rect 66026 292898 66262 293134
rect 66346 292898 66582 293134
rect 66026 266218 66262 266454
rect 66346 266218 66582 266454
rect 66026 265898 66262 266134
rect 66346 265898 66582 266134
rect 66026 239218 66262 239454
rect 66346 239218 66582 239454
rect 66026 238898 66262 239134
rect 66346 238898 66582 239134
rect 66026 212218 66262 212454
rect 66346 212218 66582 212454
rect 66026 211898 66262 212134
rect 66346 211898 66582 212134
rect 66026 185218 66262 185454
rect 66346 185218 66582 185454
rect 66026 184898 66262 185134
rect 66346 184898 66582 185134
rect 66026 158218 66262 158454
rect 66346 158218 66582 158454
rect 66026 157898 66262 158134
rect 66346 157898 66582 158134
rect 66026 131218 66262 131454
rect 66346 131218 66582 131454
rect 66026 130898 66262 131134
rect 66346 130898 66582 131134
rect 66026 104218 66262 104454
rect 66346 104218 66582 104454
rect 66026 103898 66262 104134
rect 66346 103898 66582 104134
rect 66026 77218 66262 77454
rect 66346 77218 66582 77454
rect 66026 76898 66262 77134
rect 66346 76898 66582 77134
rect 66026 50218 66262 50454
rect 66346 50218 66582 50454
rect 66026 49898 66262 50134
rect 66346 49898 66582 50134
rect 55304 26593 55540 26829
rect 55304 26273 55540 26509
rect 60778 23218 61014 23454
rect 60778 22898 61014 23134
rect 66026 23218 66262 23454
rect 66346 23218 66582 23454
rect 66026 22898 66262 23134
rect 66346 22898 66582 23134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 66026 -1542 66262 -1306
rect 66346 -1542 66582 -1306
rect 66026 -1862 66262 -1626
rect 66346 -1862 66582 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 69526 704602 69762 704838
rect 69846 704602 70082 704838
rect 69526 704282 69762 704518
rect 69846 704282 70082 704518
rect 69526 701593 69762 701829
rect 69846 701593 70082 701829
rect 69526 701273 69762 701509
rect 69846 701273 70082 701509
rect 69526 674593 69762 674829
rect 69846 674593 70082 674829
rect 69526 674273 69762 674509
rect 69846 674273 70082 674509
rect 69526 647593 69762 647829
rect 69846 647593 70082 647829
rect 69526 647273 69762 647509
rect 69846 647273 70082 647509
rect 69526 620593 69762 620829
rect 69846 620593 70082 620829
rect 69526 620273 69762 620509
rect 69846 620273 70082 620509
rect 69526 593593 69762 593829
rect 69846 593593 70082 593829
rect 69526 593273 69762 593509
rect 69846 593273 70082 593509
rect 69526 566593 69762 566829
rect 69846 566593 70082 566829
rect 69526 566273 69762 566509
rect 69846 566273 70082 566509
rect 69526 539593 69762 539829
rect 69846 539593 70082 539829
rect 69526 539273 69762 539509
rect 69846 539273 70082 539509
rect 69526 512593 69762 512829
rect 69846 512593 70082 512829
rect 69526 512273 69762 512509
rect 69846 512273 70082 512509
rect 69526 485593 69762 485829
rect 69846 485593 70082 485829
rect 69526 485273 69762 485509
rect 69846 485273 70082 485509
rect 69526 458593 69762 458829
rect 69846 458593 70082 458829
rect 69526 458273 69762 458509
rect 69846 458273 70082 458509
rect 69526 431593 69762 431829
rect 69846 431593 70082 431829
rect 69526 431273 69762 431509
rect 69846 431273 70082 431509
rect 69526 404593 69762 404829
rect 69846 404593 70082 404829
rect 69526 404273 69762 404509
rect 69846 404273 70082 404509
rect 69526 377593 69762 377829
rect 69846 377593 70082 377829
rect 69526 377273 69762 377509
rect 69846 377273 70082 377509
rect 69526 350593 69762 350829
rect 69846 350593 70082 350829
rect 69526 350273 69762 350509
rect 69846 350273 70082 350509
rect 69526 323593 69762 323829
rect 69846 323593 70082 323829
rect 69526 323273 69762 323509
rect 69846 323273 70082 323509
rect 69526 296593 69762 296829
rect 69846 296593 70082 296829
rect 69526 296273 69762 296509
rect 69846 296273 70082 296509
rect 69526 269593 69762 269829
rect 69846 269593 70082 269829
rect 69526 269273 69762 269509
rect 69846 269273 70082 269509
rect 69526 242593 69762 242829
rect 69846 242593 70082 242829
rect 69526 242273 69762 242509
rect 69846 242273 70082 242509
rect 69526 215593 69762 215829
rect 69846 215593 70082 215829
rect 69526 215273 69762 215509
rect 69846 215273 70082 215509
rect 69526 188593 69762 188829
rect 69846 188593 70082 188829
rect 69526 188273 69762 188509
rect 69846 188273 70082 188509
rect 69526 161593 69762 161829
rect 69846 161593 70082 161829
rect 69526 161273 69762 161509
rect 69846 161273 70082 161509
rect 69526 134593 69762 134829
rect 69846 134593 70082 134829
rect 69526 134273 69762 134509
rect 69846 134273 70082 134509
rect 69526 107593 69762 107829
rect 69846 107593 70082 107829
rect 69526 107273 69762 107509
rect 69846 107273 70082 107509
rect 69526 80593 69762 80829
rect 69846 80593 70082 80829
rect 69526 80273 69762 80509
rect 69846 80273 70082 80509
rect 69526 53593 69762 53829
rect 69846 53593 70082 53829
rect 69526 53273 69762 53509
rect 69846 53273 70082 53509
rect 94026 705562 94262 705798
rect 94346 705562 94582 705798
rect 94026 705242 94262 705478
rect 94346 705242 94582 705478
rect 94026 698218 94262 698454
rect 94346 698218 94582 698454
rect 94026 697898 94262 698134
rect 94346 697898 94582 698134
rect 94026 671218 94262 671454
rect 94346 671218 94582 671454
rect 94026 670898 94262 671134
rect 94346 670898 94582 671134
rect 94026 644218 94262 644454
rect 94346 644218 94582 644454
rect 94026 643898 94262 644134
rect 94346 643898 94582 644134
rect 94026 617218 94262 617454
rect 94346 617218 94582 617454
rect 94026 616898 94262 617134
rect 94346 616898 94582 617134
rect 94026 590218 94262 590454
rect 94346 590218 94582 590454
rect 94026 589898 94262 590134
rect 94346 589898 94582 590134
rect 94026 563218 94262 563454
rect 94346 563218 94582 563454
rect 94026 562898 94262 563134
rect 94346 562898 94582 563134
rect 94026 536218 94262 536454
rect 94346 536218 94582 536454
rect 94026 535898 94262 536134
rect 94346 535898 94582 536134
rect 94026 509218 94262 509454
rect 94346 509218 94582 509454
rect 94026 508898 94262 509134
rect 94346 508898 94582 509134
rect 94026 482218 94262 482454
rect 94346 482218 94582 482454
rect 94026 481898 94262 482134
rect 94346 481898 94582 482134
rect 94026 455218 94262 455454
rect 94346 455218 94582 455454
rect 94026 454898 94262 455134
rect 94346 454898 94582 455134
rect 94026 428218 94262 428454
rect 94346 428218 94582 428454
rect 94026 427898 94262 428134
rect 94346 427898 94582 428134
rect 94026 401218 94262 401454
rect 94346 401218 94582 401454
rect 94026 400898 94262 401134
rect 94346 400898 94582 401134
rect 94026 374218 94262 374454
rect 94346 374218 94582 374454
rect 94026 373898 94262 374134
rect 94346 373898 94582 374134
rect 94026 347218 94262 347454
rect 94346 347218 94582 347454
rect 94026 346898 94262 347134
rect 94346 346898 94582 347134
rect 94026 320218 94262 320454
rect 94346 320218 94582 320454
rect 94026 319898 94262 320134
rect 94346 319898 94582 320134
rect 94026 293218 94262 293454
rect 94346 293218 94582 293454
rect 94026 292898 94262 293134
rect 94346 292898 94582 293134
rect 94026 266218 94262 266454
rect 94346 266218 94582 266454
rect 94026 265898 94262 266134
rect 94346 265898 94582 266134
rect 94026 239218 94262 239454
rect 94346 239218 94582 239454
rect 94026 238898 94262 239134
rect 94346 238898 94582 239134
rect 94026 212218 94262 212454
rect 94346 212218 94582 212454
rect 94026 211898 94262 212134
rect 94346 211898 94582 212134
rect 94026 185218 94262 185454
rect 94346 185218 94582 185454
rect 94026 184898 94262 185134
rect 94346 184898 94582 185134
rect 94026 158218 94262 158454
rect 94346 158218 94582 158454
rect 94026 157898 94262 158134
rect 94346 157898 94582 158134
rect 94026 131218 94262 131454
rect 94346 131218 94582 131454
rect 94026 130898 94262 131134
rect 94346 130898 94582 131134
rect 94026 104218 94262 104454
rect 94346 104218 94582 104454
rect 94026 103898 94262 104134
rect 94346 103898 94582 104134
rect 94026 77218 94262 77454
rect 94346 77218 94582 77454
rect 94026 76898 94262 77134
rect 94346 76898 94582 77134
rect 94026 50218 94262 50454
rect 94346 50218 94582 50454
rect 94026 49898 94262 50134
rect 94346 49898 94582 50134
rect 97526 704602 97762 704838
rect 97846 704602 98082 704838
rect 97526 704282 97762 704518
rect 97846 704282 98082 704518
rect 97526 701593 97762 701829
rect 97846 701593 98082 701829
rect 97526 701273 97762 701509
rect 97846 701273 98082 701509
rect 97526 674593 97762 674829
rect 97846 674593 98082 674829
rect 97526 674273 97762 674509
rect 97846 674273 98082 674509
rect 97526 647593 97762 647829
rect 97846 647593 98082 647829
rect 97526 647273 97762 647509
rect 97846 647273 98082 647509
rect 97526 620593 97762 620829
rect 97846 620593 98082 620829
rect 97526 620273 97762 620509
rect 97846 620273 98082 620509
rect 97526 593593 97762 593829
rect 97846 593593 98082 593829
rect 97526 593273 97762 593509
rect 97846 593273 98082 593509
rect 97526 566593 97762 566829
rect 97846 566593 98082 566829
rect 97526 566273 97762 566509
rect 97846 566273 98082 566509
rect 97526 539593 97762 539829
rect 97846 539593 98082 539829
rect 97526 539273 97762 539509
rect 97846 539273 98082 539509
rect 97526 512593 97762 512829
rect 97846 512593 98082 512829
rect 97526 512273 97762 512509
rect 97846 512273 98082 512509
rect 97526 485593 97762 485829
rect 97846 485593 98082 485829
rect 97526 485273 97762 485509
rect 97846 485273 98082 485509
rect 97526 458593 97762 458829
rect 97846 458593 98082 458829
rect 97526 458273 97762 458509
rect 97846 458273 98082 458509
rect 97526 431593 97762 431829
rect 97846 431593 98082 431829
rect 97526 431273 97762 431509
rect 97846 431273 98082 431509
rect 97526 404593 97762 404829
rect 97846 404593 98082 404829
rect 97526 404273 97762 404509
rect 97846 404273 98082 404509
rect 97526 377593 97762 377829
rect 97846 377593 98082 377829
rect 97526 377273 97762 377509
rect 97846 377273 98082 377509
rect 97526 350593 97762 350829
rect 97846 350593 98082 350829
rect 97526 350273 97762 350509
rect 97846 350273 98082 350509
rect 97526 323593 97762 323829
rect 97846 323593 98082 323829
rect 97526 323273 97762 323509
rect 97846 323273 98082 323509
rect 97526 296593 97762 296829
rect 97846 296593 98082 296829
rect 97526 296273 97762 296509
rect 97846 296273 98082 296509
rect 97526 269593 97762 269829
rect 97846 269593 98082 269829
rect 97526 269273 97762 269509
rect 97846 269273 98082 269509
rect 97526 242593 97762 242829
rect 97846 242593 98082 242829
rect 97526 242273 97762 242509
rect 97846 242273 98082 242509
rect 97526 215593 97762 215829
rect 97846 215593 98082 215829
rect 97526 215273 97762 215509
rect 97846 215273 98082 215509
rect 97526 188593 97762 188829
rect 97846 188593 98082 188829
rect 97526 188273 97762 188509
rect 97846 188273 98082 188509
rect 97526 161593 97762 161829
rect 97846 161593 98082 161829
rect 97526 161273 97762 161509
rect 97846 161273 98082 161509
rect 97526 134593 97762 134829
rect 97846 134593 98082 134829
rect 97526 134273 97762 134509
rect 97846 134273 98082 134509
rect 97526 107593 97762 107829
rect 97846 107593 98082 107829
rect 97526 107273 97762 107509
rect 97846 107273 98082 107509
rect 97526 80593 97762 80829
rect 97846 80593 98082 80829
rect 97526 80273 97762 80509
rect 97846 80273 98082 80509
rect 97526 53593 97762 53829
rect 97846 53593 98082 53829
rect 97526 53273 97762 53509
rect 97846 53273 98082 53509
rect 122026 705562 122262 705798
rect 122346 705562 122582 705798
rect 122026 705242 122262 705478
rect 122346 705242 122582 705478
rect 122026 698218 122262 698454
rect 122346 698218 122582 698454
rect 122026 697898 122262 698134
rect 122346 697898 122582 698134
rect 122026 671218 122262 671454
rect 122346 671218 122582 671454
rect 122026 670898 122262 671134
rect 122346 670898 122582 671134
rect 122026 644218 122262 644454
rect 122346 644218 122582 644454
rect 122026 643898 122262 644134
rect 122346 643898 122582 644134
rect 122026 617218 122262 617454
rect 122346 617218 122582 617454
rect 122026 616898 122262 617134
rect 122346 616898 122582 617134
rect 122026 590218 122262 590454
rect 122346 590218 122582 590454
rect 122026 589898 122262 590134
rect 122346 589898 122582 590134
rect 122026 563218 122262 563454
rect 122346 563218 122582 563454
rect 122026 562898 122262 563134
rect 122346 562898 122582 563134
rect 122026 536218 122262 536454
rect 122346 536218 122582 536454
rect 122026 535898 122262 536134
rect 122346 535898 122582 536134
rect 122026 509218 122262 509454
rect 122346 509218 122582 509454
rect 122026 508898 122262 509134
rect 122346 508898 122582 509134
rect 122026 482218 122262 482454
rect 122346 482218 122582 482454
rect 122026 481898 122262 482134
rect 122346 481898 122582 482134
rect 122026 455218 122262 455454
rect 122346 455218 122582 455454
rect 122026 454898 122262 455134
rect 122346 454898 122582 455134
rect 122026 428218 122262 428454
rect 122346 428218 122582 428454
rect 122026 427898 122262 428134
rect 122346 427898 122582 428134
rect 122026 401218 122262 401454
rect 122346 401218 122582 401454
rect 122026 400898 122262 401134
rect 122346 400898 122582 401134
rect 122026 374218 122262 374454
rect 122346 374218 122582 374454
rect 122026 373898 122262 374134
rect 122346 373898 122582 374134
rect 122026 347218 122262 347454
rect 122346 347218 122582 347454
rect 122026 346898 122262 347134
rect 122346 346898 122582 347134
rect 122026 320218 122262 320454
rect 122346 320218 122582 320454
rect 122026 319898 122262 320134
rect 122346 319898 122582 320134
rect 122026 293218 122262 293454
rect 122346 293218 122582 293454
rect 122026 292898 122262 293134
rect 122346 292898 122582 293134
rect 122026 266218 122262 266454
rect 122346 266218 122582 266454
rect 122026 265898 122262 266134
rect 122346 265898 122582 266134
rect 122026 239218 122262 239454
rect 122346 239218 122582 239454
rect 122026 238898 122262 239134
rect 122346 238898 122582 239134
rect 122026 212218 122262 212454
rect 122346 212218 122582 212454
rect 122026 211898 122262 212134
rect 122346 211898 122582 212134
rect 122026 185218 122262 185454
rect 122346 185218 122582 185454
rect 122026 184898 122262 185134
rect 122346 184898 122582 185134
rect 122026 158218 122262 158454
rect 122346 158218 122582 158454
rect 122026 157898 122262 158134
rect 122346 157898 122582 158134
rect 122026 131218 122262 131454
rect 122346 131218 122582 131454
rect 122026 130898 122262 131134
rect 122346 130898 122582 131134
rect 122026 104218 122262 104454
rect 122346 104218 122582 104454
rect 122026 103898 122262 104134
rect 122346 103898 122582 104134
rect 122026 77218 122262 77454
rect 122346 77218 122582 77454
rect 122026 76898 122262 77134
rect 122346 76898 122582 77134
rect 122026 50218 122262 50454
rect 122346 50218 122582 50454
rect 122026 49898 122262 50134
rect 122346 49898 122582 50134
rect 125526 704602 125762 704838
rect 125846 704602 126082 704838
rect 125526 704282 125762 704518
rect 125846 704282 126082 704518
rect 125526 701593 125762 701829
rect 125846 701593 126082 701829
rect 125526 701273 125762 701509
rect 125846 701273 126082 701509
rect 125526 674593 125762 674829
rect 125846 674593 126082 674829
rect 125526 674273 125762 674509
rect 125846 674273 126082 674509
rect 125526 647593 125762 647829
rect 125846 647593 126082 647829
rect 125526 647273 125762 647509
rect 125846 647273 126082 647509
rect 125526 620593 125762 620829
rect 125846 620593 126082 620829
rect 125526 620273 125762 620509
rect 125846 620273 126082 620509
rect 125526 593593 125762 593829
rect 125846 593593 126082 593829
rect 125526 593273 125762 593509
rect 125846 593273 126082 593509
rect 125526 566593 125762 566829
rect 125846 566593 126082 566829
rect 125526 566273 125762 566509
rect 125846 566273 126082 566509
rect 125526 539593 125762 539829
rect 125846 539593 126082 539829
rect 125526 539273 125762 539509
rect 125846 539273 126082 539509
rect 125526 512593 125762 512829
rect 125846 512593 126082 512829
rect 125526 512273 125762 512509
rect 125846 512273 126082 512509
rect 125526 485593 125762 485829
rect 125846 485593 126082 485829
rect 125526 485273 125762 485509
rect 125846 485273 126082 485509
rect 125526 458593 125762 458829
rect 125846 458593 126082 458829
rect 125526 458273 125762 458509
rect 125846 458273 126082 458509
rect 125526 431593 125762 431829
rect 125846 431593 126082 431829
rect 125526 431273 125762 431509
rect 125846 431273 126082 431509
rect 125526 404593 125762 404829
rect 125846 404593 126082 404829
rect 125526 404273 125762 404509
rect 125846 404273 126082 404509
rect 125526 377593 125762 377829
rect 125846 377593 126082 377829
rect 125526 377273 125762 377509
rect 125846 377273 126082 377509
rect 125526 350593 125762 350829
rect 125846 350593 126082 350829
rect 125526 350273 125762 350509
rect 125846 350273 126082 350509
rect 125526 323593 125762 323829
rect 125846 323593 126082 323829
rect 125526 323273 125762 323509
rect 125846 323273 126082 323509
rect 125526 296593 125762 296829
rect 125846 296593 126082 296829
rect 125526 296273 125762 296509
rect 125846 296273 126082 296509
rect 125526 269593 125762 269829
rect 125846 269593 126082 269829
rect 125526 269273 125762 269509
rect 125846 269273 126082 269509
rect 125526 242593 125762 242829
rect 125846 242593 126082 242829
rect 125526 242273 125762 242509
rect 125846 242273 126082 242509
rect 125526 215593 125762 215829
rect 125846 215593 126082 215829
rect 125526 215273 125762 215509
rect 125846 215273 126082 215509
rect 125526 188593 125762 188829
rect 125846 188593 126082 188829
rect 125526 188273 125762 188509
rect 125846 188273 126082 188509
rect 125526 161593 125762 161829
rect 125846 161593 126082 161829
rect 125526 161273 125762 161509
rect 125846 161273 126082 161509
rect 125526 134593 125762 134829
rect 125846 134593 126082 134829
rect 125526 134273 125762 134509
rect 125846 134273 126082 134509
rect 125526 107593 125762 107829
rect 125846 107593 126082 107829
rect 125526 107273 125762 107509
rect 125846 107273 126082 107509
rect 125526 80593 125762 80829
rect 125846 80593 126082 80829
rect 125526 80273 125762 80509
rect 125846 80273 126082 80509
rect 125526 53593 125762 53829
rect 125846 53593 126082 53829
rect 125526 53273 125762 53509
rect 125846 53273 126082 53509
rect 150026 705562 150262 705798
rect 150346 705562 150582 705798
rect 150026 705242 150262 705478
rect 150346 705242 150582 705478
rect 150026 698218 150262 698454
rect 150346 698218 150582 698454
rect 150026 697898 150262 698134
rect 150346 697898 150582 698134
rect 150026 671218 150262 671454
rect 150346 671218 150582 671454
rect 150026 670898 150262 671134
rect 150346 670898 150582 671134
rect 150026 644218 150262 644454
rect 150346 644218 150582 644454
rect 150026 643898 150262 644134
rect 150346 643898 150582 644134
rect 150026 617218 150262 617454
rect 150346 617218 150582 617454
rect 150026 616898 150262 617134
rect 150346 616898 150582 617134
rect 150026 590218 150262 590454
rect 150346 590218 150582 590454
rect 150026 589898 150262 590134
rect 150346 589898 150582 590134
rect 150026 563218 150262 563454
rect 150346 563218 150582 563454
rect 150026 562898 150262 563134
rect 150346 562898 150582 563134
rect 150026 536218 150262 536454
rect 150346 536218 150582 536454
rect 150026 535898 150262 536134
rect 150346 535898 150582 536134
rect 150026 509218 150262 509454
rect 150346 509218 150582 509454
rect 150026 508898 150262 509134
rect 150346 508898 150582 509134
rect 150026 482218 150262 482454
rect 150346 482218 150582 482454
rect 150026 481898 150262 482134
rect 150346 481898 150582 482134
rect 150026 455218 150262 455454
rect 150346 455218 150582 455454
rect 150026 454898 150262 455134
rect 150346 454898 150582 455134
rect 150026 428218 150262 428454
rect 150346 428218 150582 428454
rect 150026 427898 150262 428134
rect 150346 427898 150582 428134
rect 150026 401218 150262 401454
rect 150346 401218 150582 401454
rect 150026 400898 150262 401134
rect 150346 400898 150582 401134
rect 150026 374218 150262 374454
rect 150346 374218 150582 374454
rect 150026 373898 150262 374134
rect 150346 373898 150582 374134
rect 150026 347218 150262 347454
rect 150346 347218 150582 347454
rect 150026 346898 150262 347134
rect 150346 346898 150582 347134
rect 150026 320218 150262 320454
rect 150346 320218 150582 320454
rect 150026 319898 150262 320134
rect 150346 319898 150582 320134
rect 150026 293218 150262 293454
rect 150346 293218 150582 293454
rect 150026 292898 150262 293134
rect 150346 292898 150582 293134
rect 150026 266218 150262 266454
rect 150346 266218 150582 266454
rect 150026 265898 150262 266134
rect 150346 265898 150582 266134
rect 150026 239218 150262 239454
rect 150346 239218 150582 239454
rect 150026 238898 150262 239134
rect 150346 238898 150582 239134
rect 150026 212218 150262 212454
rect 150346 212218 150582 212454
rect 150026 211898 150262 212134
rect 150346 211898 150582 212134
rect 150026 185218 150262 185454
rect 150346 185218 150582 185454
rect 150026 184898 150262 185134
rect 150346 184898 150582 185134
rect 150026 158218 150262 158454
rect 150346 158218 150582 158454
rect 150026 157898 150262 158134
rect 150346 157898 150582 158134
rect 150026 131218 150262 131454
rect 150346 131218 150582 131454
rect 150026 130898 150262 131134
rect 150346 130898 150582 131134
rect 150026 104218 150262 104454
rect 150346 104218 150582 104454
rect 150026 103898 150262 104134
rect 150346 103898 150582 104134
rect 150026 77218 150262 77454
rect 150346 77218 150582 77454
rect 150026 76898 150262 77134
rect 150346 76898 150582 77134
rect 150026 50218 150262 50454
rect 150346 50218 150582 50454
rect 150026 49898 150262 50134
rect 150346 49898 150582 50134
rect 153526 704602 153762 704838
rect 153846 704602 154082 704838
rect 153526 704282 153762 704518
rect 153846 704282 154082 704518
rect 153526 701593 153762 701829
rect 153846 701593 154082 701829
rect 153526 701273 153762 701509
rect 153846 701273 154082 701509
rect 178026 705562 178262 705798
rect 178346 705562 178582 705798
rect 178026 705242 178262 705478
rect 178346 705242 178582 705478
rect 153526 674593 153762 674829
rect 153846 674593 154082 674829
rect 153526 674273 153762 674509
rect 153846 674273 154082 674509
rect 153526 647593 153762 647829
rect 153846 647593 154082 647829
rect 153526 647273 153762 647509
rect 153846 647273 154082 647509
rect 153526 620593 153762 620829
rect 153846 620593 154082 620829
rect 153526 620273 153762 620509
rect 153846 620273 154082 620509
rect 153526 593593 153762 593829
rect 153846 593593 154082 593829
rect 153526 593273 153762 593509
rect 153846 593273 154082 593509
rect 153526 566593 153762 566829
rect 153846 566593 154082 566829
rect 153526 566273 153762 566509
rect 153846 566273 154082 566509
rect 153526 539593 153762 539829
rect 153846 539593 154082 539829
rect 153526 539273 153762 539509
rect 153846 539273 154082 539509
rect 153526 512593 153762 512829
rect 153846 512593 154082 512829
rect 153526 512273 153762 512509
rect 153846 512273 154082 512509
rect 153526 485593 153762 485829
rect 153846 485593 154082 485829
rect 153526 485273 153762 485509
rect 153846 485273 154082 485509
rect 153526 458593 153762 458829
rect 153846 458593 154082 458829
rect 153526 458273 153762 458509
rect 153846 458273 154082 458509
rect 153526 431593 153762 431829
rect 153846 431593 154082 431829
rect 153526 431273 153762 431509
rect 153846 431273 154082 431509
rect 153526 404593 153762 404829
rect 153846 404593 154082 404829
rect 153526 404273 153762 404509
rect 153846 404273 154082 404509
rect 153526 377593 153762 377829
rect 153846 377593 154082 377829
rect 153526 377273 153762 377509
rect 153846 377273 154082 377509
rect 153526 350593 153762 350829
rect 153846 350593 154082 350829
rect 153526 350273 153762 350509
rect 153846 350273 154082 350509
rect 153526 323593 153762 323829
rect 153846 323593 154082 323829
rect 153526 323273 153762 323509
rect 153846 323273 154082 323509
rect 153526 296593 153762 296829
rect 153846 296593 154082 296829
rect 153526 296273 153762 296509
rect 153846 296273 154082 296509
rect 153526 269593 153762 269829
rect 153846 269593 154082 269829
rect 153526 269273 153762 269509
rect 153846 269273 154082 269509
rect 153526 242593 153762 242829
rect 153846 242593 154082 242829
rect 153526 242273 153762 242509
rect 153846 242273 154082 242509
rect 153526 215593 153762 215829
rect 153846 215593 154082 215829
rect 153526 215273 153762 215509
rect 153846 215273 154082 215509
rect 153526 188593 153762 188829
rect 153846 188593 154082 188829
rect 153526 188273 153762 188509
rect 153846 188273 154082 188509
rect 153526 161593 153762 161829
rect 153846 161593 154082 161829
rect 153526 161273 153762 161509
rect 153846 161273 154082 161509
rect 153526 134593 153762 134829
rect 153846 134593 154082 134829
rect 153526 134273 153762 134509
rect 153846 134273 154082 134509
rect 153526 107593 153762 107829
rect 153846 107593 154082 107829
rect 153526 107273 153762 107509
rect 153846 107273 154082 107509
rect 153526 80593 153762 80829
rect 153846 80593 154082 80829
rect 153526 80273 153762 80509
rect 153846 80273 154082 80509
rect 153526 53593 153762 53829
rect 153846 53593 154082 53829
rect 153526 53273 153762 53509
rect 153846 53273 154082 53509
rect 69526 26593 69762 26829
rect 69846 26593 70082 26829
rect 69526 26273 69762 26509
rect 69846 26273 70082 26509
rect 75460 26593 75696 26829
rect 75460 26273 75696 26509
rect 76408 26593 76644 26829
rect 76408 26273 76644 26509
rect 77356 26593 77592 26829
rect 77356 26273 77592 26509
rect 78304 26593 78540 26829
rect 78304 26273 78540 26509
rect 84160 26593 84396 26829
rect 84160 26273 84396 26509
rect 88108 26593 88344 26829
rect 88108 26273 88344 26509
rect 92056 26593 92292 26829
rect 92056 26273 92292 26509
rect 96004 26593 96240 26829
rect 96004 26273 96240 26509
rect 104460 26593 104696 26829
rect 104460 26273 104696 26509
rect 105408 26593 105644 26829
rect 105408 26273 105644 26509
rect 106356 26593 106592 26829
rect 106356 26273 106592 26509
rect 107304 26593 107540 26829
rect 107304 26273 107540 26509
rect 113160 26593 113396 26829
rect 113160 26273 113396 26509
rect 117108 26593 117344 26829
rect 117108 26273 117344 26509
rect 121056 26593 121292 26829
rect 121056 26273 121292 26509
rect 125004 26593 125240 26829
rect 125004 26273 125240 26509
rect 133460 26593 133696 26829
rect 133460 26273 133696 26509
rect 134408 26593 134644 26829
rect 134408 26273 134644 26509
rect 135356 26593 135592 26829
rect 135356 26273 135592 26509
rect 136304 26593 136540 26829
rect 136304 26273 136540 26509
rect 142160 26593 142396 26829
rect 142160 26273 142396 26509
rect 146108 26593 146344 26829
rect 146108 26273 146344 26509
rect 150056 26593 150292 26829
rect 150056 26273 150292 26509
rect 154004 26593 154240 26829
rect 154004 26273 154240 26509
rect 162460 26593 162696 26829
rect 162460 26273 162696 26509
rect 163408 26593 163644 26829
rect 163408 26273 163644 26509
rect 164356 26593 164592 26829
rect 164356 26273 164592 26509
rect 165304 26593 165540 26829
rect 165304 26273 165540 26509
rect 75934 23218 76170 23454
rect 75934 22898 76170 23134
rect 76882 23218 77118 23454
rect 76882 22898 77118 23134
rect 77830 23218 78066 23454
rect 77830 22898 78066 23134
rect 86134 23218 86370 23454
rect 86134 22898 86370 23134
rect 90082 23218 90318 23454
rect 90082 22898 90318 23134
rect 94030 23218 94266 23454
rect 94030 22898 94266 23134
rect 104934 23218 105170 23454
rect 104934 22898 105170 23134
rect 105882 23218 106118 23454
rect 105882 22898 106118 23134
rect 106830 23218 107066 23454
rect 106830 22898 107066 23134
rect 115134 23218 115370 23454
rect 115134 22898 115370 23134
rect 119082 23218 119318 23454
rect 119082 22898 119318 23134
rect 123030 23218 123266 23454
rect 123030 22898 123266 23134
rect 133934 23218 134170 23454
rect 133934 22898 134170 23134
rect 134882 23218 135118 23454
rect 134882 22898 135118 23134
rect 135830 23218 136066 23454
rect 135830 22898 136066 23134
rect 144134 23218 144370 23454
rect 144134 22898 144370 23134
rect 148082 23218 148318 23454
rect 148082 22898 148318 23134
rect 152030 23218 152266 23454
rect 152030 22898 152266 23134
rect 162934 23218 163170 23454
rect 162934 22898 163170 23134
rect 163882 23218 164118 23454
rect 163882 22898 164118 23134
rect 164830 23218 165066 23454
rect 164830 22898 165066 23134
rect 178026 698218 178262 698454
rect 178346 698218 178582 698454
rect 178026 697898 178262 698134
rect 178346 697898 178582 698134
rect 178026 671218 178262 671454
rect 178346 671218 178582 671454
rect 178026 670898 178262 671134
rect 178346 670898 178582 671134
rect 178026 644218 178262 644454
rect 178346 644218 178582 644454
rect 178026 643898 178262 644134
rect 178346 643898 178582 644134
rect 178026 617218 178262 617454
rect 178346 617218 178582 617454
rect 178026 616898 178262 617134
rect 178346 616898 178582 617134
rect 178026 590218 178262 590454
rect 178346 590218 178582 590454
rect 178026 589898 178262 590134
rect 178346 589898 178582 590134
rect 178026 563218 178262 563454
rect 178346 563218 178582 563454
rect 178026 562898 178262 563134
rect 178346 562898 178582 563134
rect 178026 536218 178262 536454
rect 178346 536218 178582 536454
rect 178026 535898 178262 536134
rect 178346 535898 178582 536134
rect 178026 509218 178262 509454
rect 178346 509218 178582 509454
rect 178026 508898 178262 509134
rect 178346 508898 178582 509134
rect 178026 482218 178262 482454
rect 178346 482218 178582 482454
rect 178026 481898 178262 482134
rect 178346 481898 178582 482134
rect 178026 455218 178262 455454
rect 178346 455218 178582 455454
rect 178026 454898 178262 455134
rect 178346 454898 178582 455134
rect 178026 428218 178262 428454
rect 178346 428218 178582 428454
rect 178026 427898 178262 428134
rect 178346 427898 178582 428134
rect 178026 401218 178262 401454
rect 178346 401218 178582 401454
rect 178026 400898 178262 401134
rect 178346 400898 178582 401134
rect 178026 374218 178262 374454
rect 178346 374218 178582 374454
rect 178026 373898 178262 374134
rect 178346 373898 178582 374134
rect 178026 347218 178262 347454
rect 178346 347218 178582 347454
rect 178026 346898 178262 347134
rect 178346 346898 178582 347134
rect 178026 320218 178262 320454
rect 178346 320218 178582 320454
rect 178026 319898 178262 320134
rect 178346 319898 178582 320134
rect 178026 293218 178262 293454
rect 178346 293218 178582 293454
rect 178026 292898 178262 293134
rect 178346 292898 178582 293134
rect 178026 266218 178262 266454
rect 178346 266218 178582 266454
rect 178026 265898 178262 266134
rect 178346 265898 178582 266134
rect 178026 239218 178262 239454
rect 178346 239218 178582 239454
rect 178026 238898 178262 239134
rect 178346 238898 178582 239134
rect 178026 212218 178262 212454
rect 178346 212218 178582 212454
rect 178026 211898 178262 212134
rect 178346 211898 178582 212134
rect 178026 185218 178262 185454
rect 178346 185218 178582 185454
rect 178026 184898 178262 185134
rect 178346 184898 178582 185134
rect 178026 158218 178262 158454
rect 178346 158218 178582 158454
rect 178026 157898 178262 158134
rect 178346 157898 178582 158134
rect 178026 131218 178262 131454
rect 178346 131218 178582 131454
rect 178026 130898 178262 131134
rect 178346 130898 178582 131134
rect 178026 104218 178262 104454
rect 178346 104218 178582 104454
rect 178026 103898 178262 104134
rect 178346 103898 178582 104134
rect 178026 77218 178262 77454
rect 178346 77218 178582 77454
rect 178026 76898 178262 77134
rect 178346 76898 178582 77134
rect 178026 50218 178262 50454
rect 178346 50218 178582 50454
rect 178026 49898 178262 50134
rect 178346 49898 178582 50134
rect 181526 704602 181762 704838
rect 181846 704602 182082 704838
rect 181526 704282 181762 704518
rect 181846 704282 182082 704518
rect 181526 701593 181762 701829
rect 181846 701593 182082 701829
rect 181526 701273 181762 701509
rect 181846 701273 182082 701509
rect 181526 674593 181762 674829
rect 181846 674593 182082 674829
rect 181526 674273 181762 674509
rect 181846 674273 182082 674509
rect 181526 647593 181762 647829
rect 181846 647593 182082 647829
rect 181526 647273 181762 647509
rect 181846 647273 182082 647509
rect 181526 620593 181762 620829
rect 181846 620593 182082 620829
rect 181526 620273 181762 620509
rect 181846 620273 182082 620509
rect 181526 593593 181762 593829
rect 181846 593593 182082 593829
rect 181526 593273 181762 593509
rect 181846 593273 182082 593509
rect 181526 566593 181762 566829
rect 181846 566593 182082 566829
rect 181526 566273 181762 566509
rect 181846 566273 182082 566509
rect 181526 539593 181762 539829
rect 181846 539593 182082 539829
rect 181526 539273 181762 539509
rect 181846 539273 182082 539509
rect 181526 512593 181762 512829
rect 181846 512593 182082 512829
rect 181526 512273 181762 512509
rect 181846 512273 182082 512509
rect 181526 485593 181762 485829
rect 181846 485593 182082 485829
rect 181526 485273 181762 485509
rect 181846 485273 182082 485509
rect 181526 458593 181762 458829
rect 181846 458593 182082 458829
rect 181526 458273 181762 458509
rect 181846 458273 182082 458509
rect 181526 431593 181762 431829
rect 181846 431593 182082 431829
rect 181526 431273 181762 431509
rect 181846 431273 182082 431509
rect 181526 404593 181762 404829
rect 181846 404593 182082 404829
rect 181526 404273 181762 404509
rect 181846 404273 182082 404509
rect 181526 377593 181762 377829
rect 181846 377593 182082 377829
rect 181526 377273 181762 377509
rect 181846 377273 182082 377509
rect 181526 350593 181762 350829
rect 181846 350593 182082 350829
rect 181526 350273 181762 350509
rect 181846 350273 182082 350509
rect 181526 323593 181762 323829
rect 181846 323593 182082 323829
rect 181526 323273 181762 323509
rect 181846 323273 182082 323509
rect 181526 296593 181762 296829
rect 181846 296593 182082 296829
rect 181526 296273 181762 296509
rect 181846 296273 182082 296509
rect 181526 269593 181762 269829
rect 181846 269593 182082 269829
rect 181526 269273 181762 269509
rect 181846 269273 182082 269509
rect 181526 242593 181762 242829
rect 181846 242593 182082 242829
rect 181526 242273 181762 242509
rect 181846 242273 182082 242509
rect 181526 215593 181762 215829
rect 181846 215593 182082 215829
rect 181526 215273 181762 215509
rect 181846 215273 182082 215509
rect 181526 188593 181762 188829
rect 181846 188593 182082 188829
rect 181526 188273 181762 188509
rect 181846 188273 182082 188509
rect 181526 161593 181762 161829
rect 181846 161593 182082 161829
rect 181526 161273 181762 161509
rect 181846 161273 182082 161509
rect 181526 134593 181762 134829
rect 181846 134593 182082 134829
rect 181526 134273 181762 134509
rect 181846 134273 182082 134509
rect 181526 107593 181762 107829
rect 181846 107593 182082 107829
rect 181526 107273 181762 107509
rect 181846 107273 182082 107509
rect 181526 80593 181762 80829
rect 181846 80593 182082 80829
rect 181526 80273 181762 80509
rect 181846 80273 182082 80509
rect 206026 705562 206262 705798
rect 206346 705562 206582 705798
rect 206026 705242 206262 705478
rect 206346 705242 206582 705478
rect 206026 698218 206262 698454
rect 206346 698218 206582 698454
rect 206026 697898 206262 698134
rect 206346 697898 206582 698134
rect 206026 671218 206262 671454
rect 206346 671218 206582 671454
rect 206026 670898 206262 671134
rect 206346 670898 206582 671134
rect 206026 644218 206262 644454
rect 206346 644218 206582 644454
rect 206026 643898 206262 644134
rect 206346 643898 206582 644134
rect 206026 617218 206262 617454
rect 206346 617218 206582 617454
rect 206026 616898 206262 617134
rect 206346 616898 206582 617134
rect 206026 590218 206262 590454
rect 206346 590218 206582 590454
rect 206026 589898 206262 590134
rect 206346 589898 206582 590134
rect 206026 563218 206262 563454
rect 206346 563218 206582 563454
rect 206026 562898 206262 563134
rect 206346 562898 206582 563134
rect 206026 536218 206262 536454
rect 206346 536218 206582 536454
rect 206026 535898 206262 536134
rect 206346 535898 206582 536134
rect 206026 509218 206262 509454
rect 206346 509218 206582 509454
rect 206026 508898 206262 509134
rect 206346 508898 206582 509134
rect 206026 482218 206262 482454
rect 206346 482218 206582 482454
rect 206026 481898 206262 482134
rect 206346 481898 206582 482134
rect 206026 455218 206262 455454
rect 206346 455218 206582 455454
rect 206026 454898 206262 455134
rect 206346 454898 206582 455134
rect 206026 428218 206262 428454
rect 206346 428218 206582 428454
rect 206026 427898 206262 428134
rect 206346 427898 206582 428134
rect 206026 401218 206262 401454
rect 206346 401218 206582 401454
rect 206026 400898 206262 401134
rect 206346 400898 206582 401134
rect 206026 374218 206262 374454
rect 206346 374218 206582 374454
rect 206026 373898 206262 374134
rect 206346 373898 206582 374134
rect 206026 347218 206262 347454
rect 206346 347218 206582 347454
rect 206026 346898 206262 347134
rect 206346 346898 206582 347134
rect 206026 320218 206262 320454
rect 206346 320218 206582 320454
rect 206026 319898 206262 320134
rect 206346 319898 206582 320134
rect 206026 293218 206262 293454
rect 206346 293218 206582 293454
rect 206026 292898 206262 293134
rect 206346 292898 206582 293134
rect 206026 266218 206262 266454
rect 206346 266218 206582 266454
rect 206026 265898 206262 266134
rect 206346 265898 206582 266134
rect 206026 239218 206262 239454
rect 206346 239218 206582 239454
rect 206026 238898 206262 239134
rect 206346 238898 206582 239134
rect 206026 212218 206262 212454
rect 206346 212218 206582 212454
rect 206026 211898 206262 212134
rect 206346 211898 206582 212134
rect 206026 185218 206262 185454
rect 206346 185218 206582 185454
rect 206026 184898 206262 185134
rect 206346 184898 206582 185134
rect 206026 158218 206262 158454
rect 206346 158218 206582 158454
rect 206026 157898 206262 158134
rect 206346 157898 206582 158134
rect 206026 131218 206262 131454
rect 206346 131218 206582 131454
rect 206026 130898 206262 131134
rect 206346 130898 206582 131134
rect 206026 104218 206262 104454
rect 206346 104218 206582 104454
rect 206026 103898 206262 104134
rect 206346 103898 206582 104134
rect 206026 77218 206262 77454
rect 206346 77218 206582 77454
rect 206026 76898 206262 77134
rect 206346 76898 206582 77134
rect 209526 704602 209762 704838
rect 209846 704602 210082 704838
rect 209526 704282 209762 704518
rect 209846 704282 210082 704518
rect 209526 701593 209762 701829
rect 209846 701593 210082 701829
rect 209526 701273 209762 701509
rect 209846 701273 210082 701509
rect 209526 674593 209762 674829
rect 209846 674593 210082 674829
rect 209526 674273 209762 674509
rect 209846 674273 210082 674509
rect 209526 647593 209762 647829
rect 209846 647593 210082 647829
rect 209526 647273 209762 647509
rect 209846 647273 210082 647509
rect 209526 620593 209762 620829
rect 209846 620593 210082 620829
rect 209526 620273 209762 620509
rect 209846 620273 210082 620509
rect 209526 593593 209762 593829
rect 209846 593593 210082 593829
rect 209526 593273 209762 593509
rect 209846 593273 210082 593509
rect 209526 566593 209762 566829
rect 209846 566593 210082 566829
rect 209526 566273 209762 566509
rect 209846 566273 210082 566509
rect 209526 539593 209762 539829
rect 209846 539593 210082 539829
rect 209526 539273 209762 539509
rect 209846 539273 210082 539509
rect 209526 512593 209762 512829
rect 209846 512593 210082 512829
rect 209526 512273 209762 512509
rect 209846 512273 210082 512509
rect 209526 485593 209762 485829
rect 209846 485593 210082 485829
rect 209526 485273 209762 485509
rect 209846 485273 210082 485509
rect 209526 458593 209762 458829
rect 209846 458593 210082 458829
rect 209526 458273 209762 458509
rect 209846 458273 210082 458509
rect 209526 431593 209762 431829
rect 209846 431593 210082 431829
rect 209526 431273 209762 431509
rect 209846 431273 210082 431509
rect 209526 404593 209762 404829
rect 209846 404593 210082 404829
rect 209526 404273 209762 404509
rect 209846 404273 210082 404509
rect 209526 377593 209762 377829
rect 209846 377593 210082 377829
rect 209526 377273 209762 377509
rect 209846 377273 210082 377509
rect 209526 350593 209762 350829
rect 209846 350593 210082 350829
rect 209526 350273 209762 350509
rect 209846 350273 210082 350509
rect 209526 323593 209762 323829
rect 209846 323593 210082 323829
rect 209526 323273 209762 323509
rect 209846 323273 210082 323509
rect 209526 296593 209762 296829
rect 209846 296593 210082 296829
rect 209526 296273 209762 296509
rect 209846 296273 210082 296509
rect 209526 269593 209762 269829
rect 209846 269593 210082 269829
rect 209526 269273 209762 269509
rect 209846 269273 210082 269509
rect 209526 242593 209762 242829
rect 209846 242593 210082 242829
rect 209526 242273 209762 242509
rect 209846 242273 210082 242509
rect 209526 215593 209762 215829
rect 209846 215593 210082 215829
rect 209526 215273 209762 215509
rect 209846 215273 210082 215509
rect 209526 188593 209762 188829
rect 209846 188593 210082 188829
rect 209526 188273 209762 188509
rect 209846 188273 210082 188509
rect 209526 161593 209762 161829
rect 209846 161593 210082 161829
rect 209526 161273 209762 161509
rect 209846 161273 210082 161509
rect 209526 134593 209762 134829
rect 209846 134593 210082 134829
rect 209526 134273 209762 134509
rect 209846 134273 210082 134509
rect 209526 107593 209762 107829
rect 209846 107593 210082 107829
rect 209526 107273 209762 107509
rect 209846 107273 210082 107509
rect 209526 80593 209762 80829
rect 209846 80593 210082 80829
rect 209526 80273 209762 80509
rect 209846 80273 210082 80509
rect 234026 705562 234262 705798
rect 234346 705562 234582 705798
rect 234026 705242 234262 705478
rect 234346 705242 234582 705478
rect 234026 698218 234262 698454
rect 234346 698218 234582 698454
rect 234026 697898 234262 698134
rect 234346 697898 234582 698134
rect 234026 671218 234262 671454
rect 234346 671218 234582 671454
rect 234026 670898 234262 671134
rect 234346 670898 234582 671134
rect 234026 644218 234262 644454
rect 234346 644218 234582 644454
rect 234026 643898 234262 644134
rect 234346 643898 234582 644134
rect 234026 617218 234262 617454
rect 234346 617218 234582 617454
rect 234026 616898 234262 617134
rect 234346 616898 234582 617134
rect 234026 590218 234262 590454
rect 234346 590218 234582 590454
rect 234026 589898 234262 590134
rect 234346 589898 234582 590134
rect 234026 563218 234262 563454
rect 234346 563218 234582 563454
rect 234026 562898 234262 563134
rect 234346 562898 234582 563134
rect 234026 536218 234262 536454
rect 234346 536218 234582 536454
rect 234026 535898 234262 536134
rect 234346 535898 234582 536134
rect 234026 509218 234262 509454
rect 234346 509218 234582 509454
rect 234026 508898 234262 509134
rect 234346 508898 234582 509134
rect 234026 482218 234262 482454
rect 234346 482218 234582 482454
rect 234026 481898 234262 482134
rect 234346 481898 234582 482134
rect 234026 455218 234262 455454
rect 234346 455218 234582 455454
rect 234026 454898 234262 455134
rect 234346 454898 234582 455134
rect 234026 428218 234262 428454
rect 234346 428218 234582 428454
rect 234026 427898 234262 428134
rect 234346 427898 234582 428134
rect 234026 401218 234262 401454
rect 234346 401218 234582 401454
rect 234026 400898 234262 401134
rect 234346 400898 234582 401134
rect 234026 374218 234262 374454
rect 234346 374218 234582 374454
rect 234026 373898 234262 374134
rect 234346 373898 234582 374134
rect 234026 347218 234262 347454
rect 234346 347218 234582 347454
rect 234026 346898 234262 347134
rect 234346 346898 234582 347134
rect 234026 320218 234262 320454
rect 234346 320218 234582 320454
rect 234026 319898 234262 320134
rect 234346 319898 234582 320134
rect 234026 293218 234262 293454
rect 234346 293218 234582 293454
rect 234026 292898 234262 293134
rect 234346 292898 234582 293134
rect 234026 266218 234262 266454
rect 234346 266218 234582 266454
rect 234026 265898 234262 266134
rect 234346 265898 234582 266134
rect 234026 239218 234262 239454
rect 234346 239218 234582 239454
rect 234026 238898 234262 239134
rect 234346 238898 234582 239134
rect 234026 212218 234262 212454
rect 234346 212218 234582 212454
rect 234026 211898 234262 212134
rect 234346 211898 234582 212134
rect 234026 185218 234262 185454
rect 234346 185218 234582 185454
rect 234026 184898 234262 185134
rect 234346 184898 234582 185134
rect 234026 158218 234262 158454
rect 234346 158218 234582 158454
rect 234026 157898 234262 158134
rect 234346 157898 234582 158134
rect 234026 131218 234262 131454
rect 234346 131218 234582 131454
rect 234026 130898 234262 131134
rect 234346 130898 234582 131134
rect 234026 104218 234262 104454
rect 234346 104218 234582 104454
rect 234026 103898 234262 104134
rect 234346 103898 234582 104134
rect 234026 77218 234262 77454
rect 234346 77218 234582 77454
rect 234026 76898 234262 77134
rect 234346 76898 234582 77134
rect 237526 704602 237762 704838
rect 237846 704602 238082 704838
rect 237526 704282 237762 704518
rect 237846 704282 238082 704518
rect 237526 701593 237762 701829
rect 237846 701593 238082 701829
rect 237526 701273 237762 701509
rect 237846 701273 238082 701509
rect 237526 674593 237762 674829
rect 237846 674593 238082 674829
rect 237526 674273 237762 674509
rect 237846 674273 238082 674509
rect 237526 647593 237762 647829
rect 237846 647593 238082 647829
rect 237526 647273 237762 647509
rect 237846 647273 238082 647509
rect 237526 620593 237762 620829
rect 237846 620593 238082 620829
rect 237526 620273 237762 620509
rect 237846 620273 238082 620509
rect 237526 593593 237762 593829
rect 237846 593593 238082 593829
rect 237526 593273 237762 593509
rect 237846 593273 238082 593509
rect 237526 566593 237762 566829
rect 237846 566593 238082 566829
rect 237526 566273 237762 566509
rect 237846 566273 238082 566509
rect 237526 539593 237762 539829
rect 237846 539593 238082 539829
rect 237526 539273 237762 539509
rect 237846 539273 238082 539509
rect 237526 512593 237762 512829
rect 237846 512593 238082 512829
rect 237526 512273 237762 512509
rect 237846 512273 238082 512509
rect 237526 485593 237762 485829
rect 237846 485593 238082 485829
rect 237526 485273 237762 485509
rect 237846 485273 238082 485509
rect 237526 458593 237762 458829
rect 237846 458593 238082 458829
rect 237526 458273 237762 458509
rect 237846 458273 238082 458509
rect 237526 431593 237762 431829
rect 237846 431593 238082 431829
rect 237526 431273 237762 431509
rect 237846 431273 238082 431509
rect 237526 404593 237762 404829
rect 237846 404593 238082 404829
rect 237526 404273 237762 404509
rect 237846 404273 238082 404509
rect 237526 377593 237762 377829
rect 237846 377593 238082 377829
rect 237526 377273 237762 377509
rect 237846 377273 238082 377509
rect 237526 350593 237762 350829
rect 237846 350593 238082 350829
rect 237526 350273 237762 350509
rect 237846 350273 238082 350509
rect 237526 323593 237762 323829
rect 237846 323593 238082 323829
rect 237526 323273 237762 323509
rect 237846 323273 238082 323509
rect 237526 296593 237762 296829
rect 237846 296593 238082 296829
rect 237526 296273 237762 296509
rect 237846 296273 238082 296509
rect 237526 269593 237762 269829
rect 237846 269593 238082 269829
rect 237526 269273 237762 269509
rect 237846 269273 238082 269509
rect 237526 242593 237762 242829
rect 237846 242593 238082 242829
rect 237526 242273 237762 242509
rect 237846 242273 238082 242509
rect 237526 215593 237762 215829
rect 237846 215593 238082 215829
rect 237526 215273 237762 215509
rect 237846 215273 238082 215509
rect 237526 188593 237762 188829
rect 237846 188593 238082 188829
rect 237526 188273 237762 188509
rect 237846 188273 238082 188509
rect 237526 161593 237762 161829
rect 237846 161593 238082 161829
rect 237526 161273 237762 161509
rect 237846 161273 238082 161509
rect 237526 134593 237762 134829
rect 237846 134593 238082 134829
rect 237526 134273 237762 134509
rect 237846 134273 238082 134509
rect 237526 107593 237762 107829
rect 237846 107593 238082 107829
rect 237526 107273 237762 107509
rect 237846 107273 238082 107509
rect 237526 80593 237762 80829
rect 237846 80593 238082 80829
rect 237526 80273 237762 80509
rect 237846 80273 238082 80509
rect 262026 705562 262262 705798
rect 262346 705562 262582 705798
rect 262026 705242 262262 705478
rect 262346 705242 262582 705478
rect 262026 698218 262262 698454
rect 262346 698218 262582 698454
rect 262026 697898 262262 698134
rect 262346 697898 262582 698134
rect 262026 671218 262262 671454
rect 262346 671218 262582 671454
rect 262026 670898 262262 671134
rect 262346 670898 262582 671134
rect 262026 644218 262262 644454
rect 262346 644218 262582 644454
rect 262026 643898 262262 644134
rect 262346 643898 262582 644134
rect 262026 617218 262262 617454
rect 262346 617218 262582 617454
rect 262026 616898 262262 617134
rect 262346 616898 262582 617134
rect 262026 590218 262262 590454
rect 262346 590218 262582 590454
rect 262026 589898 262262 590134
rect 262346 589898 262582 590134
rect 262026 563218 262262 563454
rect 262346 563218 262582 563454
rect 262026 562898 262262 563134
rect 262346 562898 262582 563134
rect 262026 536218 262262 536454
rect 262346 536218 262582 536454
rect 262026 535898 262262 536134
rect 262346 535898 262582 536134
rect 262026 509218 262262 509454
rect 262346 509218 262582 509454
rect 262026 508898 262262 509134
rect 262346 508898 262582 509134
rect 262026 482218 262262 482454
rect 262346 482218 262582 482454
rect 262026 481898 262262 482134
rect 262346 481898 262582 482134
rect 262026 455218 262262 455454
rect 262346 455218 262582 455454
rect 262026 454898 262262 455134
rect 262346 454898 262582 455134
rect 262026 428218 262262 428454
rect 262346 428218 262582 428454
rect 262026 427898 262262 428134
rect 262346 427898 262582 428134
rect 262026 401218 262262 401454
rect 262346 401218 262582 401454
rect 262026 400898 262262 401134
rect 262346 400898 262582 401134
rect 262026 374218 262262 374454
rect 262346 374218 262582 374454
rect 262026 373898 262262 374134
rect 262346 373898 262582 374134
rect 262026 347218 262262 347454
rect 262346 347218 262582 347454
rect 262026 346898 262262 347134
rect 262346 346898 262582 347134
rect 262026 320218 262262 320454
rect 262346 320218 262582 320454
rect 262026 319898 262262 320134
rect 262346 319898 262582 320134
rect 262026 293218 262262 293454
rect 262346 293218 262582 293454
rect 262026 292898 262262 293134
rect 262346 292898 262582 293134
rect 262026 266218 262262 266454
rect 262346 266218 262582 266454
rect 262026 265898 262262 266134
rect 262346 265898 262582 266134
rect 262026 239218 262262 239454
rect 262346 239218 262582 239454
rect 262026 238898 262262 239134
rect 262346 238898 262582 239134
rect 262026 212218 262262 212454
rect 262346 212218 262582 212454
rect 262026 211898 262262 212134
rect 262346 211898 262582 212134
rect 262026 185218 262262 185454
rect 262346 185218 262582 185454
rect 262026 184898 262262 185134
rect 262346 184898 262582 185134
rect 262026 158218 262262 158454
rect 262346 158218 262582 158454
rect 262026 157898 262262 158134
rect 262346 157898 262582 158134
rect 262026 131218 262262 131454
rect 262346 131218 262582 131454
rect 262026 130898 262262 131134
rect 262346 130898 262582 131134
rect 262026 104218 262262 104454
rect 262346 104218 262582 104454
rect 262026 103898 262262 104134
rect 262346 103898 262582 104134
rect 262026 77218 262262 77454
rect 262346 77218 262582 77454
rect 262026 76898 262262 77134
rect 262346 76898 262582 77134
rect 265526 704602 265762 704838
rect 265846 704602 266082 704838
rect 265526 704282 265762 704518
rect 265846 704282 266082 704518
rect 265526 701593 265762 701829
rect 265846 701593 266082 701829
rect 265526 701273 265762 701509
rect 265846 701273 266082 701509
rect 265526 674593 265762 674829
rect 265846 674593 266082 674829
rect 265526 674273 265762 674509
rect 265846 674273 266082 674509
rect 265526 647593 265762 647829
rect 265846 647593 266082 647829
rect 265526 647273 265762 647509
rect 265846 647273 266082 647509
rect 265526 620593 265762 620829
rect 265846 620593 266082 620829
rect 265526 620273 265762 620509
rect 265846 620273 266082 620509
rect 265526 593593 265762 593829
rect 265846 593593 266082 593829
rect 265526 593273 265762 593509
rect 265846 593273 266082 593509
rect 265526 566593 265762 566829
rect 265846 566593 266082 566829
rect 265526 566273 265762 566509
rect 265846 566273 266082 566509
rect 265526 539593 265762 539829
rect 265846 539593 266082 539829
rect 265526 539273 265762 539509
rect 265846 539273 266082 539509
rect 265526 512593 265762 512829
rect 265846 512593 266082 512829
rect 265526 512273 265762 512509
rect 265846 512273 266082 512509
rect 265526 485593 265762 485829
rect 265846 485593 266082 485829
rect 265526 485273 265762 485509
rect 265846 485273 266082 485509
rect 265526 458593 265762 458829
rect 265846 458593 266082 458829
rect 265526 458273 265762 458509
rect 265846 458273 266082 458509
rect 265526 431593 265762 431829
rect 265846 431593 266082 431829
rect 265526 431273 265762 431509
rect 265846 431273 266082 431509
rect 265526 404593 265762 404829
rect 265846 404593 266082 404829
rect 265526 404273 265762 404509
rect 265846 404273 266082 404509
rect 265526 377593 265762 377829
rect 265846 377593 266082 377829
rect 265526 377273 265762 377509
rect 265846 377273 266082 377509
rect 265526 350593 265762 350829
rect 265846 350593 266082 350829
rect 265526 350273 265762 350509
rect 265846 350273 266082 350509
rect 265526 323593 265762 323829
rect 265846 323593 266082 323829
rect 265526 323273 265762 323509
rect 265846 323273 266082 323509
rect 265526 296593 265762 296829
rect 265846 296593 266082 296829
rect 265526 296273 265762 296509
rect 265846 296273 266082 296509
rect 265526 269593 265762 269829
rect 265846 269593 266082 269829
rect 265526 269273 265762 269509
rect 265846 269273 266082 269509
rect 265526 242593 265762 242829
rect 265846 242593 266082 242829
rect 265526 242273 265762 242509
rect 265846 242273 266082 242509
rect 265526 215593 265762 215829
rect 265846 215593 266082 215829
rect 265526 215273 265762 215509
rect 265846 215273 266082 215509
rect 265526 188593 265762 188829
rect 265846 188593 266082 188829
rect 265526 188273 265762 188509
rect 265846 188273 266082 188509
rect 265526 161593 265762 161829
rect 265846 161593 266082 161829
rect 265526 161273 265762 161509
rect 265846 161273 266082 161509
rect 265526 134593 265762 134829
rect 265846 134593 266082 134829
rect 265526 134273 265762 134509
rect 265846 134273 266082 134509
rect 265526 107593 265762 107829
rect 265846 107593 266082 107829
rect 265526 107273 265762 107509
rect 265846 107273 266082 107509
rect 265526 80593 265762 80829
rect 265846 80593 266082 80829
rect 265526 80273 265762 80509
rect 265846 80273 266082 80509
rect 290026 705562 290262 705798
rect 290346 705562 290582 705798
rect 290026 705242 290262 705478
rect 290346 705242 290582 705478
rect 290026 698218 290262 698454
rect 290346 698218 290582 698454
rect 290026 697898 290262 698134
rect 290346 697898 290582 698134
rect 290026 671218 290262 671454
rect 290346 671218 290582 671454
rect 290026 670898 290262 671134
rect 290346 670898 290582 671134
rect 290026 644218 290262 644454
rect 290346 644218 290582 644454
rect 290026 643898 290262 644134
rect 290346 643898 290582 644134
rect 290026 617218 290262 617454
rect 290346 617218 290582 617454
rect 290026 616898 290262 617134
rect 290346 616898 290582 617134
rect 290026 590218 290262 590454
rect 290346 590218 290582 590454
rect 290026 589898 290262 590134
rect 290346 589898 290582 590134
rect 290026 563218 290262 563454
rect 290346 563218 290582 563454
rect 290026 562898 290262 563134
rect 290346 562898 290582 563134
rect 290026 536218 290262 536454
rect 290346 536218 290582 536454
rect 290026 535898 290262 536134
rect 290346 535898 290582 536134
rect 290026 509218 290262 509454
rect 290346 509218 290582 509454
rect 290026 508898 290262 509134
rect 290346 508898 290582 509134
rect 290026 482218 290262 482454
rect 290346 482218 290582 482454
rect 290026 481898 290262 482134
rect 290346 481898 290582 482134
rect 290026 455218 290262 455454
rect 290346 455218 290582 455454
rect 290026 454898 290262 455134
rect 290346 454898 290582 455134
rect 290026 428218 290262 428454
rect 290346 428218 290582 428454
rect 290026 427898 290262 428134
rect 290346 427898 290582 428134
rect 290026 401218 290262 401454
rect 290346 401218 290582 401454
rect 290026 400898 290262 401134
rect 290346 400898 290582 401134
rect 290026 374218 290262 374454
rect 290346 374218 290582 374454
rect 290026 373898 290262 374134
rect 290346 373898 290582 374134
rect 290026 347218 290262 347454
rect 290346 347218 290582 347454
rect 290026 346898 290262 347134
rect 290346 346898 290582 347134
rect 290026 320218 290262 320454
rect 290346 320218 290582 320454
rect 290026 319898 290262 320134
rect 290346 319898 290582 320134
rect 290026 293218 290262 293454
rect 290346 293218 290582 293454
rect 290026 292898 290262 293134
rect 290346 292898 290582 293134
rect 290026 266218 290262 266454
rect 290346 266218 290582 266454
rect 290026 265898 290262 266134
rect 290346 265898 290582 266134
rect 290026 239218 290262 239454
rect 290346 239218 290582 239454
rect 290026 238898 290262 239134
rect 290346 238898 290582 239134
rect 290026 212218 290262 212454
rect 290346 212218 290582 212454
rect 290026 211898 290262 212134
rect 290346 211898 290582 212134
rect 290026 185218 290262 185454
rect 290346 185218 290582 185454
rect 290026 184898 290262 185134
rect 290346 184898 290582 185134
rect 290026 158218 290262 158454
rect 290346 158218 290582 158454
rect 290026 157898 290262 158134
rect 290346 157898 290582 158134
rect 290026 131218 290262 131454
rect 290346 131218 290582 131454
rect 290026 130898 290262 131134
rect 290346 130898 290582 131134
rect 290026 104218 290262 104454
rect 290346 104218 290582 104454
rect 290026 103898 290262 104134
rect 290346 103898 290582 104134
rect 290026 77218 290262 77454
rect 290346 77218 290582 77454
rect 290026 76898 290262 77134
rect 290346 76898 290582 77134
rect 293526 704602 293762 704838
rect 293846 704602 294082 704838
rect 293526 704282 293762 704518
rect 293846 704282 294082 704518
rect 293526 701593 293762 701829
rect 293846 701593 294082 701829
rect 293526 701273 293762 701509
rect 293846 701273 294082 701509
rect 293526 674593 293762 674829
rect 293846 674593 294082 674829
rect 293526 674273 293762 674509
rect 293846 674273 294082 674509
rect 293526 647593 293762 647829
rect 293846 647593 294082 647829
rect 293526 647273 293762 647509
rect 293846 647273 294082 647509
rect 293526 620593 293762 620829
rect 293846 620593 294082 620829
rect 293526 620273 293762 620509
rect 293846 620273 294082 620509
rect 293526 593593 293762 593829
rect 293846 593593 294082 593829
rect 293526 593273 293762 593509
rect 293846 593273 294082 593509
rect 293526 566593 293762 566829
rect 293846 566593 294082 566829
rect 293526 566273 293762 566509
rect 293846 566273 294082 566509
rect 293526 539593 293762 539829
rect 293846 539593 294082 539829
rect 293526 539273 293762 539509
rect 293846 539273 294082 539509
rect 293526 512593 293762 512829
rect 293846 512593 294082 512829
rect 293526 512273 293762 512509
rect 293846 512273 294082 512509
rect 293526 485593 293762 485829
rect 293846 485593 294082 485829
rect 293526 485273 293762 485509
rect 293846 485273 294082 485509
rect 293526 458593 293762 458829
rect 293846 458593 294082 458829
rect 293526 458273 293762 458509
rect 293846 458273 294082 458509
rect 293526 431593 293762 431829
rect 293846 431593 294082 431829
rect 293526 431273 293762 431509
rect 293846 431273 294082 431509
rect 293526 404593 293762 404829
rect 293846 404593 294082 404829
rect 293526 404273 293762 404509
rect 293846 404273 294082 404509
rect 293526 377593 293762 377829
rect 293846 377593 294082 377829
rect 293526 377273 293762 377509
rect 293846 377273 294082 377509
rect 293526 350593 293762 350829
rect 293846 350593 294082 350829
rect 293526 350273 293762 350509
rect 293846 350273 294082 350509
rect 293526 323593 293762 323829
rect 293846 323593 294082 323829
rect 293526 323273 293762 323509
rect 293846 323273 294082 323509
rect 293526 296593 293762 296829
rect 293846 296593 294082 296829
rect 293526 296273 293762 296509
rect 293846 296273 294082 296509
rect 293526 269593 293762 269829
rect 293846 269593 294082 269829
rect 293526 269273 293762 269509
rect 293846 269273 294082 269509
rect 293526 242593 293762 242829
rect 293846 242593 294082 242829
rect 293526 242273 293762 242509
rect 293846 242273 294082 242509
rect 293526 215593 293762 215829
rect 293846 215593 294082 215829
rect 293526 215273 293762 215509
rect 293846 215273 294082 215509
rect 293526 188593 293762 188829
rect 293846 188593 294082 188829
rect 293526 188273 293762 188509
rect 293846 188273 294082 188509
rect 293526 161593 293762 161829
rect 293846 161593 294082 161829
rect 293526 161273 293762 161509
rect 293846 161273 294082 161509
rect 293526 134593 293762 134829
rect 293846 134593 294082 134829
rect 293526 134273 293762 134509
rect 293846 134273 294082 134509
rect 293526 107593 293762 107829
rect 293846 107593 294082 107829
rect 293526 107273 293762 107509
rect 293846 107273 294082 107509
rect 293526 80593 293762 80829
rect 293846 80593 294082 80829
rect 293526 80273 293762 80509
rect 293846 80273 294082 80509
rect 318026 705562 318262 705798
rect 318346 705562 318582 705798
rect 318026 705242 318262 705478
rect 318346 705242 318582 705478
rect 318026 698218 318262 698454
rect 318346 698218 318582 698454
rect 318026 697898 318262 698134
rect 318346 697898 318582 698134
rect 318026 671218 318262 671454
rect 318346 671218 318582 671454
rect 318026 670898 318262 671134
rect 318346 670898 318582 671134
rect 318026 644218 318262 644454
rect 318346 644218 318582 644454
rect 318026 643898 318262 644134
rect 318346 643898 318582 644134
rect 318026 617218 318262 617454
rect 318346 617218 318582 617454
rect 318026 616898 318262 617134
rect 318346 616898 318582 617134
rect 318026 590218 318262 590454
rect 318346 590218 318582 590454
rect 318026 589898 318262 590134
rect 318346 589898 318582 590134
rect 318026 563218 318262 563454
rect 318346 563218 318582 563454
rect 318026 562898 318262 563134
rect 318346 562898 318582 563134
rect 318026 536218 318262 536454
rect 318346 536218 318582 536454
rect 318026 535898 318262 536134
rect 318346 535898 318582 536134
rect 318026 509218 318262 509454
rect 318346 509218 318582 509454
rect 318026 508898 318262 509134
rect 318346 508898 318582 509134
rect 318026 482218 318262 482454
rect 318346 482218 318582 482454
rect 318026 481898 318262 482134
rect 318346 481898 318582 482134
rect 318026 455218 318262 455454
rect 318346 455218 318582 455454
rect 318026 454898 318262 455134
rect 318346 454898 318582 455134
rect 318026 428218 318262 428454
rect 318346 428218 318582 428454
rect 318026 427898 318262 428134
rect 318346 427898 318582 428134
rect 318026 401218 318262 401454
rect 318346 401218 318582 401454
rect 318026 400898 318262 401134
rect 318346 400898 318582 401134
rect 318026 374218 318262 374454
rect 318346 374218 318582 374454
rect 318026 373898 318262 374134
rect 318346 373898 318582 374134
rect 318026 347218 318262 347454
rect 318346 347218 318582 347454
rect 318026 346898 318262 347134
rect 318346 346898 318582 347134
rect 318026 320218 318262 320454
rect 318346 320218 318582 320454
rect 318026 319898 318262 320134
rect 318346 319898 318582 320134
rect 318026 293218 318262 293454
rect 318346 293218 318582 293454
rect 318026 292898 318262 293134
rect 318346 292898 318582 293134
rect 318026 266218 318262 266454
rect 318346 266218 318582 266454
rect 318026 265898 318262 266134
rect 318346 265898 318582 266134
rect 318026 239218 318262 239454
rect 318346 239218 318582 239454
rect 318026 238898 318262 239134
rect 318346 238898 318582 239134
rect 318026 212218 318262 212454
rect 318346 212218 318582 212454
rect 318026 211898 318262 212134
rect 318346 211898 318582 212134
rect 318026 185218 318262 185454
rect 318346 185218 318582 185454
rect 318026 184898 318262 185134
rect 318346 184898 318582 185134
rect 318026 158218 318262 158454
rect 318346 158218 318582 158454
rect 318026 157898 318262 158134
rect 318346 157898 318582 158134
rect 318026 131218 318262 131454
rect 318346 131218 318582 131454
rect 318026 130898 318262 131134
rect 318346 130898 318582 131134
rect 318026 104218 318262 104454
rect 318346 104218 318582 104454
rect 318026 103898 318262 104134
rect 318346 103898 318582 104134
rect 318026 77218 318262 77454
rect 318346 77218 318582 77454
rect 318026 76898 318262 77134
rect 318346 76898 318582 77134
rect 321526 704602 321762 704838
rect 321846 704602 322082 704838
rect 321526 704282 321762 704518
rect 321846 704282 322082 704518
rect 321526 701593 321762 701829
rect 321846 701593 322082 701829
rect 321526 701273 321762 701509
rect 321846 701273 322082 701509
rect 321526 674593 321762 674829
rect 321846 674593 322082 674829
rect 321526 674273 321762 674509
rect 321846 674273 322082 674509
rect 321526 647593 321762 647829
rect 321846 647593 322082 647829
rect 321526 647273 321762 647509
rect 321846 647273 322082 647509
rect 321526 620593 321762 620829
rect 321846 620593 322082 620829
rect 321526 620273 321762 620509
rect 321846 620273 322082 620509
rect 321526 593593 321762 593829
rect 321846 593593 322082 593829
rect 321526 593273 321762 593509
rect 321846 593273 322082 593509
rect 321526 566593 321762 566829
rect 321846 566593 322082 566829
rect 321526 566273 321762 566509
rect 321846 566273 322082 566509
rect 321526 539593 321762 539829
rect 321846 539593 322082 539829
rect 321526 539273 321762 539509
rect 321846 539273 322082 539509
rect 321526 512593 321762 512829
rect 321846 512593 322082 512829
rect 321526 512273 321762 512509
rect 321846 512273 322082 512509
rect 321526 485593 321762 485829
rect 321846 485593 322082 485829
rect 321526 485273 321762 485509
rect 321846 485273 322082 485509
rect 321526 458593 321762 458829
rect 321846 458593 322082 458829
rect 321526 458273 321762 458509
rect 321846 458273 322082 458509
rect 321526 431593 321762 431829
rect 321846 431593 322082 431829
rect 321526 431273 321762 431509
rect 321846 431273 322082 431509
rect 321526 404593 321762 404829
rect 321846 404593 322082 404829
rect 321526 404273 321762 404509
rect 321846 404273 322082 404509
rect 321526 377593 321762 377829
rect 321846 377593 322082 377829
rect 321526 377273 321762 377509
rect 321846 377273 322082 377509
rect 321526 350593 321762 350829
rect 321846 350593 322082 350829
rect 321526 350273 321762 350509
rect 321846 350273 322082 350509
rect 321526 323593 321762 323829
rect 321846 323593 322082 323829
rect 321526 323273 321762 323509
rect 321846 323273 322082 323509
rect 321526 296593 321762 296829
rect 321846 296593 322082 296829
rect 321526 296273 321762 296509
rect 321846 296273 322082 296509
rect 321526 269593 321762 269829
rect 321846 269593 322082 269829
rect 321526 269273 321762 269509
rect 321846 269273 322082 269509
rect 321526 242593 321762 242829
rect 321846 242593 322082 242829
rect 321526 242273 321762 242509
rect 321846 242273 322082 242509
rect 321526 215593 321762 215829
rect 321846 215593 322082 215829
rect 321526 215273 321762 215509
rect 321846 215273 322082 215509
rect 321526 188593 321762 188829
rect 321846 188593 322082 188829
rect 321526 188273 321762 188509
rect 321846 188273 322082 188509
rect 321526 161593 321762 161829
rect 321846 161593 322082 161829
rect 321526 161273 321762 161509
rect 321846 161273 322082 161509
rect 321526 134593 321762 134829
rect 321846 134593 322082 134829
rect 321526 134273 321762 134509
rect 321846 134273 322082 134509
rect 321526 107593 321762 107829
rect 321846 107593 322082 107829
rect 321526 107273 321762 107509
rect 321846 107273 322082 107509
rect 321526 80593 321762 80829
rect 321846 80593 322082 80829
rect 321526 80273 321762 80509
rect 321846 80273 322082 80509
rect 346026 705562 346262 705798
rect 346346 705562 346582 705798
rect 346026 705242 346262 705478
rect 346346 705242 346582 705478
rect 346026 698218 346262 698454
rect 346346 698218 346582 698454
rect 346026 697898 346262 698134
rect 346346 697898 346582 698134
rect 346026 671218 346262 671454
rect 346346 671218 346582 671454
rect 346026 670898 346262 671134
rect 346346 670898 346582 671134
rect 346026 644218 346262 644454
rect 346346 644218 346582 644454
rect 346026 643898 346262 644134
rect 346346 643898 346582 644134
rect 346026 617218 346262 617454
rect 346346 617218 346582 617454
rect 346026 616898 346262 617134
rect 346346 616898 346582 617134
rect 346026 590218 346262 590454
rect 346346 590218 346582 590454
rect 346026 589898 346262 590134
rect 346346 589898 346582 590134
rect 346026 563218 346262 563454
rect 346346 563218 346582 563454
rect 346026 562898 346262 563134
rect 346346 562898 346582 563134
rect 346026 536218 346262 536454
rect 346346 536218 346582 536454
rect 346026 535898 346262 536134
rect 346346 535898 346582 536134
rect 346026 509218 346262 509454
rect 346346 509218 346582 509454
rect 346026 508898 346262 509134
rect 346346 508898 346582 509134
rect 346026 482218 346262 482454
rect 346346 482218 346582 482454
rect 346026 481898 346262 482134
rect 346346 481898 346582 482134
rect 346026 455218 346262 455454
rect 346346 455218 346582 455454
rect 346026 454898 346262 455134
rect 346346 454898 346582 455134
rect 346026 428218 346262 428454
rect 346346 428218 346582 428454
rect 346026 427898 346262 428134
rect 346346 427898 346582 428134
rect 346026 401218 346262 401454
rect 346346 401218 346582 401454
rect 346026 400898 346262 401134
rect 346346 400898 346582 401134
rect 346026 374218 346262 374454
rect 346346 374218 346582 374454
rect 346026 373898 346262 374134
rect 346346 373898 346582 374134
rect 346026 347218 346262 347454
rect 346346 347218 346582 347454
rect 346026 346898 346262 347134
rect 346346 346898 346582 347134
rect 346026 320218 346262 320454
rect 346346 320218 346582 320454
rect 346026 319898 346262 320134
rect 346346 319898 346582 320134
rect 346026 293218 346262 293454
rect 346346 293218 346582 293454
rect 346026 292898 346262 293134
rect 346346 292898 346582 293134
rect 346026 266218 346262 266454
rect 346346 266218 346582 266454
rect 346026 265898 346262 266134
rect 346346 265898 346582 266134
rect 346026 239218 346262 239454
rect 346346 239218 346582 239454
rect 346026 238898 346262 239134
rect 346346 238898 346582 239134
rect 346026 212218 346262 212454
rect 346346 212218 346582 212454
rect 346026 211898 346262 212134
rect 346346 211898 346582 212134
rect 346026 185218 346262 185454
rect 346346 185218 346582 185454
rect 346026 184898 346262 185134
rect 346346 184898 346582 185134
rect 346026 158218 346262 158454
rect 346346 158218 346582 158454
rect 346026 157898 346262 158134
rect 346346 157898 346582 158134
rect 346026 131218 346262 131454
rect 346346 131218 346582 131454
rect 346026 130898 346262 131134
rect 346346 130898 346582 131134
rect 346026 104218 346262 104454
rect 346346 104218 346582 104454
rect 346026 103898 346262 104134
rect 346346 103898 346582 104134
rect 346026 77218 346262 77454
rect 346346 77218 346582 77454
rect 346026 76898 346262 77134
rect 346346 76898 346582 77134
rect 349526 704602 349762 704838
rect 349846 704602 350082 704838
rect 349526 704282 349762 704518
rect 349846 704282 350082 704518
rect 349526 701593 349762 701829
rect 349846 701593 350082 701829
rect 349526 701273 349762 701509
rect 349846 701273 350082 701509
rect 349526 674593 349762 674829
rect 349846 674593 350082 674829
rect 349526 674273 349762 674509
rect 349846 674273 350082 674509
rect 349526 647593 349762 647829
rect 349846 647593 350082 647829
rect 349526 647273 349762 647509
rect 349846 647273 350082 647509
rect 349526 620593 349762 620829
rect 349846 620593 350082 620829
rect 349526 620273 349762 620509
rect 349846 620273 350082 620509
rect 349526 593593 349762 593829
rect 349846 593593 350082 593829
rect 349526 593273 349762 593509
rect 349846 593273 350082 593509
rect 349526 566593 349762 566829
rect 349846 566593 350082 566829
rect 349526 566273 349762 566509
rect 349846 566273 350082 566509
rect 349526 539593 349762 539829
rect 349846 539593 350082 539829
rect 349526 539273 349762 539509
rect 349846 539273 350082 539509
rect 349526 512593 349762 512829
rect 349846 512593 350082 512829
rect 349526 512273 349762 512509
rect 349846 512273 350082 512509
rect 349526 485593 349762 485829
rect 349846 485593 350082 485829
rect 349526 485273 349762 485509
rect 349846 485273 350082 485509
rect 349526 458593 349762 458829
rect 349846 458593 350082 458829
rect 349526 458273 349762 458509
rect 349846 458273 350082 458509
rect 349526 431593 349762 431829
rect 349846 431593 350082 431829
rect 349526 431273 349762 431509
rect 349846 431273 350082 431509
rect 349526 404593 349762 404829
rect 349846 404593 350082 404829
rect 349526 404273 349762 404509
rect 349846 404273 350082 404509
rect 349526 377593 349762 377829
rect 349846 377593 350082 377829
rect 349526 377273 349762 377509
rect 349846 377273 350082 377509
rect 349526 350593 349762 350829
rect 349846 350593 350082 350829
rect 349526 350273 349762 350509
rect 349846 350273 350082 350509
rect 349526 323593 349762 323829
rect 349846 323593 350082 323829
rect 349526 323273 349762 323509
rect 349846 323273 350082 323509
rect 349526 296593 349762 296829
rect 349846 296593 350082 296829
rect 349526 296273 349762 296509
rect 349846 296273 350082 296509
rect 349526 269593 349762 269829
rect 349846 269593 350082 269829
rect 349526 269273 349762 269509
rect 349846 269273 350082 269509
rect 349526 242593 349762 242829
rect 349846 242593 350082 242829
rect 349526 242273 349762 242509
rect 349846 242273 350082 242509
rect 349526 215593 349762 215829
rect 349846 215593 350082 215829
rect 349526 215273 349762 215509
rect 349846 215273 350082 215509
rect 349526 188593 349762 188829
rect 349846 188593 350082 188829
rect 349526 188273 349762 188509
rect 349846 188273 350082 188509
rect 349526 161593 349762 161829
rect 349846 161593 350082 161829
rect 349526 161273 349762 161509
rect 349846 161273 350082 161509
rect 349526 134593 349762 134829
rect 349846 134593 350082 134829
rect 349526 134273 349762 134509
rect 349846 134273 350082 134509
rect 349526 107593 349762 107829
rect 349846 107593 350082 107829
rect 349526 107273 349762 107509
rect 349846 107273 350082 107509
rect 349526 80593 349762 80829
rect 349846 80593 350082 80829
rect 349526 80273 349762 80509
rect 349846 80273 350082 80509
rect 374026 705562 374262 705798
rect 374346 705562 374582 705798
rect 374026 705242 374262 705478
rect 374346 705242 374582 705478
rect 374026 698218 374262 698454
rect 374346 698218 374582 698454
rect 374026 697898 374262 698134
rect 374346 697898 374582 698134
rect 374026 671218 374262 671454
rect 374346 671218 374582 671454
rect 374026 670898 374262 671134
rect 374346 670898 374582 671134
rect 374026 644218 374262 644454
rect 374346 644218 374582 644454
rect 374026 643898 374262 644134
rect 374346 643898 374582 644134
rect 374026 617218 374262 617454
rect 374346 617218 374582 617454
rect 374026 616898 374262 617134
rect 374346 616898 374582 617134
rect 374026 590218 374262 590454
rect 374346 590218 374582 590454
rect 374026 589898 374262 590134
rect 374346 589898 374582 590134
rect 374026 563218 374262 563454
rect 374346 563218 374582 563454
rect 374026 562898 374262 563134
rect 374346 562898 374582 563134
rect 374026 536218 374262 536454
rect 374346 536218 374582 536454
rect 374026 535898 374262 536134
rect 374346 535898 374582 536134
rect 374026 509218 374262 509454
rect 374346 509218 374582 509454
rect 374026 508898 374262 509134
rect 374346 508898 374582 509134
rect 374026 482218 374262 482454
rect 374346 482218 374582 482454
rect 374026 481898 374262 482134
rect 374346 481898 374582 482134
rect 374026 455218 374262 455454
rect 374346 455218 374582 455454
rect 374026 454898 374262 455134
rect 374346 454898 374582 455134
rect 374026 428218 374262 428454
rect 374346 428218 374582 428454
rect 374026 427898 374262 428134
rect 374346 427898 374582 428134
rect 374026 401218 374262 401454
rect 374346 401218 374582 401454
rect 374026 400898 374262 401134
rect 374346 400898 374582 401134
rect 374026 374218 374262 374454
rect 374346 374218 374582 374454
rect 374026 373898 374262 374134
rect 374346 373898 374582 374134
rect 374026 347218 374262 347454
rect 374346 347218 374582 347454
rect 374026 346898 374262 347134
rect 374346 346898 374582 347134
rect 374026 320218 374262 320454
rect 374346 320218 374582 320454
rect 374026 319898 374262 320134
rect 374346 319898 374582 320134
rect 374026 293218 374262 293454
rect 374346 293218 374582 293454
rect 374026 292898 374262 293134
rect 374346 292898 374582 293134
rect 374026 266218 374262 266454
rect 374346 266218 374582 266454
rect 374026 265898 374262 266134
rect 374346 265898 374582 266134
rect 374026 239218 374262 239454
rect 374346 239218 374582 239454
rect 374026 238898 374262 239134
rect 374346 238898 374582 239134
rect 374026 212218 374262 212454
rect 374346 212218 374582 212454
rect 374026 211898 374262 212134
rect 374346 211898 374582 212134
rect 374026 185218 374262 185454
rect 374346 185218 374582 185454
rect 374026 184898 374262 185134
rect 374346 184898 374582 185134
rect 374026 158218 374262 158454
rect 374346 158218 374582 158454
rect 374026 157898 374262 158134
rect 374346 157898 374582 158134
rect 374026 131218 374262 131454
rect 374346 131218 374582 131454
rect 374026 130898 374262 131134
rect 374346 130898 374582 131134
rect 374026 104218 374262 104454
rect 374346 104218 374582 104454
rect 374026 103898 374262 104134
rect 374346 103898 374582 104134
rect 374026 77218 374262 77454
rect 374346 77218 374582 77454
rect 374026 76898 374262 77134
rect 374346 76898 374582 77134
rect 377526 704602 377762 704838
rect 377846 704602 378082 704838
rect 377526 704282 377762 704518
rect 377846 704282 378082 704518
rect 377526 701593 377762 701829
rect 377846 701593 378082 701829
rect 377526 701273 377762 701509
rect 377846 701273 378082 701509
rect 402026 705562 402262 705798
rect 402346 705562 402582 705798
rect 402026 705242 402262 705478
rect 402346 705242 402582 705478
rect 377526 674593 377762 674829
rect 377846 674593 378082 674829
rect 377526 674273 377762 674509
rect 377846 674273 378082 674509
rect 377526 647593 377762 647829
rect 377846 647593 378082 647829
rect 377526 647273 377762 647509
rect 377846 647273 378082 647509
rect 377526 620593 377762 620829
rect 377846 620593 378082 620829
rect 377526 620273 377762 620509
rect 377846 620273 378082 620509
rect 377526 593593 377762 593829
rect 377846 593593 378082 593829
rect 377526 593273 377762 593509
rect 377846 593273 378082 593509
rect 377526 566593 377762 566829
rect 377846 566593 378082 566829
rect 377526 566273 377762 566509
rect 377846 566273 378082 566509
rect 377526 539593 377762 539829
rect 377846 539593 378082 539829
rect 377526 539273 377762 539509
rect 377846 539273 378082 539509
rect 377526 512593 377762 512829
rect 377846 512593 378082 512829
rect 377526 512273 377762 512509
rect 377846 512273 378082 512509
rect 377526 485593 377762 485829
rect 377846 485593 378082 485829
rect 377526 485273 377762 485509
rect 377846 485273 378082 485509
rect 377526 458593 377762 458829
rect 377846 458593 378082 458829
rect 377526 458273 377762 458509
rect 377846 458273 378082 458509
rect 377526 431593 377762 431829
rect 377846 431593 378082 431829
rect 377526 431273 377762 431509
rect 377846 431273 378082 431509
rect 377526 404593 377762 404829
rect 377846 404593 378082 404829
rect 377526 404273 377762 404509
rect 377846 404273 378082 404509
rect 377526 377593 377762 377829
rect 377846 377593 378082 377829
rect 377526 377273 377762 377509
rect 377846 377273 378082 377509
rect 377526 350593 377762 350829
rect 377846 350593 378082 350829
rect 377526 350273 377762 350509
rect 377846 350273 378082 350509
rect 377526 323593 377762 323829
rect 377846 323593 378082 323829
rect 377526 323273 377762 323509
rect 377846 323273 378082 323509
rect 377526 296593 377762 296829
rect 377846 296593 378082 296829
rect 377526 296273 377762 296509
rect 377846 296273 378082 296509
rect 377526 269593 377762 269829
rect 377846 269593 378082 269829
rect 377526 269273 377762 269509
rect 377846 269273 378082 269509
rect 377526 242593 377762 242829
rect 377846 242593 378082 242829
rect 377526 242273 377762 242509
rect 377846 242273 378082 242509
rect 377526 215593 377762 215829
rect 377846 215593 378082 215829
rect 377526 215273 377762 215509
rect 377846 215273 378082 215509
rect 377526 188593 377762 188829
rect 377846 188593 378082 188829
rect 377526 188273 377762 188509
rect 377846 188273 378082 188509
rect 377526 161593 377762 161829
rect 377846 161593 378082 161829
rect 377526 161273 377762 161509
rect 377846 161273 378082 161509
rect 377526 134593 377762 134829
rect 377846 134593 378082 134829
rect 377526 134273 377762 134509
rect 377846 134273 378082 134509
rect 377526 107593 377762 107829
rect 377846 107593 378082 107829
rect 377526 107273 377762 107509
rect 377846 107273 378082 107509
rect 377526 80593 377762 80829
rect 377846 80593 378082 80829
rect 377526 80273 377762 80509
rect 377846 80273 378082 80509
rect 181526 53593 181762 53829
rect 181846 53593 182082 53829
rect 181526 53273 181762 53509
rect 181846 53273 182082 53509
rect 192960 53593 193196 53829
rect 192960 53273 193196 53509
rect 196908 53593 197144 53829
rect 196908 53273 197144 53509
rect 200856 53593 201092 53829
rect 200856 53273 201092 53509
rect 204804 53593 205040 53829
rect 204804 53273 205040 53509
rect 213260 53593 213496 53829
rect 213260 53273 213496 53509
rect 214208 53593 214444 53829
rect 214208 53273 214444 53509
rect 215156 53593 215392 53829
rect 215156 53273 215392 53509
rect 216104 53593 216340 53829
rect 216104 53273 216340 53509
rect 221960 53593 222196 53829
rect 221960 53273 222196 53509
rect 225908 53593 226144 53829
rect 225908 53273 226144 53509
rect 229856 53593 230092 53829
rect 229856 53273 230092 53509
rect 233804 53593 234040 53829
rect 233804 53273 234040 53509
rect 242260 53593 242496 53829
rect 242260 53273 242496 53509
rect 243208 53593 243444 53829
rect 243208 53273 243444 53509
rect 244156 53593 244392 53829
rect 244156 53273 244392 53509
rect 245104 53593 245340 53829
rect 245104 53273 245340 53509
rect 194934 50218 195170 50454
rect 194934 49898 195170 50134
rect 198882 50218 199118 50454
rect 198882 49898 199118 50134
rect 202830 50218 203066 50454
rect 202830 49898 203066 50134
rect 213734 50218 213970 50454
rect 213734 49898 213970 50134
rect 214682 50218 214918 50454
rect 214682 49898 214918 50134
rect 215630 50218 215866 50454
rect 215630 49898 215866 50134
rect 223934 50218 224170 50454
rect 223934 49898 224170 50134
rect 227882 50218 228118 50454
rect 227882 49898 228118 50134
rect 231830 50218 232066 50454
rect 231830 49898 232066 50134
rect 242734 50218 242970 50454
rect 242734 49898 242970 50134
rect 243682 50218 243918 50454
rect 243682 49898 243918 50134
rect 244630 50218 244866 50454
rect 244630 49898 244866 50134
rect 250960 53593 251196 53829
rect 250960 53273 251196 53509
rect 254908 53593 255144 53829
rect 254908 53273 255144 53509
rect 258856 53593 259092 53829
rect 258856 53273 259092 53509
rect 262804 53593 263040 53829
rect 262804 53273 263040 53509
rect 271260 53593 271496 53829
rect 271260 53273 271496 53509
rect 272208 53593 272444 53829
rect 272208 53273 272444 53509
rect 273156 53593 273392 53829
rect 273156 53273 273392 53509
rect 274104 53593 274340 53829
rect 274104 53273 274340 53509
rect 252934 50218 253170 50454
rect 252934 49898 253170 50134
rect 256882 50218 257118 50454
rect 256882 49898 257118 50134
rect 260830 50218 261066 50454
rect 260830 49898 261066 50134
rect 271734 50218 271970 50454
rect 271734 49898 271970 50134
rect 272682 50218 272918 50454
rect 272682 49898 272918 50134
rect 273630 50218 273866 50454
rect 273630 49898 273866 50134
rect 279960 53593 280196 53829
rect 279960 53273 280196 53509
rect 283908 53593 284144 53829
rect 283908 53273 284144 53509
rect 287856 53593 288092 53829
rect 287856 53273 288092 53509
rect 291804 53593 292040 53829
rect 291804 53273 292040 53509
rect 300260 53593 300496 53829
rect 300260 53273 300496 53509
rect 301208 53593 301444 53829
rect 301208 53273 301444 53509
rect 302156 53593 302392 53829
rect 302156 53273 302392 53509
rect 303104 53593 303340 53829
rect 303104 53273 303340 53509
rect 281934 50218 282170 50454
rect 281934 49898 282170 50134
rect 285882 50218 286118 50454
rect 285882 49898 286118 50134
rect 289830 50218 290066 50454
rect 289830 49898 290066 50134
rect 300734 50218 300970 50454
rect 300734 49898 300970 50134
rect 301682 50218 301918 50454
rect 301682 49898 301918 50134
rect 302630 50218 302866 50454
rect 302630 49898 302866 50134
rect 308960 53593 309196 53829
rect 308960 53273 309196 53509
rect 312908 53593 313144 53829
rect 312908 53273 313144 53509
rect 316856 53593 317092 53829
rect 316856 53273 317092 53509
rect 320804 53593 321040 53829
rect 320804 53273 321040 53509
rect 329260 53593 329496 53829
rect 329260 53273 329496 53509
rect 330208 53593 330444 53829
rect 330208 53273 330444 53509
rect 331156 53593 331392 53829
rect 331156 53273 331392 53509
rect 332104 53593 332340 53829
rect 332104 53273 332340 53509
rect 310934 50218 311170 50454
rect 310934 49898 311170 50134
rect 314882 50218 315118 50454
rect 314882 49898 315118 50134
rect 318830 50218 319066 50454
rect 318830 49898 319066 50134
rect 329734 50218 329970 50454
rect 329734 49898 329970 50134
rect 330682 50218 330918 50454
rect 330682 49898 330918 50134
rect 331630 50218 331866 50454
rect 331630 49898 331866 50134
rect 337960 53593 338196 53829
rect 337960 53273 338196 53509
rect 341908 53593 342144 53829
rect 341908 53273 342144 53509
rect 345856 53593 346092 53829
rect 345856 53273 346092 53509
rect 349804 53593 350040 53829
rect 349804 53273 350040 53509
rect 358260 53593 358496 53829
rect 358260 53273 358496 53509
rect 359208 53593 359444 53829
rect 359208 53273 359444 53509
rect 360156 53593 360392 53829
rect 360156 53273 360392 53509
rect 361104 53593 361340 53829
rect 361104 53273 361340 53509
rect 339934 50218 340170 50454
rect 339934 49898 340170 50134
rect 343882 50218 344118 50454
rect 343882 49898 344118 50134
rect 347830 50218 348066 50454
rect 347830 49898 348066 50134
rect 358734 50218 358970 50454
rect 358734 49898 358970 50134
rect 359682 50218 359918 50454
rect 359682 49898 359918 50134
rect 360630 50218 360866 50454
rect 360630 49898 360866 50134
rect 366960 53593 367196 53829
rect 366960 53273 367196 53509
rect 370908 53593 371144 53829
rect 370908 53273 371144 53509
rect 374856 53593 375092 53829
rect 374856 53273 375092 53509
rect 378804 53593 379040 53829
rect 378804 53273 379040 53509
rect 387260 53593 387496 53829
rect 387260 53273 387496 53509
rect 388208 53593 388444 53829
rect 388208 53273 388444 53509
rect 389156 53593 389392 53829
rect 389156 53273 389392 53509
rect 390104 53593 390340 53829
rect 390104 53273 390340 53509
rect 368934 50218 369170 50454
rect 368934 49898 369170 50134
rect 372882 50218 373118 50454
rect 372882 49898 373118 50134
rect 376830 50218 377066 50454
rect 376830 49898 377066 50134
rect 387734 50218 387970 50454
rect 387734 49898 387970 50134
rect 388682 50218 388918 50454
rect 388682 49898 388918 50134
rect 389630 50218 389866 50454
rect 389630 49898 389866 50134
rect 395960 53593 396196 53829
rect 395960 53273 396196 53509
rect 171160 26593 171396 26829
rect 171160 26273 171396 26509
rect 175108 26593 175344 26829
rect 175108 26273 175344 26509
rect 179056 26593 179292 26829
rect 179056 26273 179292 26509
rect 183004 26593 183240 26829
rect 183004 26273 183240 26509
rect 191460 26593 191696 26829
rect 191460 26273 191696 26509
rect 192408 26593 192644 26829
rect 192408 26273 192644 26509
rect 193356 26593 193592 26829
rect 193356 26273 193592 26509
rect 194304 26593 194540 26829
rect 194304 26273 194540 26509
rect 200160 26593 200396 26829
rect 200160 26273 200396 26509
rect 204108 26593 204344 26829
rect 204108 26273 204344 26509
rect 208056 26593 208292 26829
rect 208056 26273 208292 26509
rect 212004 26593 212240 26829
rect 212004 26273 212240 26509
rect 220460 26593 220696 26829
rect 220460 26273 220696 26509
rect 221408 26593 221644 26829
rect 221408 26273 221644 26509
rect 222356 26593 222592 26829
rect 222356 26273 222592 26509
rect 223304 26593 223540 26829
rect 223304 26273 223540 26509
rect 229160 26593 229396 26829
rect 229160 26273 229396 26509
rect 233108 26593 233344 26829
rect 233108 26273 233344 26509
rect 237056 26593 237292 26829
rect 237056 26273 237292 26509
rect 241004 26593 241240 26829
rect 241004 26273 241240 26509
rect 249460 26593 249696 26829
rect 249460 26273 249696 26509
rect 250408 26593 250644 26829
rect 250408 26273 250644 26509
rect 251356 26593 251592 26829
rect 251356 26273 251592 26509
rect 252304 26593 252540 26829
rect 252304 26273 252540 26509
rect 258160 26593 258396 26829
rect 258160 26273 258396 26509
rect 262108 26593 262344 26829
rect 262108 26273 262344 26509
rect 266056 26593 266292 26829
rect 266056 26273 266292 26509
rect 270004 26593 270240 26829
rect 270004 26273 270240 26509
rect 278460 26593 278696 26829
rect 278460 26273 278696 26509
rect 279408 26593 279644 26829
rect 279408 26273 279644 26509
rect 280356 26593 280592 26829
rect 280356 26273 280592 26509
rect 281304 26593 281540 26829
rect 281304 26273 281540 26509
rect 287160 26593 287396 26829
rect 287160 26273 287396 26509
rect 291108 26593 291344 26829
rect 291108 26273 291344 26509
rect 295056 26593 295292 26829
rect 295056 26273 295292 26509
rect 299004 26593 299240 26829
rect 299004 26273 299240 26509
rect 307460 26593 307696 26829
rect 307460 26273 307696 26509
rect 308408 26593 308644 26829
rect 308408 26273 308644 26509
rect 309356 26593 309592 26829
rect 309356 26273 309592 26509
rect 310304 26593 310540 26829
rect 310304 26273 310540 26509
rect 316160 26593 316396 26829
rect 316160 26273 316396 26509
rect 320108 26593 320344 26829
rect 320108 26273 320344 26509
rect 324056 26593 324292 26829
rect 324056 26273 324292 26509
rect 328004 26593 328240 26829
rect 328004 26273 328240 26509
rect 336460 26593 336696 26829
rect 336460 26273 336696 26509
rect 337408 26593 337644 26829
rect 337408 26273 337644 26509
rect 338356 26593 338592 26829
rect 338356 26273 338592 26509
rect 339304 26593 339540 26829
rect 339304 26273 339540 26509
rect 345160 26593 345396 26829
rect 345160 26273 345396 26509
rect 349108 26593 349344 26829
rect 349108 26273 349344 26509
rect 353056 26593 353292 26829
rect 353056 26273 353292 26509
rect 357004 26593 357240 26829
rect 357004 26273 357240 26509
rect 365460 26593 365696 26829
rect 365460 26273 365696 26509
rect 366408 26593 366644 26829
rect 366408 26273 366644 26509
rect 367356 26593 367592 26829
rect 367356 26273 367592 26509
rect 368304 26593 368540 26829
rect 368304 26273 368540 26509
rect 374160 26593 374396 26829
rect 374160 26273 374396 26509
rect 378108 26593 378344 26829
rect 378108 26273 378344 26509
rect 382056 26593 382292 26829
rect 382056 26273 382292 26509
rect 386004 26593 386240 26829
rect 386004 26273 386240 26509
rect 394460 26593 394696 26829
rect 394460 26273 394696 26509
rect 395408 26593 395644 26829
rect 395408 26273 395644 26509
rect 396356 26593 396592 26829
rect 396356 26273 396592 26509
rect 397304 26593 397540 26829
rect 397304 26273 397540 26509
rect 173134 23218 173370 23454
rect 173134 22898 173370 23134
rect 177082 23218 177318 23454
rect 177082 22898 177318 23134
rect 181030 23218 181266 23454
rect 181030 22898 181266 23134
rect 191934 23218 192170 23454
rect 191934 22898 192170 23134
rect 192882 23218 193118 23454
rect 192882 22898 193118 23134
rect 193830 23218 194066 23454
rect 193830 22898 194066 23134
rect 202134 23218 202370 23454
rect 202134 22898 202370 23134
rect 206082 23218 206318 23454
rect 206082 22898 206318 23134
rect 210030 23218 210266 23454
rect 210030 22898 210266 23134
rect 220934 23218 221170 23454
rect 220934 22898 221170 23134
rect 221882 23218 222118 23454
rect 221882 22898 222118 23134
rect 222830 23218 223066 23454
rect 222830 22898 223066 23134
rect 231134 23218 231370 23454
rect 231134 22898 231370 23134
rect 235082 23218 235318 23454
rect 235082 22898 235318 23134
rect 239030 23218 239266 23454
rect 239030 22898 239266 23134
rect 249934 23218 250170 23454
rect 249934 22898 250170 23134
rect 250882 23218 251118 23454
rect 250882 22898 251118 23134
rect 251830 23218 252066 23454
rect 251830 22898 252066 23134
rect 260134 23218 260370 23454
rect 260134 22898 260370 23134
rect 264082 23218 264318 23454
rect 264082 22898 264318 23134
rect 268030 23218 268266 23454
rect 268030 22898 268266 23134
rect 278934 23218 279170 23454
rect 278934 22898 279170 23134
rect 279882 23218 280118 23454
rect 279882 22898 280118 23134
rect 280830 23218 281066 23454
rect 280830 22898 281066 23134
rect 289134 23218 289370 23454
rect 289134 22898 289370 23134
rect 293082 23218 293318 23454
rect 293082 22898 293318 23134
rect 297030 23218 297266 23454
rect 297030 22898 297266 23134
rect 307934 23218 308170 23454
rect 307934 22898 308170 23134
rect 308882 23218 309118 23454
rect 308882 22898 309118 23134
rect 309830 23218 310066 23454
rect 309830 22898 310066 23134
rect 318134 23218 318370 23454
rect 318134 22898 318370 23134
rect 322082 23218 322318 23454
rect 322082 22898 322318 23134
rect 326030 23218 326266 23454
rect 326030 22898 326266 23134
rect 336934 23218 337170 23454
rect 336934 22898 337170 23134
rect 337882 23218 338118 23454
rect 337882 22898 338118 23134
rect 338830 23218 339066 23454
rect 338830 22898 339066 23134
rect 347134 23218 347370 23454
rect 347134 22898 347370 23134
rect 351082 23218 351318 23454
rect 351082 22898 351318 23134
rect 355030 23218 355266 23454
rect 355030 22898 355266 23134
rect 365934 23218 366170 23454
rect 365934 22898 366170 23134
rect 366882 23218 367118 23454
rect 366882 22898 367118 23134
rect 367830 23218 368066 23454
rect 367830 22898 368066 23134
rect 376134 23218 376370 23454
rect 376134 22898 376370 23134
rect 380082 23218 380318 23454
rect 380082 22898 380318 23134
rect 384030 23218 384266 23454
rect 384030 22898 384266 23134
rect 394934 23218 395170 23454
rect 394934 22898 395170 23134
rect 395882 23218 396118 23454
rect 395882 22898 396118 23134
rect 396830 23218 397066 23454
rect 396830 22898 397066 23134
rect 402026 698218 402262 698454
rect 402346 698218 402582 698454
rect 402026 697898 402262 698134
rect 402346 697898 402582 698134
rect 402026 671218 402262 671454
rect 402346 671218 402582 671454
rect 402026 670898 402262 671134
rect 402346 670898 402582 671134
rect 402026 644218 402262 644454
rect 402346 644218 402582 644454
rect 402026 643898 402262 644134
rect 402346 643898 402582 644134
rect 402026 617218 402262 617454
rect 402346 617218 402582 617454
rect 402026 616898 402262 617134
rect 402346 616898 402582 617134
rect 402026 590218 402262 590454
rect 402346 590218 402582 590454
rect 402026 589898 402262 590134
rect 402346 589898 402582 590134
rect 402026 563218 402262 563454
rect 402346 563218 402582 563454
rect 402026 562898 402262 563134
rect 402346 562898 402582 563134
rect 402026 536218 402262 536454
rect 402346 536218 402582 536454
rect 402026 535898 402262 536134
rect 402346 535898 402582 536134
rect 402026 509218 402262 509454
rect 402346 509218 402582 509454
rect 402026 508898 402262 509134
rect 402346 508898 402582 509134
rect 402026 482218 402262 482454
rect 402346 482218 402582 482454
rect 402026 481898 402262 482134
rect 402346 481898 402582 482134
rect 402026 455218 402262 455454
rect 402346 455218 402582 455454
rect 402026 454898 402262 455134
rect 402346 454898 402582 455134
rect 402026 428218 402262 428454
rect 402346 428218 402582 428454
rect 402026 427898 402262 428134
rect 402346 427898 402582 428134
rect 402026 401218 402262 401454
rect 402346 401218 402582 401454
rect 402026 400898 402262 401134
rect 402346 400898 402582 401134
rect 402026 374218 402262 374454
rect 402346 374218 402582 374454
rect 402026 373898 402262 374134
rect 402346 373898 402582 374134
rect 402026 347218 402262 347454
rect 402346 347218 402582 347454
rect 402026 346898 402262 347134
rect 402346 346898 402582 347134
rect 402026 320218 402262 320454
rect 402346 320218 402582 320454
rect 402026 319898 402262 320134
rect 402346 319898 402582 320134
rect 402026 293218 402262 293454
rect 402346 293218 402582 293454
rect 402026 292898 402262 293134
rect 402346 292898 402582 293134
rect 402026 266218 402262 266454
rect 402346 266218 402582 266454
rect 402026 265898 402262 266134
rect 402346 265898 402582 266134
rect 402026 239218 402262 239454
rect 402346 239218 402582 239454
rect 402026 238898 402262 239134
rect 402346 238898 402582 239134
rect 402026 212218 402262 212454
rect 402346 212218 402582 212454
rect 402026 211898 402262 212134
rect 402346 211898 402582 212134
rect 402026 185218 402262 185454
rect 402346 185218 402582 185454
rect 402026 184898 402262 185134
rect 402346 184898 402582 185134
rect 402026 158218 402262 158454
rect 402346 158218 402582 158454
rect 402026 157898 402262 158134
rect 402346 157898 402582 158134
rect 402026 131218 402262 131454
rect 402346 131218 402582 131454
rect 402026 130898 402262 131134
rect 402346 130898 402582 131134
rect 402026 104218 402262 104454
rect 402346 104218 402582 104454
rect 402026 103898 402262 104134
rect 402346 103898 402582 104134
rect 402026 77218 402262 77454
rect 402346 77218 402582 77454
rect 402026 76898 402262 77134
rect 402346 76898 402582 77134
rect 405526 704602 405762 704838
rect 405846 704602 406082 704838
rect 405526 704282 405762 704518
rect 405846 704282 406082 704518
rect 405526 701593 405762 701829
rect 405846 701593 406082 701829
rect 405526 701273 405762 701509
rect 405846 701273 406082 701509
rect 430026 705562 430262 705798
rect 430346 705562 430582 705798
rect 430026 705242 430262 705478
rect 430346 705242 430582 705478
rect 405526 674593 405762 674829
rect 405846 674593 406082 674829
rect 405526 674273 405762 674509
rect 405846 674273 406082 674509
rect 405526 647593 405762 647829
rect 405846 647593 406082 647829
rect 405526 647273 405762 647509
rect 405846 647273 406082 647509
rect 405526 620593 405762 620829
rect 405846 620593 406082 620829
rect 405526 620273 405762 620509
rect 405846 620273 406082 620509
rect 405526 593593 405762 593829
rect 405846 593593 406082 593829
rect 405526 593273 405762 593509
rect 405846 593273 406082 593509
rect 405526 566593 405762 566829
rect 405846 566593 406082 566829
rect 405526 566273 405762 566509
rect 405846 566273 406082 566509
rect 405526 539593 405762 539829
rect 405846 539593 406082 539829
rect 405526 539273 405762 539509
rect 405846 539273 406082 539509
rect 405526 512593 405762 512829
rect 405846 512593 406082 512829
rect 405526 512273 405762 512509
rect 405846 512273 406082 512509
rect 405526 485593 405762 485829
rect 405846 485593 406082 485829
rect 405526 485273 405762 485509
rect 405846 485273 406082 485509
rect 405526 458593 405762 458829
rect 405846 458593 406082 458829
rect 405526 458273 405762 458509
rect 405846 458273 406082 458509
rect 405526 431593 405762 431829
rect 405846 431593 406082 431829
rect 405526 431273 405762 431509
rect 405846 431273 406082 431509
rect 405526 404593 405762 404829
rect 405846 404593 406082 404829
rect 405526 404273 405762 404509
rect 405846 404273 406082 404509
rect 405526 377593 405762 377829
rect 405846 377593 406082 377829
rect 405526 377273 405762 377509
rect 405846 377273 406082 377509
rect 405526 350593 405762 350829
rect 405846 350593 406082 350829
rect 405526 350273 405762 350509
rect 405846 350273 406082 350509
rect 405526 323593 405762 323829
rect 405846 323593 406082 323829
rect 405526 323273 405762 323509
rect 405846 323273 406082 323509
rect 405526 296593 405762 296829
rect 405846 296593 406082 296829
rect 405526 296273 405762 296509
rect 405846 296273 406082 296509
rect 405526 269593 405762 269829
rect 405846 269593 406082 269829
rect 405526 269273 405762 269509
rect 405846 269273 406082 269509
rect 405526 242593 405762 242829
rect 405846 242593 406082 242829
rect 405526 242273 405762 242509
rect 405846 242273 406082 242509
rect 405526 215593 405762 215829
rect 405846 215593 406082 215829
rect 405526 215273 405762 215509
rect 405846 215273 406082 215509
rect 405526 188593 405762 188829
rect 405846 188593 406082 188829
rect 405526 188273 405762 188509
rect 405846 188273 406082 188509
rect 405526 161593 405762 161829
rect 405846 161593 406082 161829
rect 405526 161273 405762 161509
rect 405846 161273 406082 161509
rect 405526 134593 405762 134829
rect 405846 134593 406082 134829
rect 405526 134273 405762 134509
rect 405846 134273 406082 134509
rect 405526 107593 405762 107829
rect 405846 107593 406082 107829
rect 405526 107273 405762 107509
rect 405846 107273 406082 107509
rect 405526 80593 405762 80829
rect 405846 80593 406082 80829
rect 405526 80273 405762 80509
rect 405846 80273 406082 80509
rect 399908 53593 400144 53829
rect 399908 53273 400144 53509
rect 403856 53593 404092 53829
rect 403856 53273 404092 53509
rect 407804 53593 408040 53829
rect 407804 53273 408040 53509
rect 416260 53593 416496 53829
rect 416260 53273 416496 53509
rect 417208 53593 417444 53829
rect 417208 53273 417444 53509
rect 418156 53593 418392 53829
rect 418156 53273 418392 53509
rect 419104 53593 419340 53829
rect 419104 53273 419340 53509
rect 397934 50218 398170 50454
rect 397934 49898 398170 50134
rect 401882 50218 402118 50454
rect 401882 49898 402118 50134
rect 405830 50218 406066 50454
rect 405830 49898 406066 50134
rect 416734 50218 416970 50454
rect 416734 49898 416970 50134
rect 417682 50218 417918 50454
rect 417682 49898 417918 50134
rect 418630 50218 418866 50454
rect 418630 49898 418866 50134
rect 424960 53593 425196 53829
rect 424960 53273 425196 53509
rect 428908 53593 429144 53829
rect 428908 53273 429144 53509
rect 426934 50218 427170 50454
rect 426934 49898 427170 50134
rect 403160 26593 403396 26829
rect 403160 26273 403396 26509
rect 407108 26593 407344 26829
rect 407108 26273 407344 26509
rect 411056 26593 411292 26829
rect 411056 26273 411292 26509
rect 415004 26593 415240 26829
rect 415004 26273 415240 26509
rect 423460 26593 423696 26829
rect 423460 26273 423696 26509
rect 424408 26593 424644 26829
rect 424408 26273 424644 26509
rect 425356 26593 425592 26829
rect 425356 26273 425592 26509
rect 426304 26593 426540 26829
rect 426304 26273 426540 26509
rect 405134 23218 405370 23454
rect 405134 22898 405370 23134
rect 409082 23218 409318 23454
rect 409082 22898 409318 23134
rect 413030 23218 413266 23454
rect 413030 22898 413266 23134
rect 423934 23218 424170 23454
rect 423934 22898 424170 23134
rect 424882 23218 425118 23454
rect 424882 22898 425118 23134
rect 425830 23218 426066 23454
rect 425830 22898 426066 23134
rect 430026 698218 430262 698454
rect 430346 698218 430582 698454
rect 430026 697898 430262 698134
rect 430346 697898 430582 698134
rect 430026 671218 430262 671454
rect 430346 671218 430582 671454
rect 430026 670898 430262 671134
rect 430346 670898 430582 671134
rect 430026 644218 430262 644454
rect 430346 644218 430582 644454
rect 430026 643898 430262 644134
rect 430346 643898 430582 644134
rect 430026 617218 430262 617454
rect 430346 617218 430582 617454
rect 430026 616898 430262 617134
rect 430346 616898 430582 617134
rect 430026 590218 430262 590454
rect 430346 590218 430582 590454
rect 430026 589898 430262 590134
rect 430346 589898 430582 590134
rect 430026 563218 430262 563454
rect 430346 563218 430582 563454
rect 430026 562898 430262 563134
rect 430346 562898 430582 563134
rect 430026 536218 430262 536454
rect 430346 536218 430582 536454
rect 430026 535898 430262 536134
rect 430346 535898 430582 536134
rect 430026 509218 430262 509454
rect 430346 509218 430582 509454
rect 430026 508898 430262 509134
rect 430346 508898 430582 509134
rect 430026 482218 430262 482454
rect 430346 482218 430582 482454
rect 430026 481898 430262 482134
rect 430346 481898 430582 482134
rect 430026 455218 430262 455454
rect 430346 455218 430582 455454
rect 430026 454898 430262 455134
rect 430346 454898 430582 455134
rect 430026 428218 430262 428454
rect 430346 428218 430582 428454
rect 430026 427898 430262 428134
rect 430346 427898 430582 428134
rect 430026 401218 430262 401454
rect 430346 401218 430582 401454
rect 430026 400898 430262 401134
rect 430346 400898 430582 401134
rect 430026 374218 430262 374454
rect 430346 374218 430582 374454
rect 430026 373898 430262 374134
rect 430346 373898 430582 374134
rect 430026 347218 430262 347454
rect 430346 347218 430582 347454
rect 430026 346898 430262 347134
rect 430346 346898 430582 347134
rect 430026 320218 430262 320454
rect 430346 320218 430582 320454
rect 430026 319898 430262 320134
rect 430346 319898 430582 320134
rect 430026 293218 430262 293454
rect 430346 293218 430582 293454
rect 430026 292898 430262 293134
rect 430346 292898 430582 293134
rect 430026 266218 430262 266454
rect 430346 266218 430582 266454
rect 430026 265898 430262 266134
rect 430346 265898 430582 266134
rect 430026 239218 430262 239454
rect 430346 239218 430582 239454
rect 430026 238898 430262 239134
rect 430346 238898 430582 239134
rect 430026 212218 430262 212454
rect 430346 212218 430582 212454
rect 430026 211898 430262 212134
rect 430346 211898 430582 212134
rect 430026 185218 430262 185454
rect 430346 185218 430582 185454
rect 430026 184898 430262 185134
rect 430346 184898 430582 185134
rect 430026 158218 430262 158454
rect 430346 158218 430582 158454
rect 430026 157898 430262 158134
rect 430346 157898 430582 158134
rect 430026 131218 430262 131454
rect 430346 131218 430582 131454
rect 430026 130898 430262 131134
rect 430346 130898 430582 131134
rect 430026 104218 430262 104454
rect 430346 104218 430582 104454
rect 430026 103898 430262 104134
rect 430346 103898 430582 104134
rect 430026 77218 430262 77454
rect 430346 77218 430582 77454
rect 430026 76898 430262 77134
rect 430346 76898 430582 77134
rect 433526 704602 433762 704838
rect 433846 704602 434082 704838
rect 433526 704282 433762 704518
rect 433846 704282 434082 704518
rect 433526 701593 433762 701829
rect 433846 701593 434082 701829
rect 433526 701273 433762 701509
rect 433846 701273 434082 701509
rect 433526 674593 433762 674829
rect 433846 674593 434082 674829
rect 433526 674273 433762 674509
rect 433846 674273 434082 674509
rect 433526 647593 433762 647829
rect 433846 647593 434082 647829
rect 433526 647273 433762 647509
rect 433846 647273 434082 647509
rect 433526 620593 433762 620829
rect 433846 620593 434082 620829
rect 433526 620273 433762 620509
rect 433846 620273 434082 620509
rect 433526 593593 433762 593829
rect 433846 593593 434082 593829
rect 433526 593273 433762 593509
rect 433846 593273 434082 593509
rect 433526 566593 433762 566829
rect 433846 566593 434082 566829
rect 433526 566273 433762 566509
rect 433846 566273 434082 566509
rect 433526 539593 433762 539829
rect 433846 539593 434082 539829
rect 433526 539273 433762 539509
rect 433846 539273 434082 539509
rect 433526 512593 433762 512829
rect 433846 512593 434082 512829
rect 433526 512273 433762 512509
rect 433846 512273 434082 512509
rect 433526 485593 433762 485829
rect 433846 485593 434082 485829
rect 433526 485273 433762 485509
rect 433846 485273 434082 485509
rect 433526 458593 433762 458829
rect 433846 458593 434082 458829
rect 433526 458273 433762 458509
rect 433846 458273 434082 458509
rect 433526 431593 433762 431829
rect 433846 431593 434082 431829
rect 433526 431273 433762 431509
rect 433846 431273 434082 431509
rect 433526 404593 433762 404829
rect 433846 404593 434082 404829
rect 433526 404273 433762 404509
rect 433846 404273 434082 404509
rect 433526 377593 433762 377829
rect 433846 377593 434082 377829
rect 433526 377273 433762 377509
rect 433846 377273 434082 377509
rect 433526 350593 433762 350829
rect 433846 350593 434082 350829
rect 433526 350273 433762 350509
rect 433846 350273 434082 350509
rect 433526 323593 433762 323829
rect 433846 323593 434082 323829
rect 433526 323273 433762 323509
rect 433846 323273 434082 323509
rect 433526 296593 433762 296829
rect 433846 296593 434082 296829
rect 433526 296273 433762 296509
rect 433846 296273 434082 296509
rect 433526 269593 433762 269829
rect 433846 269593 434082 269829
rect 433526 269273 433762 269509
rect 433846 269273 434082 269509
rect 433526 242593 433762 242829
rect 433846 242593 434082 242829
rect 433526 242273 433762 242509
rect 433846 242273 434082 242509
rect 433526 215593 433762 215829
rect 433846 215593 434082 215829
rect 433526 215273 433762 215509
rect 433846 215273 434082 215509
rect 433526 188593 433762 188829
rect 433846 188593 434082 188829
rect 433526 188273 433762 188509
rect 433846 188273 434082 188509
rect 433526 161593 433762 161829
rect 433846 161593 434082 161829
rect 433526 161273 433762 161509
rect 433846 161273 434082 161509
rect 433526 134593 433762 134829
rect 433846 134593 434082 134829
rect 433526 134273 433762 134509
rect 433846 134273 434082 134509
rect 433526 107593 433762 107829
rect 433846 107593 434082 107829
rect 433526 107273 433762 107509
rect 433846 107273 434082 107509
rect 433526 80593 433762 80829
rect 433846 80593 434082 80829
rect 433526 80273 433762 80509
rect 433846 80273 434082 80509
rect 458026 705562 458262 705798
rect 458346 705562 458582 705798
rect 458026 705242 458262 705478
rect 458346 705242 458582 705478
rect 458026 698218 458262 698454
rect 458346 698218 458582 698454
rect 458026 697898 458262 698134
rect 458346 697898 458582 698134
rect 458026 671218 458262 671454
rect 458346 671218 458582 671454
rect 458026 670898 458262 671134
rect 458346 670898 458582 671134
rect 458026 644218 458262 644454
rect 458346 644218 458582 644454
rect 458026 643898 458262 644134
rect 458346 643898 458582 644134
rect 458026 617218 458262 617454
rect 458346 617218 458582 617454
rect 458026 616898 458262 617134
rect 458346 616898 458582 617134
rect 458026 590218 458262 590454
rect 458346 590218 458582 590454
rect 458026 589898 458262 590134
rect 458346 589898 458582 590134
rect 458026 563218 458262 563454
rect 458346 563218 458582 563454
rect 458026 562898 458262 563134
rect 458346 562898 458582 563134
rect 458026 536218 458262 536454
rect 458346 536218 458582 536454
rect 458026 535898 458262 536134
rect 458346 535898 458582 536134
rect 458026 509218 458262 509454
rect 458346 509218 458582 509454
rect 458026 508898 458262 509134
rect 458346 508898 458582 509134
rect 458026 482218 458262 482454
rect 458346 482218 458582 482454
rect 458026 481898 458262 482134
rect 458346 481898 458582 482134
rect 458026 455218 458262 455454
rect 458346 455218 458582 455454
rect 458026 454898 458262 455134
rect 458346 454898 458582 455134
rect 458026 428218 458262 428454
rect 458346 428218 458582 428454
rect 458026 427898 458262 428134
rect 458346 427898 458582 428134
rect 458026 401218 458262 401454
rect 458346 401218 458582 401454
rect 458026 400898 458262 401134
rect 458346 400898 458582 401134
rect 458026 374218 458262 374454
rect 458346 374218 458582 374454
rect 458026 373898 458262 374134
rect 458346 373898 458582 374134
rect 458026 347218 458262 347454
rect 458346 347218 458582 347454
rect 458026 346898 458262 347134
rect 458346 346898 458582 347134
rect 458026 320218 458262 320454
rect 458346 320218 458582 320454
rect 458026 319898 458262 320134
rect 458346 319898 458582 320134
rect 458026 293218 458262 293454
rect 458346 293218 458582 293454
rect 458026 292898 458262 293134
rect 458346 292898 458582 293134
rect 458026 266218 458262 266454
rect 458346 266218 458582 266454
rect 458026 265898 458262 266134
rect 458346 265898 458582 266134
rect 458026 239218 458262 239454
rect 458346 239218 458582 239454
rect 458026 238898 458262 239134
rect 458346 238898 458582 239134
rect 458026 212218 458262 212454
rect 458346 212218 458582 212454
rect 458026 211898 458262 212134
rect 458346 211898 458582 212134
rect 458026 185218 458262 185454
rect 458346 185218 458582 185454
rect 458026 184898 458262 185134
rect 458346 184898 458582 185134
rect 458026 158218 458262 158454
rect 458346 158218 458582 158454
rect 458026 157898 458262 158134
rect 458346 157898 458582 158134
rect 458026 131218 458262 131454
rect 458346 131218 458582 131454
rect 458026 130898 458262 131134
rect 458346 130898 458582 131134
rect 458026 104218 458262 104454
rect 458346 104218 458582 104454
rect 458026 103898 458262 104134
rect 458346 103898 458582 104134
rect 458026 77218 458262 77454
rect 458346 77218 458582 77454
rect 458026 76898 458262 77134
rect 458346 76898 458582 77134
rect 461526 704602 461762 704838
rect 461846 704602 462082 704838
rect 461526 704282 461762 704518
rect 461846 704282 462082 704518
rect 461526 701593 461762 701829
rect 461846 701593 462082 701829
rect 461526 701273 461762 701509
rect 461846 701273 462082 701509
rect 461526 674593 461762 674829
rect 461846 674593 462082 674829
rect 461526 674273 461762 674509
rect 461846 674273 462082 674509
rect 461526 647593 461762 647829
rect 461846 647593 462082 647829
rect 461526 647273 461762 647509
rect 461846 647273 462082 647509
rect 461526 620593 461762 620829
rect 461846 620593 462082 620829
rect 461526 620273 461762 620509
rect 461846 620273 462082 620509
rect 461526 593593 461762 593829
rect 461846 593593 462082 593829
rect 461526 593273 461762 593509
rect 461846 593273 462082 593509
rect 461526 566593 461762 566829
rect 461846 566593 462082 566829
rect 461526 566273 461762 566509
rect 461846 566273 462082 566509
rect 461526 539593 461762 539829
rect 461846 539593 462082 539829
rect 461526 539273 461762 539509
rect 461846 539273 462082 539509
rect 461526 512593 461762 512829
rect 461846 512593 462082 512829
rect 461526 512273 461762 512509
rect 461846 512273 462082 512509
rect 461526 485593 461762 485829
rect 461846 485593 462082 485829
rect 461526 485273 461762 485509
rect 461846 485273 462082 485509
rect 461526 458593 461762 458829
rect 461846 458593 462082 458829
rect 461526 458273 461762 458509
rect 461846 458273 462082 458509
rect 461526 431593 461762 431829
rect 461846 431593 462082 431829
rect 461526 431273 461762 431509
rect 461846 431273 462082 431509
rect 461526 404593 461762 404829
rect 461846 404593 462082 404829
rect 461526 404273 461762 404509
rect 461846 404273 462082 404509
rect 461526 377593 461762 377829
rect 461846 377593 462082 377829
rect 461526 377273 461762 377509
rect 461846 377273 462082 377509
rect 461526 350593 461762 350829
rect 461846 350593 462082 350829
rect 461526 350273 461762 350509
rect 461846 350273 462082 350509
rect 461526 323593 461762 323829
rect 461846 323593 462082 323829
rect 461526 323273 461762 323509
rect 461846 323273 462082 323509
rect 461526 296593 461762 296829
rect 461846 296593 462082 296829
rect 461526 296273 461762 296509
rect 461846 296273 462082 296509
rect 461526 269593 461762 269829
rect 461846 269593 462082 269829
rect 461526 269273 461762 269509
rect 461846 269273 462082 269509
rect 461526 242593 461762 242829
rect 461846 242593 462082 242829
rect 461526 242273 461762 242509
rect 461846 242273 462082 242509
rect 461526 215593 461762 215829
rect 461846 215593 462082 215829
rect 461526 215273 461762 215509
rect 461846 215273 462082 215509
rect 461526 188593 461762 188829
rect 461846 188593 462082 188829
rect 461526 188273 461762 188509
rect 461846 188273 462082 188509
rect 461526 161593 461762 161829
rect 461846 161593 462082 161829
rect 461526 161273 461762 161509
rect 461846 161273 462082 161509
rect 461526 134593 461762 134829
rect 461846 134593 462082 134829
rect 461526 134273 461762 134509
rect 461846 134273 462082 134509
rect 461526 107593 461762 107829
rect 461846 107593 462082 107829
rect 461526 107273 461762 107509
rect 461846 107273 462082 107509
rect 461526 80593 461762 80829
rect 461846 80593 462082 80829
rect 461526 80273 461762 80509
rect 461846 80273 462082 80509
rect 486026 705562 486262 705798
rect 486346 705562 486582 705798
rect 486026 705242 486262 705478
rect 486346 705242 486582 705478
rect 486026 698218 486262 698454
rect 486346 698218 486582 698454
rect 486026 697898 486262 698134
rect 486346 697898 486582 698134
rect 486026 671218 486262 671454
rect 486346 671218 486582 671454
rect 486026 670898 486262 671134
rect 486346 670898 486582 671134
rect 486026 644218 486262 644454
rect 486346 644218 486582 644454
rect 486026 643898 486262 644134
rect 486346 643898 486582 644134
rect 486026 617218 486262 617454
rect 486346 617218 486582 617454
rect 486026 616898 486262 617134
rect 486346 616898 486582 617134
rect 486026 590218 486262 590454
rect 486346 590218 486582 590454
rect 486026 589898 486262 590134
rect 486346 589898 486582 590134
rect 486026 563218 486262 563454
rect 486346 563218 486582 563454
rect 486026 562898 486262 563134
rect 486346 562898 486582 563134
rect 486026 536218 486262 536454
rect 486346 536218 486582 536454
rect 486026 535898 486262 536134
rect 486346 535898 486582 536134
rect 486026 509218 486262 509454
rect 486346 509218 486582 509454
rect 486026 508898 486262 509134
rect 486346 508898 486582 509134
rect 486026 482218 486262 482454
rect 486346 482218 486582 482454
rect 486026 481898 486262 482134
rect 486346 481898 486582 482134
rect 486026 455218 486262 455454
rect 486346 455218 486582 455454
rect 486026 454898 486262 455134
rect 486346 454898 486582 455134
rect 486026 428218 486262 428454
rect 486346 428218 486582 428454
rect 486026 427898 486262 428134
rect 486346 427898 486582 428134
rect 486026 401218 486262 401454
rect 486346 401218 486582 401454
rect 486026 400898 486262 401134
rect 486346 400898 486582 401134
rect 486026 374218 486262 374454
rect 486346 374218 486582 374454
rect 486026 373898 486262 374134
rect 486346 373898 486582 374134
rect 486026 347218 486262 347454
rect 486346 347218 486582 347454
rect 486026 346898 486262 347134
rect 486346 346898 486582 347134
rect 486026 320218 486262 320454
rect 486346 320218 486582 320454
rect 486026 319898 486262 320134
rect 486346 319898 486582 320134
rect 486026 293218 486262 293454
rect 486346 293218 486582 293454
rect 486026 292898 486262 293134
rect 486346 292898 486582 293134
rect 486026 266218 486262 266454
rect 486346 266218 486582 266454
rect 486026 265898 486262 266134
rect 486346 265898 486582 266134
rect 486026 239218 486262 239454
rect 486346 239218 486582 239454
rect 486026 238898 486262 239134
rect 486346 238898 486582 239134
rect 486026 212218 486262 212454
rect 486346 212218 486582 212454
rect 486026 211898 486262 212134
rect 486346 211898 486582 212134
rect 486026 185218 486262 185454
rect 486346 185218 486582 185454
rect 486026 184898 486262 185134
rect 486346 184898 486582 185134
rect 486026 158218 486262 158454
rect 486346 158218 486582 158454
rect 486026 157898 486262 158134
rect 486346 157898 486582 158134
rect 486026 131218 486262 131454
rect 486346 131218 486582 131454
rect 486026 130898 486262 131134
rect 486346 130898 486582 131134
rect 486026 104218 486262 104454
rect 486346 104218 486582 104454
rect 486026 103898 486262 104134
rect 486346 103898 486582 104134
rect 486026 77218 486262 77454
rect 486346 77218 486582 77454
rect 486026 76898 486262 77134
rect 486346 76898 486582 77134
rect 489526 704602 489762 704838
rect 489846 704602 490082 704838
rect 489526 704282 489762 704518
rect 489846 704282 490082 704518
rect 489526 701593 489762 701829
rect 489846 701593 490082 701829
rect 489526 701273 489762 701509
rect 489846 701273 490082 701509
rect 489526 674593 489762 674829
rect 489846 674593 490082 674829
rect 489526 674273 489762 674509
rect 489846 674273 490082 674509
rect 489526 647593 489762 647829
rect 489846 647593 490082 647829
rect 489526 647273 489762 647509
rect 489846 647273 490082 647509
rect 489526 620593 489762 620829
rect 489846 620593 490082 620829
rect 489526 620273 489762 620509
rect 489846 620273 490082 620509
rect 489526 593593 489762 593829
rect 489846 593593 490082 593829
rect 489526 593273 489762 593509
rect 489846 593273 490082 593509
rect 489526 566593 489762 566829
rect 489846 566593 490082 566829
rect 489526 566273 489762 566509
rect 489846 566273 490082 566509
rect 489526 539593 489762 539829
rect 489846 539593 490082 539829
rect 489526 539273 489762 539509
rect 489846 539273 490082 539509
rect 489526 512593 489762 512829
rect 489846 512593 490082 512829
rect 489526 512273 489762 512509
rect 489846 512273 490082 512509
rect 489526 485593 489762 485829
rect 489846 485593 490082 485829
rect 489526 485273 489762 485509
rect 489846 485273 490082 485509
rect 489526 458593 489762 458829
rect 489846 458593 490082 458829
rect 489526 458273 489762 458509
rect 489846 458273 490082 458509
rect 489526 431593 489762 431829
rect 489846 431593 490082 431829
rect 489526 431273 489762 431509
rect 489846 431273 490082 431509
rect 489526 404593 489762 404829
rect 489846 404593 490082 404829
rect 489526 404273 489762 404509
rect 489846 404273 490082 404509
rect 489526 377593 489762 377829
rect 489846 377593 490082 377829
rect 489526 377273 489762 377509
rect 489846 377273 490082 377509
rect 489526 350593 489762 350829
rect 489846 350593 490082 350829
rect 489526 350273 489762 350509
rect 489846 350273 490082 350509
rect 489526 323593 489762 323829
rect 489846 323593 490082 323829
rect 489526 323273 489762 323509
rect 489846 323273 490082 323509
rect 489526 296593 489762 296829
rect 489846 296593 490082 296829
rect 489526 296273 489762 296509
rect 489846 296273 490082 296509
rect 489526 269593 489762 269829
rect 489846 269593 490082 269829
rect 489526 269273 489762 269509
rect 489846 269273 490082 269509
rect 489526 242593 489762 242829
rect 489846 242593 490082 242829
rect 489526 242273 489762 242509
rect 489846 242273 490082 242509
rect 489526 215593 489762 215829
rect 489846 215593 490082 215829
rect 489526 215273 489762 215509
rect 489846 215273 490082 215509
rect 489526 188593 489762 188829
rect 489846 188593 490082 188829
rect 489526 188273 489762 188509
rect 489846 188273 490082 188509
rect 489526 161593 489762 161829
rect 489846 161593 490082 161829
rect 489526 161273 489762 161509
rect 489846 161273 490082 161509
rect 489526 134593 489762 134829
rect 489846 134593 490082 134829
rect 489526 134273 489762 134509
rect 489846 134273 490082 134509
rect 489526 107593 489762 107829
rect 489846 107593 490082 107829
rect 489526 107273 489762 107509
rect 489846 107273 490082 107509
rect 489526 80593 489762 80829
rect 489846 80593 490082 80829
rect 489526 80273 489762 80509
rect 489846 80273 490082 80509
rect 514026 705562 514262 705798
rect 514346 705562 514582 705798
rect 514026 705242 514262 705478
rect 514346 705242 514582 705478
rect 514026 698218 514262 698454
rect 514346 698218 514582 698454
rect 514026 697898 514262 698134
rect 514346 697898 514582 698134
rect 514026 671218 514262 671454
rect 514346 671218 514582 671454
rect 514026 670898 514262 671134
rect 514346 670898 514582 671134
rect 514026 644218 514262 644454
rect 514346 644218 514582 644454
rect 514026 643898 514262 644134
rect 514346 643898 514582 644134
rect 514026 617218 514262 617454
rect 514346 617218 514582 617454
rect 514026 616898 514262 617134
rect 514346 616898 514582 617134
rect 514026 590218 514262 590454
rect 514346 590218 514582 590454
rect 514026 589898 514262 590134
rect 514346 589898 514582 590134
rect 514026 563218 514262 563454
rect 514346 563218 514582 563454
rect 514026 562898 514262 563134
rect 514346 562898 514582 563134
rect 514026 536218 514262 536454
rect 514346 536218 514582 536454
rect 514026 535898 514262 536134
rect 514346 535898 514582 536134
rect 514026 509218 514262 509454
rect 514346 509218 514582 509454
rect 514026 508898 514262 509134
rect 514346 508898 514582 509134
rect 514026 482218 514262 482454
rect 514346 482218 514582 482454
rect 514026 481898 514262 482134
rect 514346 481898 514582 482134
rect 514026 455218 514262 455454
rect 514346 455218 514582 455454
rect 514026 454898 514262 455134
rect 514346 454898 514582 455134
rect 514026 428218 514262 428454
rect 514346 428218 514582 428454
rect 514026 427898 514262 428134
rect 514346 427898 514582 428134
rect 514026 401218 514262 401454
rect 514346 401218 514582 401454
rect 514026 400898 514262 401134
rect 514346 400898 514582 401134
rect 514026 374218 514262 374454
rect 514346 374218 514582 374454
rect 514026 373898 514262 374134
rect 514346 373898 514582 374134
rect 514026 347218 514262 347454
rect 514346 347218 514582 347454
rect 514026 346898 514262 347134
rect 514346 346898 514582 347134
rect 514026 320218 514262 320454
rect 514346 320218 514582 320454
rect 514026 319898 514262 320134
rect 514346 319898 514582 320134
rect 514026 293218 514262 293454
rect 514346 293218 514582 293454
rect 514026 292898 514262 293134
rect 514346 292898 514582 293134
rect 514026 266218 514262 266454
rect 514346 266218 514582 266454
rect 514026 265898 514262 266134
rect 514346 265898 514582 266134
rect 514026 239218 514262 239454
rect 514346 239218 514582 239454
rect 514026 238898 514262 239134
rect 514346 238898 514582 239134
rect 514026 212218 514262 212454
rect 514346 212218 514582 212454
rect 514026 211898 514262 212134
rect 514346 211898 514582 212134
rect 514026 185218 514262 185454
rect 514346 185218 514582 185454
rect 514026 184898 514262 185134
rect 514346 184898 514582 185134
rect 514026 158218 514262 158454
rect 514346 158218 514582 158454
rect 514026 157898 514262 158134
rect 514346 157898 514582 158134
rect 514026 131218 514262 131454
rect 514346 131218 514582 131454
rect 514026 130898 514262 131134
rect 514346 130898 514582 131134
rect 514026 104218 514262 104454
rect 514346 104218 514582 104454
rect 514026 103898 514262 104134
rect 514346 103898 514582 104134
rect 514026 77218 514262 77454
rect 514346 77218 514582 77454
rect 514026 76898 514262 77134
rect 514346 76898 514582 77134
rect 517526 704602 517762 704838
rect 517846 704602 518082 704838
rect 517526 704282 517762 704518
rect 517846 704282 518082 704518
rect 517526 701593 517762 701829
rect 517846 701593 518082 701829
rect 517526 701273 517762 701509
rect 517846 701273 518082 701509
rect 542026 705562 542262 705798
rect 542346 705562 542582 705798
rect 542026 705242 542262 705478
rect 542346 705242 542582 705478
rect 517526 674593 517762 674829
rect 517846 674593 518082 674829
rect 517526 674273 517762 674509
rect 517846 674273 518082 674509
rect 517526 647593 517762 647829
rect 517846 647593 518082 647829
rect 517526 647273 517762 647509
rect 517846 647273 518082 647509
rect 517526 620593 517762 620829
rect 517846 620593 518082 620829
rect 517526 620273 517762 620509
rect 517846 620273 518082 620509
rect 517526 593593 517762 593829
rect 517846 593593 518082 593829
rect 517526 593273 517762 593509
rect 517846 593273 518082 593509
rect 517526 566593 517762 566829
rect 517846 566593 518082 566829
rect 517526 566273 517762 566509
rect 517846 566273 518082 566509
rect 517526 539593 517762 539829
rect 517846 539593 518082 539829
rect 517526 539273 517762 539509
rect 517846 539273 518082 539509
rect 517526 512593 517762 512829
rect 517846 512593 518082 512829
rect 517526 512273 517762 512509
rect 517846 512273 518082 512509
rect 517526 485593 517762 485829
rect 517846 485593 518082 485829
rect 517526 485273 517762 485509
rect 517846 485273 518082 485509
rect 517526 458593 517762 458829
rect 517846 458593 518082 458829
rect 517526 458273 517762 458509
rect 517846 458273 518082 458509
rect 517526 431593 517762 431829
rect 517846 431593 518082 431829
rect 517526 431273 517762 431509
rect 517846 431273 518082 431509
rect 517526 404593 517762 404829
rect 517846 404593 518082 404829
rect 517526 404273 517762 404509
rect 517846 404273 518082 404509
rect 517526 377593 517762 377829
rect 517846 377593 518082 377829
rect 517526 377273 517762 377509
rect 517846 377273 518082 377509
rect 517526 350593 517762 350829
rect 517846 350593 518082 350829
rect 517526 350273 517762 350509
rect 517846 350273 518082 350509
rect 517526 323593 517762 323829
rect 517846 323593 518082 323829
rect 517526 323273 517762 323509
rect 517846 323273 518082 323509
rect 517526 296593 517762 296829
rect 517846 296593 518082 296829
rect 517526 296273 517762 296509
rect 517846 296273 518082 296509
rect 517526 269593 517762 269829
rect 517846 269593 518082 269829
rect 517526 269273 517762 269509
rect 517846 269273 518082 269509
rect 517526 242593 517762 242829
rect 517846 242593 518082 242829
rect 517526 242273 517762 242509
rect 517846 242273 518082 242509
rect 517526 215593 517762 215829
rect 517846 215593 518082 215829
rect 517526 215273 517762 215509
rect 517846 215273 518082 215509
rect 517526 188593 517762 188829
rect 517846 188593 518082 188829
rect 517526 188273 517762 188509
rect 517846 188273 518082 188509
rect 517526 161593 517762 161829
rect 517846 161593 518082 161829
rect 517526 161273 517762 161509
rect 517846 161273 518082 161509
rect 517526 134593 517762 134829
rect 517846 134593 518082 134829
rect 517526 134273 517762 134509
rect 517846 134273 518082 134509
rect 517526 107593 517762 107829
rect 517846 107593 518082 107829
rect 517526 107273 517762 107509
rect 517846 107273 518082 107509
rect 517526 80593 517762 80829
rect 517846 80593 518082 80829
rect 517526 80273 517762 80509
rect 517846 80273 518082 80509
rect 432856 53593 433092 53829
rect 432856 53273 433092 53509
rect 436804 53593 437040 53829
rect 436804 53273 437040 53509
rect 445260 53593 445496 53829
rect 445260 53273 445496 53509
rect 446208 53593 446444 53829
rect 446208 53273 446444 53509
rect 447156 53593 447392 53829
rect 447156 53273 447392 53509
rect 448104 53593 448340 53829
rect 448104 53273 448340 53509
rect 453960 53593 454196 53829
rect 453960 53273 454196 53509
rect 457908 53593 458144 53829
rect 457908 53273 458144 53509
rect 461856 53593 462092 53829
rect 461856 53273 462092 53509
rect 465804 53593 466040 53829
rect 465804 53273 466040 53509
rect 474260 53593 474496 53829
rect 474260 53273 474496 53509
rect 475208 53593 475444 53829
rect 475208 53273 475444 53509
rect 476156 53593 476392 53829
rect 476156 53273 476392 53509
rect 477104 53593 477340 53829
rect 477104 53273 477340 53509
rect 482960 53593 483196 53829
rect 482960 53273 483196 53509
rect 486908 53593 487144 53829
rect 486908 53273 487144 53509
rect 490856 53593 491092 53829
rect 490856 53273 491092 53509
rect 494804 53593 495040 53829
rect 494804 53273 495040 53509
rect 503260 53593 503496 53829
rect 503260 53273 503496 53509
rect 504208 53593 504444 53829
rect 504208 53273 504444 53509
rect 505156 53593 505392 53829
rect 505156 53273 505392 53509
rect 506104 53593 506340 53829
rect 506104 53273 506340 53509
rect 511960 53593 512196 53829
rect 511960 53273 512196 53509
rect 515908 53593 516144 53829
rect 515908 53273 516144 53509
rect 519856 53593 520092 53829
rect 519856 53273 520092 53509
rect 523804 53593 524040 53829
rect 523804 53273 524040 53509
rect 430882 50218 431118 50454
rect 430882 49898 431118 50134
rect 434830 50218 435066 50454
rect 434830 49898 435066 50134
rect 445734 50218 445970 50454
rect 445734 49898 445970 50134
rect 446682 50218 446918 50454
rect 446682 49898 446918 50134
rect 447630 50218 447866 50454
rect 447630 49898 447866 50134
rect 455934 50218 456170 50454
rect 455934 49898 456170 50134
rect 459882 50218 460118 50454
rect 459882 49898 460118 50134
rect 463830 50218 464066 50454
rect 463830 49898 464066 50134
rect 474734 50218 474970 50454
rect 474734 49898 474970 50134
rect 475682 50218 475918 50454
rect 475682 49898 475918 50134
rect 476630 50218 476866 50454
rect 476630 49898 476866 50134
rect 484934 50218 485170 50454
rect 484934 49898 485170 50134
rect 488882 50218 489118 50454
rect 488882 49898 489118 50134
rect 492830 50218 493066 50454
rect 492830 49898 493066 50134
rect 503734 50218 503970 50454
rect 503734 49898 503970 50134
rect 504682 50218 504918 50454
rect 504682 49898 504918 50134
rect 505630 50218 505866 50454
rect 505630 49898 505866 50134
rect 513934 50218 514170 50454
rect 513934 49898 514170 50134
rect 517882 50218 518118 50454
rect 517882 49898 518118 50134
rect 521830 50218 522066 50454
rect 521830 49898 522066 50134
rect 432160 26593 432396 26829
rect 432160 26273 432396 26509
rect 436108 26593 436344 26829
rect 436108 26273 436344 26509
rect 440056 26593 440292 26829
rect 440056 26273 440292 26509
rect 444004 26593 444240 26829
rect 444004 26273 444240 26509
rect 452460 26593 452696 26829
rect 452460 26273 452696 26509
rect 453408 26593 453644 26829
rect 453408 26273 453644 26509
rect 454356 26593 454592 26829
rect 454356 26273 454592 26509
rect 455304 26593 455540 26829
rect 455304 26273 455540 26509
rect 461160 26593 461396 26829
rect 461160 26273 461396 26509
rect 465108 26593 465344 26829
rect 465108 26273 465344 26509
rect 469056 26593 469292 26829
rect 469056 26273 469292 26509
rect 473004 26593 473240 26829
rect 473004 26273 473240 26509
rect 481460 26593 481696 26829
rect 481460 26273 481696 26509
rect 482408 26593 482644 26829
rect 482408 26273 482644 26509
rect 483356 26593 483592 26829
rect 483356 26273 483592 26509
rect 484304 26593 484540 26829
rect 484304 26273 484540 26509
rect 490160 26593 490396 26829
rect 490160 26273 490396 26509
rect 494108 26593 494344 26829
rect 494108 26273 494344 26509
rect 498056 26593 498292 26829
rect 498056 26273 498292 26509
rect 502004 26593 502240 26829
rect 502004 26273 502240 26509
rect 510460 26593 510696 26829
rect 510460 26273 510696 26509
rect 511408 26593 511644 26829
rect 511408 26273 511644 26509
rect 512356 26593 512592 26829
rect 512356 26273 512592 26509
rect 513304 26593 513540 26829
rect 513304 26273 513540 26509
rect 519160 26593 519396 26829
rect 519160 26273 519396 26509
rect 523108 26593 523344 26829
rect 523108 26273 523344 26509
rect 527056 26593 527292 26829
rect 527056 26273 527292 26509
rect 434134 23218 434370 23454
rect 434134 22898 434370 23134
rect 438082 23218 438318 23454
rect 438082 22898 438318 23134
rect 442030 23218 442266 23454
rect 442030 22898 442266 23134
rect 452934 23218 453170 23454
rect 452934 22898 453170 23134
rect 453882 23218 454118 23454
rect 453882 22898 454118 23134
rect 454830 23218 455066 23454
rect 454830 22898 455066 23134
rect 463134 23218 463370 23454
rect 463134 22898 463370 23134
rect 467082 23218 467318 23454
rect 467082 22898 467318 23134
rect 471030 23218 471266 23454
rect 471030 22898 471266 23134
rect 481934 23218 482170 23454
rect 481934 22898 482170 23134
rect 482882 23218 483118 23454
rect 482882 22898 483118 23134
rect 483830 23218 484066 23454
rect 483830 22898 484066 23134
rect 492134 23218 492370 23454
rect 492134 22898 492370 23134
rect 496082 23218 496318 23454
rect 496082 22898 496318 23134
rect 500030 23218 500266 23454
rect 500030 22898 500266 23134
rect 510934 23218 511170 23454
rect 510934 22898 511170 23134
rect 511882 23218 512118 23454
rect 511882 22898 512118 23134
rect 512830 23218 513066 23454
rect 512830 22898 513066 23134
rect 521134 23218 521370 23454
rect 521134 22898 521370 23134
rect 525082 23218 525318 23454
rect 525082 22898 525318 23134
rect 542026 698218 542262 698454
rect 542346 698218 542582 698454
rect 542026 697898 542262 698134
rect 542346 697898 542582 698134
rect 542026 671218 542262 671454
rect 542346 671218 542582 671454
rect 542026 670898 542262 671134
rect 542346 670898 542582 671134
rect 542026 644218 542262 644454
rect 542346 644218 542582 644454
rect 542026 643898 542262 644134
rect 542346 643898 542582 644134
rect 542026 617218 542262 617454
rect 542346 617218 542582 617454
rect 542026 616898 542262 617134
rect 542346 616898 542582 617134
rect 542026 590218 542262 590454
rect 542346 590218 542582 590454
rect 542026 589898 542262 590134
rect 542346 589898 542582 590134
rect 542026 563218 542262 563454
rect 542346 563218 542582 563454
rect 542026 562898 542262 563134
rect 542346 562898 542582 563134
rect 542026 536218 542262 536454
rect 542346 536218 542582 536454
rect 542026 535898 542262 536134
rect 542346 535898 542582 536134
rect 542026 509218 542262 509454
rect 542346 509218 542582 509454
rect 542026 508898 542262 509134
rect 542346 508898 542582 509134
rect 542026 482218 542262 482454
rect 542346 482218 542582 482454
rect 542026 481898 542262 482134
rect 542346 481898 542582 482134
rect 542026 455218 542262 455454
rect 542346 455218 542582 455454
rect 542026 454898 542262 455134
rect 542346 454898 542582 455134
rect 542026 428218 542262 428454
rect 542346 428218 542582 428454
rect 542026 427898 542262 428134
rect 542346 427898 542582 428134
rect 542026 401218 542262 401454
rect 542346 401218 542582 401454
rect 542026 400898 542262 401134
rect 542346 400898 542582 401134
rect 542026 374218 542262 374454
rect 542346 374218 542582 374454
rect 542026 373898 542262 374134
rect 542346 373898 542582 374134
rect 542026 347218 542262 347454
rect 542346 347218 542582 347454
rect 542026 346898 542262 347134
rect 542346 346898 542582 347134
rect 542026 320218 542262 320454
rect 542346 320218 542582 320454
rect 542026 319898 542262 320134
rect 542346 319898 542582 320134
rect 542026 293218 542262 293454
rect 542346 293218 542582 293454
rect 542026 292898 542262 293134
rect 542346 292898 542582 293134
rect 542026 266218 542262 266454
rect 542346 266218 542582 266454
rect 542026 265898 542262 266134
rect 542346 265898 542582 266134
rect 542026 239218 542262 239454
rect 542346 239218 542582 239454
rect 542026 238898 542262 239134
rect 542346 238898 542582 239134
rect 542026 212218 542262 212454
rect 542346 212218 542582 212454
rect 542026 211898 542262 212134
rect 542346 211898 542582 212134
rect 542026 185218 542262 185454
rect 542346 185218 542582 185454
rect 542026 184898 542262 185134
rect 542346 184898 542582 185134
rect 542026 158218 542262 158454
rect 542346 158218 542582 158454
rect 542026 157898 542262 158134
rect 542346 157898 542582 158134
rect 542026 131218 542262 131454
rect 542346 131218 542582 131454
rect 542026 130898 542262 131134
rect 542346 130898 542582 131134
rect 542026 104218 542262 104454
rect 542346 104218 542582 104454
rect 542026 103898 542262 104134
rect 542346 103898 542582 104134
rect 542026 77218 542262 77454
rect 542346 77218 542582 77454
rect 542026 76898 542262 77134
rect 542346 76898 542582 77134
rect 545526 704602 545762 704838
rect 545846 704602 546082 704838
rect 545526 704282 545762 704518
rect 545846 704282 546082 704518
rect 545526 701593 545762 701829
rect 545846 701593 546082 701829
rect 545526 701273 545762 701509
rect 545846 701273 546082 701509
rect 570026 705562 570262 705798
rect 570346 705562 570582 705798
rect 570026 705242 570262 705478
rect 570346 705242 570582 705478
rect 545526 674593 545762 674829
rect 545846 674593 546082 674829
rect 545526 674273 545762 674509
rect 545846 674273 546082 674509
rect 545526 647593 545762 647829
rect 545846 647593 546082 647829
rect 545526 647273 545762 647509
rect 545846 647273 546082 647509
rect 545526 620593 545762 620829
rect 545846 620593 546082 620829
rect 545526 620273 545762 620509
rect 545846 620273 546082 620509
rect 545526 593593 545762 593829
rect 545846 593593 546082 593829
rect 545526 593273 545762 593509
rect 545846 593273 546082 593509
rect 545526 566593 545762 566829
rect 545846 566593 546082 566829
rect 545526 566273 545762 566509
rect 545846 566273 546082 566509
rect 545526 539593 545762 539829
rect 545846 539593 546082 539829
rect 545526 539273 545762 539509
rect 545846 539273 546082 539509
rect 545526 512593 545762 512829
rect 545846 512593 546082 512829
rect 545526 512273 545762 512509
rect 545846 512273 546082 512509
rect 545526 485593 545762 485829
rect 545846 485593 546082 485829
rect 545526 485273 545762 485509
rect 545846 485273 546082 485509
rect 545526 458593 545762 458829
rect 545846 458593 546082 458829
rect 545526 458273 545762 458509
rect 545846 458273 546082 458509
rect 545526 431593 545762 431829
rect 545846 431593 546082 431829
rect 545526 431273 545762 431509
rect 545846 431273 546082 431509
rect 545526 404593 545762 404829
rect 545846 404593 546082 404829
rect 545526 404273 545762 404509
rect 545846 404273 546082 404509
rect 545526 377593 545762 377829
rect 545846 377593 546082 377829
rect 545526 377273 545762 377509
rect 545846 377273 546082 377509
rect 545526 350593 545762 350829
rect 545846 350593 546082 350829
rect 545526 350273 545762 350509
rect 545846 350273 546082 350509
rect 545526 323593 545762 323829
rect 545846 323593 546082 323829
rect 545526 323273 545762 323509
rect 545846 323273 546082 323509
rect 545526 296593 545762 296829
rect 545846 296593 546082 296829
rect 545526 296273 545762 296509
rect 545846 296273 546082 296509
rect 545526 269593 545762 269829
rect 545846 269593 546082 269829
rect 545526 269273 545762 269509
rect 545846 269273 546082 269509
rect 545526 242593 545762 242829
rect 545846 242593 546082 242829
rect 545526 242273 545762 242509
rect 545846 242273 546082 242509
rect 545526 215593 545762 215829
rect 545846 215593 546082 215829
rect 545526 215273 545762 215509
rect 545846 215273 546082 215509
rect 545526 188593 545762 188829
rect 545846 188593 546082 188829
rect 545526 188273 545762 188509
rect 545846 188273 546082 188509
rect 545526 161593 545762 161829
rect 545846 161593 546082 161829
rect 545526 161273 545762 161509
rect 545846 161273 546082 161509
rect 545526 134593 545762 134829
rect 545846 134593 546082 134829
rect 545526 134273 545762 134509
rect 545846 134273 546082 134509
rect 545526 107593 545762 107829
rect 545846 107593 546082 107829
rect 545526 107273 545762 107509
rect 545846 107273 546082 107509
rect 545526 80593 545762 80829
rect 545846 80593 546082 80829
rect 545526 80273 545762 80509
rect 545846 80273 546082 80509
rect 532260 53593 532496 53829
rect 532260 53273 532496 53509
rect 533208 53593 533444 53829
rect 533208 53273 533444 53509
rect 534156 53593 534392 53829
rect 534156 53273 534392 53509
rect 535104 53593 535340 53829
rect 535104 53273 535340 53509
rect 540960 53593 541196 53829
rect 540960 53273 541196 53509
rect 544908 53593 545144 53829
rect 544908 53273 545144 53509
rect 548856 53593 549092 53829
rect 548856 53273 549092 53509
rect 552804 53593 553040 53829
rect 552804 53273 553040 53509
rect 532734 50218 532970 50454
rect 532734 49898 532970 50134
rect 533682 50218 533918 50454
rect 533682 49898 533918 50134
rect 534630 50218 534866 50454
rect 534630 49898 534866 50134
rect 542934 50218 543170 50454
rect 542934 49898 543170 50134
rect 546882 50218 547118 50454
rect 546882 49898 547118 50134
rect 550830 50218 551066 50454
rect 550830 49898 551066 50134
rect 531004 26593 531240 26829
rect 531004 26273 531240 26509
rect 539460 26593 539696 26829
rect 539460 26273 539696 26509
rect 540408 26593 540644 26829
rect 540408 26273 540644 26509
rect 541356 26593 541592 26829
rect 541356 26273 541592 26509
rect 542304 26593 542540 26829
rect 542304 26273 542540 26509
rect 548160 26593 548396 26829
rect 548160 26273 548396 26509
rect 552108 26593 552344 26829
rect 552108 26273 552344 26509
rect 556056 26593 556292 26829
rect 556056 26273 556292 26509
rect 529030 23218 529266 23454
rect 529030 22898 529266 23134
rect 539934 23218 540170 23454
rect 539934 22898 540170 23134
rect 540882 23218 541118 23454
rect 540882 22898 541118 23134
rect 541830 23218 542066 23454
rect 541830 22898 542066 23134
rect 550134 23218 550370 23454
rect 550134 22898 550370 23134
rect 554082 23218 554318 23454
rect 554082 22898 554318 23134
rect 558030 23218 558266 23454
rect 558030 22898 558266 23134
rect 570026 698218 570262 698454
rect 570346 698218 570582 698454
rect 570026 697898 570262 698134
rect 570346 697898 570582 698134
rect 570026 671218 570262 671454
rect 570346 671218 570582 671454
rect 570026 670898 570262 671134
rect 570346 670898 570582 671134
rect 570026 644218 570262 644454
rect 570346 644218 570582 644454
rect 570026 643898 570262 644134
rect 570346 643898 570582 644134
rect 570026 617218 570262 617454
rect 570346 617218 570582 617454
rect 570026 616898 570262 617134
rect 570346 616898 570582 617134
rect 570026 590218 570262 590454
rect 570346 590218 570582 590454
rect 570026 589898 570262 590134
rect 570346 589898 570582 590134
rect 570026 563218 570262 563454
rect 570346 563218 570582 563454
rect 570026 562898 570262 563134
rect 570346 562898 570582 563134
rect 570026 536218 570262 536454
rect 570346 536218 570582 536454
rect 570026 535898 570262 536134
rect 570346 535898 570582 536134
rect 570026 509218 570262 509454
rect 570346 509218 570582 509454
rect 570026 508898 570262 509134
rect 570346 508898 570582 509134
rect 570026 482218 570262 482454
rect 570346 482218 570582 482454
rect 570026 481898 570262 482134
rect 570346 481898 570582 482134
rect 570026 455218 570262 455454
rect 570346 455218 570582 455454
rect 570026 454898 570262 455134
rect 570346 454898 570582 455134
rect 570026 428218 570262 428454
rect 570346 428218 570582 428454
rect 570026 427898 570262 428134
rect 570346 427898 570582 428134
rect 570026 401218 570262 401454
rect 570346 401218 570582 401454
rect 570026 400898 570262 401134
rect 570346 400898 570582 401134
rect 570026 374218 570262 374454
rect 570346 374218 570582 374454
rect 570026 373898 570262 374134
rect 570346 373898 570582 374134
rect 570026 347218 570262 347454
rect 570346 347218 570582 347454
rect 570026 346898 570262 347134
rect 570346 346898 570582 347134
rect 570026 320218 570262 320454
rect 570346 320218 570582 320454
rect 570026 319898 570262 320134
rect 570346 319898 570582 320134
rect 570026 293218 570262 293454
rect 570346 293218 570582 293454
rect 570026 292898 570262 293134
rect 570346 292898 570582 293134
rect 570026 266218 570262 266454
rect 570346 266218 570582 266454
rect 570026 265898 570262 266134
rect 570346 265898 570582 266134
rect 570026 239218 570262 239454
rect 570346 239218 570582 239454
rect 570026 238898 570262 239134
rect 570346 238898 570582 239134
rect 570026 212218 570262 212454
rect 570346 212218 570582 212454
rect 570026 211898 570262 212134
rect 570346 211898 570582 212134
rect 570026 185218 570262 185454
rect 570346 185218 570582 185454
rect 570026 184898 570262 185134
rect 570346 184898 570582 185134
rect 570026 158218 570262 158454
rect 570346 158218 570582 158454
rect 570026 157898 570262 158134
rect 570346 157898 570582 158134
rect 570026 131218 570262 131454
rect 570346 131218 570582 131454
rect 570026 130898 570262 131134
rect 570346 130898 570582 131134
rect 570026 104218 570262 104454
rect 570346 104218 570582 104454
rect 570026 103898 570262 104134
rect 570346 103898 570582 104134
rect 570026 77218 570262 77454
rect 570346 77218 570582 77454
rect 570026 76898 570262 77134
rect 570346 76898 570582 77134
rect 561260 53593 561496 53829
rect 561260 53273 561496 53509
rect 562208 53593 562444 53829
rect 562208 53273 562444 53509
rect 563156 53593 563392 53829
rect 563156 53273 563392 53509
rect 564104 53593 564340 53829
rect 564104 53273 564340 53509
rect 561734 50218 561970 50454
rect 561734 49898 561970 50134
rect 562682 50218 562918 50454
rect 562682 49898 562918 50134
rect 563630 50218 563866 50454
rect 563630 49898 563866 50134
rect 570026 50218 570262 50454
rect 570346 50218 570582 50454
rect 570026 49898 570262 50134
rect 570346 49898 570582 50134
rect 560004 26593 560240 26829
rect 560004 26273 560240 26509
rect 570026 23218 570262 23454
rect 570346 23218 570582 23454
rect 570026 22898 570262 23134
rect 570346 22898 570582 23134
rect 69526 -582 69762 -346
rect 69846 -582 70082 -346
rect 69526 -902 69762 -666
rect 69846 -902 70082 -666
rect 570026 -1542 570262 -1306
rect 570346 -1542 570582 -1306
rect 570026 -1862 570262 -1626
rect 570346 -1862 570582 -1626
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 573526 704602 573762 704838
rect 573846 704602 574082 704838
rect 573526 704282 573762 704518
rect 573846 704282 574082 704518
rect 573526 701593 573762 701829
rect 573846 701593 574082 701829
rect 573526 701273 573762 701509
rect 573846 701273 574082 701509
rect 573526 674593 573762 674829
rect 573846 674593 574082 674829
rect 573526 674273 573762 674509
rect 573846 674273 574082 674509
rect 573526 647593 573762 647829
rect 573846 647593 574082 647829
rect 573526 647273 573762 647509
rect 573846 647273 574082 647509
rect 573526 620593 573762 620829
rect 573846 620593 574082 620829
rect 573526 620273 573762 620509
rect 573846 620273 574082 620509
rect 573526 593593 573762 593829
rect 573846 593593 574082 593829
rect 573526 593273 573762 593509
rect 573846 593273 574082 593509
rect 573526 566593 573762 566829
rect 573846 566593 574082 566829
rect 573526 566273 573762 566509
rect 573846 566273 574082 566509
rect 573526 539593 573762 539829
rect 573846 539593 574082 539829
rect 573526 539273 573762 539509
rect 573846 539273 574082 539509
rect 573526 512593 573762 512829
rect 573846 512593 574082 512829
rect 573526 512273 573762 512509
rect 573846 512273 574082 512509
rect 573526 485593 573762 485829
rect 573846 485593 574082 485829
rect 573526 485273 573762 485509
rect 573846 485273 574082 485509
rect 573526 458593 573762 458829
rect 573846 458593 574082 458829
rect 573526 458273 573762 458509
rect 573846 458273 574082 458509
rect 573526 431593 573762 431829
rect 573846 431593 574082 431829
rect 573526 431273 573762 431509
rect 573846 431273 574082 431509
rect 573526 404593 573762 404829
rect 573846 404593 574082 404829
rect 573526 404273 573762 404509
rect 573846 404273 574082 404509
rect 573526 377593 573762 377829
rect 573846 377593 574082 377829
rect 573526 377273 573762 377509
rect 573846 377273 574082 377509
rect 573526 350593 573762 350829
rect 573846 350593 574082 350829
rect 573526 350273 573762 350509
rect 573846 350273 574082 350509
rect 573526 323593 573762 323829
rect 573846 323593 574082 323829
rect 573526 323273 573762 323509
rect 573846 323273 574082 323509
rect 573526 296593 573762 296829
rect 573846 296593 574082 296829
rect 573526 296273 573762 296509
rect 573846 296273 574082 296509
rect 573526 269593 573762 269829
rect 573846 269593 574082 269829
rect 573526 269273 573762 269509
rect 573846 269273 574082 269509
rect 573526 242593 573762 242829
rect 573846 242593 574082 242829
rect 573526 242273 573762 242509
rect 573846 242273 574082 242509
rect 573526 215593 573762 215829
rect 573846 215593 574082 215829
rect 573526 215273 573762 215509
rect 573846 215273 574082 215509
rect 573526 188593 573762 188829
rect 573846 188593 574082 188829
rect 573526 188273 573762 188509
rect 573846 188273 574082 188509
rect 573526 161593 573762 161829
rect 573846 161593 574082 161829
rect 573526 161273 573762 161509
rect 573846 161273 574082 161509
rect 573526 134593 573762 134829
rect 573846 134593 574082 134829
rect 573526 134273 573762 134509
rect 573846 134273 574082 134509
rect 573526 107593 573762 107829
rect 573846 107593 574082 107829
rect 573526 107273 573762 107509
rect 573846 107273 574082 107509
rect 573526 80593 573762 80829
rect 573846 80593 574082 80829
rect 573526 80273 573762 80509
rect 573846 80273 574082 80509
rect 573526 53593 573762 53829
rect 573846 53593 574082 53829
rect 573526 53273 573762 53509
rect 573846 53273 574082 53509
rect 573526 26593 573762 26829
rect 573846 26593 574082 26829
rect 573526 26273 573762 26509
rect 573846 26273 574082 26509
rect 573526 -582 573762 -346
rect 573846 -582 574082 -346
rect 573526 -902 573762 -666
rect 573846 -902 574082 -666
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 701593 585578 701829
rect 585662 701593 585898 701829
rect 585342 701273 585578 701509
rect 585662 701273 585898 701509
rect 585342 674593 585578 674829
rect 585662 674593 585898 674829
rect 585342 674273 585578 674509
rect 585662 674273 585898 674509
rect 585342 647593 585578 647829
rect 585662 647593 585898 647829
rect 585342 647273 585578 647509
rect 585662 647273 585898 647509
rect 585342 620593 585578 620829
rect 585662 620593 585898 620829
rect 585342 620273 585578 620509
rect 585662 620273 585898 620509
rect 585342 593593 585578 593829
rect 585662 593593 585898 593829
rect 585342 593273 585578 593509
rect 585662 593273 585898 593509
rect 585342 566593 585578 566829
rect 585662 566593 585898 566829
rect 585342 566273 585578 566509
rect 585662 566273 585898 566509
rect 585342 539593 585578 539829
rect 585662 539593 585898 539829
rect 585342 539273 585578 539509
rect 585662 539273 585898 539509
rect 585342 512593 585578 512829
rect 585662 512593 585898 512829
rect 585342 512273 585578 512509
rect 585662 512273 585898 512509
rect 585342 485593 585578 485829
rect 585662 485593 585898 485829
rect 585342 485273 585578 485509
rect 585662 485273 585898 485509
rect 585342 458593 585578 458829
rect 585662 458593 585898 458829
rect 585342 458273 585578 458509
rect 585662 458273 585898 458509
rect 585342 431593 585578 431829
rect 585662 431593 585898 431829
rect 585342 431273 585578 431509
rect 585662 431273 585898 431509
rect 585342 404593 585578 404829
rect 585662 404593 585898 404829
rect 585342 404273 585578 404509
rect 585662 404273 585898 404509
rect 585342 377593 585578 377829
rect 585662 377593 585898 377829
rect 585342 377273 585578 377509
rect 585662 377273 585898 377509
rect 585342 350593 585578 350829
rect 585662 350593 585898 350829
rect 585342 350273 585578 350509
rect 585662 350273 585898 350509
rect 585342 323593 585578 323829
rect 585662 323593 585898 323829
rect 585342 323273 585578 323509
rect 585662 323273 585898 323509
rect 585342 296593 585578 296829
rect 585662 296593 585898 296829
rect 585342 296273 585578 296509
rect 585662 296273 585898 296509
rect 585342 269593 585578 269829
rect 585662 269593 585898 269829
rect 585342 269273 585578 269509
rect 585662 269273 585898 269509
rect 585342 242593 585578 242829
rect 585662 242593 585898 242829
rect 585342 242273 585578 242509
rect 585662 242273 585898 242509
rect 585342 215593 585578 215829
rect 585662 215593 585898 215829
rect 585342 215273 585578 215509
rect 585662 215273 585898 215509
rect 585342 188593 585578 188829
rect 585662 188593 585898 188829
rect 585342 188273 585578 188509
rect 585662 188273 585898 188509
rect 585342 161593 585578 161829
rect 585662 161593 585898 161829
rect 585342 161273 585578 161509
rect 585662 161273 585898 161509
rect 585342 134593 585578 134829
rect 585662 134593 585898 134829
rect 585342 134273 585578 134509
rect 585662 134273 585898 134509
rect 585342 107593 585578 107829
rect 585662 107593 585898 107829
rect 585342 107273 585578 107509
rect 585662 107273 585898 107509
rect 585342 80593 585578 80829
rect 585662 80593 585898 80829
rect 585342 80273 585578 80509
rect 585662 80273 585898 80509
rect 585342 53593 585578 53829
rect 585662 53593 585898 53829
rect 585342 53273 585578 53509
rect 585662 53273 585898 53509
rect 585342 26593 585578 26829
rect 585662 26593 585898 26829
rect 585342 26273 585578 26509
rect 585662 26273 585898 26509
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 698218 586538 698454
rect 586622 698218 586858 698454
rect 586302 697898 586538 698134
rect 586622 697898 586858 698134
rect 586302 671218 586538 671454
rect 586622 671218 586858 671454
rect 586302 670898 586538 671134
rect 586622 670898 586858 671134
rect 586302 644218 586538 644454
rect 586622 644218 586858 644454
rect 586302 643898 586538 644134
rect 586622 643898 586858 644134
rect 586302 617218 586538 617454
rect 586622 617218 586858 617454
rect 586302 616898 586538 617134
rect 586622 616898 586858 617134
rect 586302 590218 586538 590454
rect 586622 590218 586858 590454
rect 586302 589898 586538 590134
rect 586622 589898 586858 590134
rect 586302 563218 586538 563454
rect 586622 563218 586858 563454
rect 586302 562898 586538 563134
rect 586622 562898 586858 563134
rect 586302 536218 586538 536454
rect 586622 536218 586858 536454
rect 586302 535898 586538 536134
rect 586622 535898 586858 536134
rect 586302 509218 586538 509454
rect 586622 509218 586858 509454
rect 586302 508898 586538 509134
rect 586622 508898 586858 509134
rect 586302 482218 586538 482454
rect 586622 482218 586858 482454
rect 586302 481898 586538 482134
rect 586622 481898 586858 482134
rect 586302 455218 586538 455454
rect 586622 455218 586858 455454
rect 586302 454898 586538 455134
rect 586622 454898 586858 455134
rect 586302 428218 586538 428454
rect 586622 428218 586858 428454
rect 586302 427898 586538 428134
rect 586622 427898 586858 428134
rect 586302 401218 586538 401454
rect 586622 401218 586858 401454
rect 586302 400898 586538 401134
rect 586622 400898 586858 401134
rect 586302 374218 586538 374454
rect 586622 374218 586858 374454
rect 586302 373898 586538 374134
rect 586622 373898 586858 374134
rect 586302 347218 586538 347454
rect 586622 347218 586858 347454
rect 586302 346898 586538 347134
rect 586622 346898 586858 347134
rect 586302 320218 586538 320454
rect 586622 320218 586858 320454
rect 586302 319898 586538 320134
rect 586622 319898 586858 320134
rect 586302 293218 586538 293454
rect 586622 293218 586858 293454
rect 586302 292898 586538 293134
rect 586622 292898 586858 293134
rect 586302 266218 586538 266454
rect 586622 266218 586858 266454
rect 586302 265898 586538 266134
rect 586622 265898 586858 266134
rect 586302 239218 586538 239454
rect 586622 239218 586858 239454
rect 586302 238898 586538 239134
rect 586622 238898 586858 239134
rect 586302 212218 586538 212454
rect 586622 212218 586858 212454
rect 586302 211898 586538 212134
rect 586622 211898 586858 212134
rect 586302 185218 586538 185454
rect 586622 185218 586858 185454
rect 586302 184898 586538 185134
rect 586622 184898 586858 185134
rect 586302 158218 586538 158454
rect 586622 158218 586858 158454
rect 586302 157898 586538 158134
rect 586622 157898 586858 158134
rect 586302 131218 586538 131454
rect 586622 131218 586858 131454
rect 586302 130898 586538 131134
rect 586622 130898 586858 131134
rect 586302 104218 586538 104454
rect 586622 104218 586858 104454
rect 586302 103898 586538 104134
rect 586622 103898 586858 104134
rect 586302 77218 586538 77454
rect 586622 77218 586858 77454
rect 586302 76898 586538 77134
rect 586622 76898 586858 77134
rect 586302 50218 586538 50454
rect 586622 50218 586858 50454
rect 586302 49898 586538 50134
rect 586622 49898 586858 50134
rect 586302 23218 586538 23454
rect 586622 23218 586858 23454
rect 586302 22898 586538 23134
rect 586622 22898 586858 23134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 38026 705798
rect 38262 705562 38346 705798
rect 38582 705562 66026 705798
rect 66262 705562 66346 705798
rect 66582 705562 94026 705798
rect 94262 705562 94346 705798
rect 94582 705562 122026 705798
rect 122262 705562 122346 705798
rect 122582 705562 150026 705798
rect 150262 705562 150346 705798
rect 150582 705562 178026 705798
rect 178262 705562 178346 705798
rect 178582 705562 206026 705798
rect 206262 705562 206346 705798
rect 206582 705562 234026 705798
rect 234262 705562 234346 705798
rect 234582 705562 262026 705798
rect 262262 705562 262346 705798
rect 262582 705562 290026 705798
rect 290262 705562 290346 705798
rect 290582 705562 318026 705798
rect 318262 705562 318346 705798
rect 318582 705562 346026 705798
rect 346262 705562 346346 705798
rect 346582 705562 374026 705798
rect 374262 705562 374346 705798
rect 374582 705562 402026 705798
rect 402262 705562 402346 705798
rect 402582 705562 430026 705798
rect 430262 705562 430346 705798
rect 430582 705562 458026 705798
rect 458262 705562 458346 705798
rect 458582 705562 486026 705798
rect 486262 705562 486346 705798
rect 486582 705562 514026 705798
rect 514262 705562 514346 705798
rect 514582 705562 542026 705798
rect 542262 705562 542346 705798
rect 542582 705562 570026 705798
rect 570262 705562 570346 705798
rect 570582 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 38026 705478
rect 38262 705242 38346 705478
rect 38582 705242 66026 705478
rect 66262 705242 66346 705478
rect 66582 705242 94026 705478
rect 94262 705242 94346 705478
rect 94582 705242 122026 705478
rect 122262 705242 122346 705478
rect 122582 705242 150026 705478
rect 150262 705242 150346 705478
rect 150582 705242 178026 705478
rect 178262 705242 178346 705478
rect 178582 705242 206026 705478
rect 206262 705242 206346 705478
rect 206582 705242 234026 705478
rect 234262 705242 234346 705478
rect 234582 705242 262026 705478
rect 262262 705242 262346 705478
rect 262582 705242 290026 705478
rect 290262 705242 290346 705478
rect 290582 705242 318026 705478
rect 318262 705242 318346 705478
rect 318582 705242 346026 705478
rect 346262 705242 346346 705478
rect 346582 705242 374026 705478
rect 374262 705242 374346 705478
rect 374582 705242 402026 705478
rect 402262 705242 402346 705478
rect 402582 705242 430026 705478
rect 430262 705242 430346 705478
rect 430582 705242 458026 705478
rect 458262 705242 458346 705478
rect 458582 705242 486026 705478
rect 486262 705242 486346 705478
rect 486582 705242 514026 705478
rect 514262 705242 514346 705478
rect 514582 705242 542026 705478
rect 542262 705242 542346 705478
rect 542582 705242 570026 705478
rect 570262 705242 570346 705478
rect 570582 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 41526 704838
rect 41762 704602 41846 704838
rect 42082 704602 69526 704838
rect 69762 704602 69846 704838
rect 70082 704602 97526 704838
rect 97762 704602 97846 704838
rect 98082 704602 125526 704838
rect 125762 704602 125846 704838
rect 126082 704602 153526 704838
rect 153762 704602 153846 704838
rect 154082 704602 181526 704838
rect 181762 704602 181846 704838
rect 182082 704602 209526 704838
rect 209762 704602 209846 704838
rect 210082 704602 237526 704838
rect 237762 704602 237846 704838
rect 238082 704602 265526 704838
rect 265762 704602 265846 704838
rect 266082 704602 293526 704838
rect 293762 704602 293846 704838
rect 294082 704602 321526 704838
rect 321762 704602 321846 704838
rect 322082 704602 349526 704838
rect 349762 704602 349846 704838
rect 350082 704602 377526 704838
rect 377762 704602 377846 704838
rect 378082 704602 405526 704838
rect 405762 704602 405846 704838
rect 406082 704602 433526 704838
rect 433762 704602 433846 704838
rect 434082 704602 461526 704838
rect 461762 704602 461846 704838
rect 462082 704602 489526 704838
rect 489762 704602 489846 704838
rect 490082 704602 517526 704838
rect 517762 704602 517846 704838
rect 518082 704602 545526 704838
rect 545762 704602 545846 704838
rect 546082 704602 573526 704838
rect 573762 704602 573846 704838
rect 574082 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 41526 704518
rect 41762 704282 41846 704518
rect 42082 704282 69526 704518
rect 69762 704282 69846 704518
rect 70082 704282 97526 704518
rect 97762 704282 97846 704518
rect 98082 704282 125526 704518
rect 125762 704282 125846 704518
rect 126082 704282 153526 704518
rect 153762 704282 153846 704518
rect 154082 704282 181526 704518
rect 181762 704282 181846 704518
rect 182082 704282 209526 704518
rect 209762 704282 209846 704518
rect 210082 704282 237526 704518
rect 237762 704282 237846 704518
rect 238082 704282 265526 704518
rect 265762 704282 265846 704518
rect 266082 704282 293526 704518
rect 293762 704282 293846 704518
rect 294082 704282 321526 704518
rect 321762 704282 321846 704518
rect 322082 704282 349526 704518
rect 349762 704282 349846 704518
rect 350082 704282 377526 704518
rect 377762 704282 377846 704518
rect 378082 704282 405526 704518
rect 405762 704282 405846 704518
rect 406082 704282 433526 704518
rect 433762 704282 433846 704518
rect 434082 704282 461526 704518
rect 461762 704282 461846 704518
rect 462082 704282 489526 704518
rect 489762 704282 489846 704518
rect 490082 704282 517526 704518
rect 517762 704282 517846 704518
rect 518082 704282 545526 704518
rect 545762 704282 545846 704518
rect 546082 704282 573526 704518
rect 573762 704282 573846 704518
rect 574082 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 701829 592650 701861
rect -8726 701593 -1974 701829
rect -1738 701593 -1654 701829
rect -1418 701593 41526 701829
rect 41762 701593 41846 701829
rect 42082 701593 69526 701829
rect 69762 701593 69846 701829
rect 70082 701593 97526 701829
rect 97762 701593 97846 701829
rect 98082 701593 125526 701829
rect 125762 701593 125846 701829
rect 126082 701593 153526 701829
rect 153762 701593 153846 701829
rect 154082 701593 181526 701829
rect 181762 701593 181846 701829
rect 182082 701593 209526 701829
rect 209762 701593 209846 701829
rect 210082 701593 237526 701829
rect 237762 701593 237846 701829
rect 238082 701593 265526 701829
rect 265762 701593 265846 701829
rect 266082 701593 293526 701829
rect 293762 701593 293846 701829
rect 294082 701593 321526 701829
rect 321762 701593 321846 701829
rect 322082 701593 349526 701829
rect 349762 701593 349846 701829
rect 350082 701593 377526 701829
rect 377762 701593 377846 701829
rect 378082 701593 405526 701829
rect 405762 701593 405846 701829
rect 406082 701593 433526 701829
rect 433762 701593 433846 701829
rect 434082 701593 461526 701829
rect 461762 701593 461846 701829
rect 462082 701593 489526 701829
rect 489762 701593 489846 701829
rect 490082 701593 517526 701829
rect 517762 701593 517846 701829
rect 518082 701593 545526 701829
rect 545762 701593 545846 701829
rect 546082 701593 573526 701829
rect 573762 701593 573846 701829
rect 574082 701593 585342 701829
rect 585578 701593 585662 701829
rect 585898 701593 592650 701829
rect -8726 701509 592650 701593
rect -8726 701273 -1974 701509
rect -1738 701273 -1654 701509
rect -1418 701273 41526 701509
rect 41762 701273 41846 701509
rect 42082 701273 69526 701509
rect 69762 701273 69846 701509
rect 70082 701273 97526 701509
rect 97762 701273 97846 701509
rect 98082 701273 125526 701509
rect 125762 701273 125846 701509
rect 126082 701273 153526 701509
rect 153762 701273 153846 701509
rect 154082 701273 181526 701509
rect 181762 701273 181846 701509
rect 182082 701273 209526 701509
rect 209762 701273 209846 701509
rect 210082 701273 237526 701509
rect 237762 701273 237846 701509
rect 238082 701273 265526 701509
rect 265762 701273 265846 701509
rect 266082 701273 293526 701509
rect 293762 701273 293846 701509
rect 294082 701273 321526 701509
rect 321762 701273 321846 701509
rect 322082 701273 349526 701509
rect 349762 701273 349846 701509
rect 350082 701273 377526 701509
rect 377762 701273 377846 701509
rect 378082 701273 405526 701509
rect 405762 701273 405846 701509
rect 406082 701273 433526 701509
rect 433762 701273 433846 701509
rect 434082 701273 461526 701509
rect 461762 701273 461846 701509
rect 462082 701273 489526 701509
rect 489762 701273 489846 701509
rect 490082 701273 517526 701509
rect 517762 701273 517846 701509
rect 518082 701273 545526 701509
rect 545762 701273 545846 701509
rect 546082 701273 573526 701509
rect 573762 701273 573846 701509
rect 574082 701273 585342 701509
rect 585578 701273 585662 701509
rect 585898 701273 592650 701509
rect -8726 701241 592650 701273
rect -8726 698454 592650 698486
rect -8726 698218 -2934 698454
rect -2698 698218 -2614 698454
rect -2378 698218 38026 698454
rect 38262 698218 38346 698454
rect 38582 698218 66026 698454
rect 66262 698218 66346 698454
rect 66582 698218 94026 698454
rect 94262 698218 94346 698454
rect 94582 698218 122026 698454
rect 122262 698218 122346 698454
rect 122582 698218 150026 698454
rect 150262 698218 150346 698454
rect 150582 698218 178026 698454
rect 178262 698218 178346 698454
rect 178582 698218 206026 698454
rect 206262 698218 206346 698454
rect 206582 698218 234026 698454
rect 234262 698218 234346 698454
rect 234582 698218 262026 698454
rect 262262 698218 262346 698454
rect 262582 698218 290026 698454
rect 290262 698218 290346 698454
rect 290582 698218 318026 698454
rect 318262 698218 318346 698454
rect 318582 698218 346026 698454
rect 346262 698218 346346 698454
rect 346582 698218 374026 698454
rect 374262 698218 374346 698454
rect 374582 698218 402026 698454
rect 402262 698218 402346 698454
rect 402582 698218 430026 698454
rect 430262 698218 430346 698454
rect 430582 698218 458026 698454
rect 458262 698218 458346 698454
rect 458582 698218 486026 698454
rect 486262 698218 486346 698454
rect 486582 698218 514026 698454
rect 514262 698218 514346 698454
rect 514582 698218 542026 698454
rect 542262 698218 542346 698454
rect 542582 698218 570026 698454
rect 570262 698218 570346 698454
rect 570582 698218 586302 698454
rect 586538 698218 586622 698454
rect 586858 698218 592650 698454
rect -8726 698134 592650 698218
rect -8726 697898 -2934 698134
rect -2698 697898 -2614 698134
rect -2378 697898 38026 698134
rect 38262 697898 38346 698134
rect 38582 697898 66026 698134
rect 66262 697898 66346 698134
rect 66582 697898 94026 698134
rect 94262 697898 94346 698134
rect 94582 697898 122026 698134
rect 122262 697898 122346 698134
rect 122582 697898 150026 698134
rect 150262 697898 150346 698134
rect 150582 697898 178026 698134
rect 178262 697898 178346 698134
rect 178582 697898 206026 698134
rect 206262 697898 206346 698134
rect 206582 697898 234026 698134
rect 234262 697898 234346 698134
rect 234582 697898 262026 698134
rect 262262 697898 262346 698134
rect 262582 697898 290026 698134
rect 290262 697898 290346 698134
rect 290582 697898 318026 698134
rect 318262 697898 318346 698134
rect 318582 697898 346026 698134
rect 346262 697898 346346 698134
rect 346582 697898 374026 698134
rect 374262 697898 374346 698134
rect 374582 697898 402026 698134
rect 402262 697898 402346 698134
rect 402582 697898 430026 698134
rect 430262 697898 430346 698134
rect 430582 697898 458026 698134
rect 458262 697898 458346 698134
rect 458582 697898 486026 698134
rect 486262 697898 486346 698134
rect 486582 697898 514026 698134
rect 514262 697898 514346 698134
rect 514582 697898 542026 698134
rect 542262 697898 542346 698134
rect 542582 697898 570026 698134
rect 570262 697898 570346 698134
rect 570582 697898 586302 698134
rect 586538 697898 586622 698134
rect 586858 697898 592650 698134
rect -8726 697866 592650 697898
rect -8726 674829 592650 674861
rect -8726 674593 -1974 674829
rect -1738 674593 -1654 674829
rect -1418 674593 41526 674829
rect 41762 674593 41846 674829
rect 42082 674593 69526 674829
rect 69762 674593 69846 674829
rect 70082 674593 97526 674829
rect 97762 674593 97846 674829
rect 98082 674593 125526 674829
rect 125762 674593 125846 674829
rect 126082 674593 153526 674829
rect 153762 674593 153846 674829
rect 154082 674593 181526 674829
rect 181762 674593 181846 674829
rect 182082 674593 209526 674829
rect 209762 674593 209846 674829
rect 210082 674593 237526 674829
rect 237762 674593 237846 674829
rect 238082 674593 265526 674829
rect 265762 674593 265846 674829
rect 266082 674593 293526 674829
rect 293762 674593 293846 674829
rect 294082 674593 321526 674829
rect 321762 674593 321846 674829
rect 322082 674593 349526 674829
rect 349762 674593 349846 674829
rect 350082 674593 377526 674829
rect 377762 674593 377846 674829
rect 378082 674593 405526 674829
rect 405762 674593 405846 674829
rect 406082 674593 433526 674829
rect 433762 674593 433846 674829
rect 434082 674593 461526 674829
rect 461762 674593 461846 674829
rect 462082 674593 489526 674829
rect 489762 674593 489846 674829
rect 490082 674593 517526 674829
rect 517762 674593 517846 674829
rect 518082 674593 545526 674829
rect 545762 674593 545846 674829
rect 546082 674593 573526 674829
rect 573762 674593 573846 674829
rect 574082 674593 585342 674829
rect 585578 674593 585662 674829
rect 585898 674593 592650 674829
rect -8726 674509 592650 674593
rect -8726 674273 -1974 674509
rect -1738 674273 -1654 674509
rect -1418 674273 41526 674509
rect 41762 674273 41846 674509
rect 42082 674273 69526 674509
rect 69762 674273 69846 674509
rect 70082 674273 97526 674509
rect 97762 674273 97846 674509
rect 98082 674273 125526 674509
rect 125762 674273 125846 674509
rect 126082 674273 153526 674509
rect 153762 674273 153846 674509
rect 154082 674273 181526 674509
rect 181762 674273 181846 674509
rect 182082 674273 209526 674509
rect 209762 674273 209846 674509
rect 210082 674273 237526 674509
rect 237762 674273 237846 674509
rect 238082 674273 265526 674509
rect 265762 674273 265846 674509
rect 266082 674273 293526 674509
rect 293762 674273 293846 674509
rect 294082 674273 321526 674509
rect 321762 674273 321846 674509
rect 322082 674273 349526 674509
rect 349762 674273 349846 674509
rect 350082 674273 377526 674509
rect 377762 674273 377846 674509
rect 378082 674273 405526 674509
rect 405762 674273 405846 674509
rect 406082 674273 433526 674509
rect 433762 674273 433846 674509
rect 434082 674273 461526 674509
rect 461762 674273 461846 674509
rect 462082 674273 489526 674509
rect 489762 674273 489846 674509
rect 490082 674273 517526 674509
rect 517762 674273 517846 674509
rect 518082 674273 545526 674509
rect 545762 674273 545846 674509
rect 546082 674273 573526 674509
rect 573762 674273 573846 674509
rect 574082 674273 585342 674509
rect 585578 674273 585662 674509
rect 585898 674273 592650 674509
rect -8726 674241 592650 674273
rect -8726 671454 592650 671486
rect -8726 671218 -2934 671454
rect -2698 671218 -2614 671454
rect -2378 671218 38026 671454
rect 38262 671218 38346 671454
rect 38582 671218 66026 671454
rect 66262 671218 66346 671454
rect 66582 671218 94026 671454
rect 94262 671218 94346 671454
rect 94582 671218 122026 671454
rect 122262 671218 122346 671454
rect 122582 671218 150026 671454
rect 150262 671218 150346 671454
rect 150582 671218 178026 671454
rect 178262 671218 178346 671454
rect 178582 671218 206026 671454
rect 206262 671218 206346 671454
rect 206582 671218 234026 671454
rect 234262 671218 234346 671454
rect 234582 671218 262026 671454
rect 262262 671218 262346 671454
rect 262582 671218 290026 671454
rect 290262 671218 290346 671454
rect 290582 671218 318026 671454
rect 318262 671218 318346 671454
rect 318582 671218 346026 671454
rect 346262 671218 346346 671454
rect 346582 671218 374026 671454
rect 374262 671218 374346 671454
rect 374582 671218 402026 671454
rect 402262 671218 402346 671454
rect 402582 671218 430026 671454
rect 430262 671218 430346 671454
rect 430582 671218 458026 671454
rect 458262 671218 458346 671454
rect 458582 671218 486026 671454
rect 486262 671218 486346 671454
rect 486582 671218 514026 671454
rect 514262 671218 514346 671454
rect 514582 671218 542026 671454
rect 542262 671218 542346 671454
rect 542582 671218 570026 671454
rect 570262 671218 570346 671454
rect 570582 671218 586302 671454
rect 586538 671218 586622 671454
rect 586858 671218 592650 671454
rect -8726 671134 592650 671218
rect -8726 670898 -2934 671134
rect -2698 670898 -2614 671134
rect -2378 670898 38026 671134
rect 38262 670898 38346 671134
rect 38582 670898 66026 671134
rect 66262 670898 66346 671134
rect 66582 670898 94026 671134
rect 94262 670898 94346 671134
rect 94582 670898 122026 671134
rect 122262 670898 122346 671134
rect 122582 670898 150026 671134
rect 150262 670898 150346 671134
rect 150582 670898 178026 671134
rect 178262 670898 178346 671134
rect 178582 670898 206026 671134
rect 206262 670898 206346 671134
rect 206582 670898 234026 671134
rect 234262 670898 234346 671134
rect 234582 670898 262026 671134
rect 262262 670898 262346 671134
rect 262582 670898 290026 671134
rect 290262 670898 290346 671134
rect 290582 670898 318026 671134
rect 318262 670898 318346 671134
rect 318582 670898 346026 671134
rect 346262 670898 346346 671134
rect 346582 670898 374026 671134
rect 374262 670898 374346 671134
rect 374582 670898 402026 671134
rect 402262 670898 402346 671134
rect 402582 670898 430026 671134
rect 430262 670898 430346 671134
rect 430582 670898 458026 671134
rect 458262 670898 458346 671134
rect 458582 670898 486026 671134
rect 486262 670898 486346 671134
rect 486582 670898 514026 671134
rect 514262 670898 514346 671134
rect 514582 670898 542026 671134
rect 542262 670898 542346 671134
rect 542582 670898 570026 671134
rect 570262 670898 570346 671134
rect 570582 670898 586302 671134
rect 586538 670898 586622 671134
rect 586858 670898 592650 671134
rect -8726 670866 592650 670898
rect -8726 647829 592650 647861
rect -8726 647593 -1974 647829
rect -1738 647593 -1654 647829
rect -1418 647593 41526 647829
rect 41762 647593 41846 647829
rect 42082 647593 69526 647829
rect 69762 647593 69846 647829
rect 70082 647593 97526 647829
rect 97762 647593 97846 647829
rect 98082 647593 125526 647829
rect 125762 647593 125846 647829
rect 126082 647593 153526 647829
rect 153762 647593 153846 647829
rect 154082 647593 181526 647829
rect 181762 647593 181846 647829
rect 182082 647593 209526 647829
rect 209762 647593 209846 647829
rect 210082 647593 237526 647829
rect 237762 647593 237846 647829
rect 238082 647593 265526 647829
rect 265762 647593 265846 647829
rect 266082 647593 293526 647829
rect 293762 647593 293846 647829
rect 294082 647593 321526 647829
rect 321762 647593 321846 647829
rect 322082 647593 349526 647829
rect 349762 647593 349846 647829
rect 350082 647593 377526 647829
rect 377762 647593 377846 647829
rect 378082 647593 405526 647829
rect 405762 647593 405846 647829
rect 406082 647593 433526 647829
rect 433762 647593 433846 647829
rect 434082 647593 461526 647829
rect 461762 647593 461846 647829
rect 462082 647593 489526 647829
rect 489762 647593 489846 647829
rect 490082 647593 517526 647829
rect 517762 647593 517846 647829
rect 518082 647593 545526 647829
rect 545762 647593 545846 647829
rect 546082 647593 573526 647829
rect 573762 647593 573846 647829
rect 574082 647593 585342 647829
rect 585578 647593 585662 647829
rect 585898 647593 592650 647829
rect -8726 647509 592650 647593
rect -8726 647273 -1974 647509
rect -1738 647273 -1654 647509
rect -1418 647273 41526 647509
rect 41762 647273 41846 647509
rect 42082 647273 69526 647509
rect 69762 647273 69846 647509
rect 70082 647273 97526 647509
rect 97762 647273 97846 647509
rect 98082 647273 125526 647509
rect 125762 647273 125846 647509
rect 126082 647273 153526 647509
rect 153762 647273 153846 647509
rect 154082 647273 181526 647509
rect 181762 647273 181846 647509
rect 182082 647273 209526 647509
rect 209762 647273 209846 647509
rect 210082 647273 237526 647509
rect 237762 647273 237846 647509
rect 238082 647273 265526 647509
rect 265762 647273 265846 647509
rect 266082 647273 293526 647509
rect 293762 647273 293846 647509
rect 294082 647273 321526 647509
rect 321762 647273 321846 647509
rect 322082 647273 349526 647509
rect 349762 647273 349846 647509
rect 350082 647273 377526 647509
rect 377762 647273 377846 647509
rect 378082 647273 405526 647509
rect 405762 647273 405846 647509
rect 406082 647273 433526 647509
rect 433762 647273 433846 647509
rect 434082 647273 461526 647509
rect 461762 647273 461846 647509
rect 462082 647273 489526 647509
rect 489762 647273 489846 647509
rect 490082 647273 517526 647509
rect 517762 647273 517846 647509
rect 518082 647273 545526 647509
rect 545762 647273 545846 647509
rect 546082 647273 573526 647509
rect 573762 647273 573846 647509
rect 574082 647273 585342 647509
rect 585578 647273 585662 647509
rect 585898 647273 592650 647509
rect -8726 647241 592650 647273
rect -8726 644454 592650 644486
rect -8726 644218 -2934 644454
rect -2698 644218 -2614 644454
rect -2378 644218 38026 644454
rect 38262 644218 38346 644454
rect 38582 644218 66026 644454
rect 66262 644218 66346 644454
rect 66582 644218 94026 644454
rect 94262 644218 94346 644454
rect 94582 644218 122026 644454
rect 122262 644218 122346 644454
rect 122582 644218 150026 644454
rect 150262 644218 150346 644454
rect 150582 644218 178026 644454
rect 178262 644218 178346 644454
rect 178582 644218 206026 644454
rect 206262 644218 206346 644454
rect 206582 644218 234026 644454
rect 234262 644218 234346 644454
rect 234582 644218 262026 644454
rect 262262 644218 262346 644454
rect 262582 644218 290026 644454
rect 290262 644218 290346 644454
rect 290582 644218 318026 644454
rect 318262 644218 318346 644454
rect 318582 644218 346026 644454
rect 346262 644218 346346 644454
rect 346582 644218 374026 644454
rect 374262 644218 374346 644454
rect 374582 644218 402026 644454
rect 402262 644218 402346 644454
rect 402582 644218 430026 644454
rect 430262 644218 430346 644454
rect 430582 644218 458026 644454
rect 458262 644218 458346 644454
rect 458582 644218 486026 644454
rect 486262 644218 486346 644454
rect 486582 644218 514026 644454
rect 514262 644218 514346 644454
rect 514582 644218 542026 644454
rect 542262 644218 542346 644454
rect 542582 644218 570026 644454
rect 570262 644218 570346 644454
rect 570582 644218 586302 644454
rect 586538 644218 586622 644454
rect 586858 644218 592650 644454
rect -8726 644134 592650 644218
rect -8726 643898 -2934 644134
rect -2698 643898 -2614 644134
rect -2378 643898 38026 644134
rect 38262 643898 38346 644134
rect 38582 643898 66026 644134
rect 66262 643898 66346 644134
rect 66582 643898 94026 644134
rect 94262 643898 94346 644134
rect 94582 643898 122026 644134
rect 122262 643898 122346 644134
rect 122582 643898 150026 644134
rect 150262 643898 150346 644134
rect 150582 643898 178026 644134
rect 178262 643898 178346 644134
rect 178582 643898 206026 644134
rect 206262 643898 206346 644134
rect 206582 643898 234026 644134
rect 234262 643898 234346 644134
rect 234582 643898 262026 644134
rect 262262 643898 262346 644134
rect 262582 643898 290026 644134
rect 290262 643898 290346 644134
rect 290582 643898 318026 644134
rect 318262 643898 318346 644134
rect 318582 643898 346026 644134
rect 346262 643898 346346 644134
rect 346582 643898 374026 644134
rect 374262 643898 374346 644134
rect 374582 643898 402026 644134
rect 402262 643898 402346 644134
rect 402582 643898 430026 644134
rect 430262 643898 430346 644134
rect 430582 643898 458026 644134
rect 458262 643898 458346 644134
rect 458582 643898 486026 644134
rect 486262 643898 486346 644134
rect 486582 643898 514026 644134
rect 514262 643898 514346 644134
rect 514582 643898 542026 644134
rect 542262 643898 542346 644134
rect 542582 643898 570026 644134
rect 570262 643898 570346 644134
rect 570582 643898 586302 644134
rect 586538 643898 586622 644134
rect 586858 643898 592650 644134
rect -8726 643866 592650 643898
rect -8726 620829 592650 620861
rect -8726 620593 -1974 620829
rect -1738 620593 -1654 620829
rect -1418 620593 41526 620829
rect 41762 620593 41846 620829
rect 42082 620593 69526 620829
rect 69762 620593 69846 620829
rect 70082 620593 97526 620829
rect 97762 620593 97846 620829
rect 98082 620593 125526 620829
rect 125762 620593 125846 620829
rect 126082 620593 153526 620829
rect 153762 620593 153846 620829
rect 154082 620593 181526 620829
rect 181762 620593 181846 620829
rect 182082 620593 209526 620829
rect 209762 620593 209846 620829
rect 210082 620593 237526 620829
rect 237762 620593 237846 620829
rect 238082 620593 265526 620829
rect 265762 620593 265846 620829
rect 266082 620593 293526 620829
rect 293762 620593 293846 620829
rect 294082 620593 321526 620829
rect 321762 620593 321846 620829
rect 322082 620593 349526 620829
rect 349762 620593 349846 620829
rect 350082 620593 377526 620829
rect 377762 620593 377846 620829
rect 378082 620593 405526 620829
rect 405762 620593 405846 620829
rect 406082 620593 433526 620829
rect 433762 620593 433846 620829
rect 434082 620593 461526 620829
rect 461762 620593 461846 620829
rect 462082 620593 489526 620829
rect 489762 620593 489846 620829
rect 490082 620593 517526 620829
rect 517762 620593 517846 620829
rect 518082 620593 545526 620829
rect 545762 620593 545846 620829
rect 546082 620593 573526 620829
rect 573762 620593 573846 620829
rect 574082 620593 585342 620829
rect 585578 620593 585662 620829
rect 585898 620593 592650 620829
rect -8726 620509 592650 620593
rect -8726 620273 -1974 620509
rect -1738 620273 -1654 620509
rect -1418 620273 41526 620509
rect 41762 620273 41846 620509
rect 42082 620273 69526 620509
rect 69762 620273 69846 620509
rect 70082 620273 97526 620509
rect 97762 620273 97846 620509
rect 98082 620273 125526 620509
rect 125762 620273 125846 620509
rect 126082 620273 153526 620509
rect 153762 620273 153846 620509
rect 154082 620273 181526 620509
rect 181762 620273 181846 620509
rect 182082 620273 209526 620509
rect 209762 620273 209846 620509
rect 210082 620273 237526 620509
rect 237762 620273 237846 620509
rect 238082 620273 265526 620509
rect 265762 620273 265846 620509
rect 266082 620273 293526 620509
rect 293762 620273 293846 620509
rect 294082 620273 321526 620509
rect 321762 620273 321846 620509
rect 322082 620273 349526 620509
rect 349762 620273 349846 620509
rect 350082 620273 377526 620509
rect 377762 620273 377846 620509
rect 378082 620273 405526 620509
rect 405762 620273 405846 620509
rect 406082 620273 433526 620509
rect 433762 620273 433846 620509
rect 434082 620273 461526 620509
rect 461762 620273 461846 620509
rect 462082 620273 489526 620509
rect 489762 620273 489846 620509
rect 490082 620273 517526 620509
rect 517762 620273 517846 620509
rect 518082 620273 545526 620509
rect 545762 620273 545846 620509
rect 546082 620273 573526 620509
rect 573762 620273 573846 620509
rect 574082 620273 585342 620509
rect 585578 620273 585662 620509
rect 585898 620273 592650 620509
rect -8726 620241 592650 620273
rect -8726 617454 592650 617486
rect -8726 617218 -2934 617454
rect -2698 617218 -2614 617454
rect -2378 617218 38026 617454
rect 38262 617218 38346 617454
rect 38582 617218 66026 617454
rect 66262 617218 66346 617454
rect 66582 617218 94026 617454
rect 94262 617218 94346 617454
rect 94582 617218 122026 617454
rect 122262 617218 122346 617454
rect 122582 617218 150026 617454
rect 150262 617218 150346 617454
rect 150582 617218 178026 617454
rect 178262 617218 178346 617454
rect 178582 617218 206026 617454
rect 206262 617218 206346 617454
rect 206582 617218 234026 617454
rect 234262 617218 234346 617454
rect 234582 617218 262026 617454
rect 262262 617218 262346 617454
rect 262582 617218 290026 617454
rect 290262 617218 290346 617454
rect 290582 617218 318026 617454
rect 318262 617218 318346 617454
rect 318582 617218 346026 617454
rect 346262 617218 346346 617454
rect 346582 617218 374026 617454
rect 374262 617218 374346 617454
rect 374582 617218 402026 617454
rect 402262 617218 402346 617454
rect 402582 617218 430026 617454
rect 430262 617218 430346 617454
rect 430582 617218 458026 617454
rect 458262 617218 458346 617454
rect 458582 617218 486026 617454
rect 486262 617218 486346 617454
rect 486582 617218 514026 617454
rect 514262 617218 514346 617454
rect 514582 617218 542026 617454
rect 542262 617218 542346 617454
rect 542582 617218 570026 617454
rect 570262 617218 570346 617454
rect 570582 617218 586302 617454
rect 586538 617218 586622 617454
rect 586858 617218 592650 617454
rect -8726 617134 592650 617218
rect -8726 616898 -2934 617134
rect -2698 616898 -2614 617134
rect -2378 616898 38026 617134
rect 38262 616898 38346 617134
rect 38582 616898 66026 617134
rect 66262 616898 66346 617134
rect 66582 616898 94026 617134
rect 94262 616898 94346 617134
rect 94582 616898 122026 617134
rect 122262 616898 122346 617134
rect 122582 616898 150026 617134
rect 150262 616898 150346 617134
rect 150582 616898 178026 617134
rect 178262 616898 178346 617134
rect 178582 616898 206026 617134
rect 206262 616898 206346 617134
rect 206582 616898 234026 617134
rect 234262 616898 234346 617134
rect 234582 616898 262026 617134
rect 262262 616898 262346 617134
rect 262582 616898 290026 617134
rect 290262 616898 290346 617134
rect 290582 616898 318026 617134
rect 318262 616898 318346 617134
rect 318582 616898 346026 617134
rect 346262 616898 346346 617134
rect 346582 616898 374026 617134
rect 374262 616898 374346 617134
rect 374582 616898 402026 617134
rect 402262 616898 402346 617134
rect 402582 616898 430026 617134
rect 430262 616898 430346 617134
rect 430582 616898 458026 617134
rect 458262 616898 458346 617134
rect 458582 616898 486026 617134
rect 486262 616898 486346 617134
rect 486582 616898 514026 617134
rect 514262 616898 514346 617134
rect 514582 616898 542026 617134
rect 542262 616898 542346 617134
rect 542582 616898 570026 617134
rect 570262 616898 570346 617134
rect 570582 616898 586302 617134
rect 586538 616898 586622 617134
rect 586858 616898 592650 617134
rect -8726 616866 592650 616898
rect -8726 593829 592650 593861
rect -8726 593593 -1974 593829
rect -1738 593593 -1654 593829
rect -1418 593593 41526 593829
rect 41762 593593 41846 593829
rect 42082 593593 69526 593829
rect 69762 593593 69846 593829
rect 70082 593593 97526 593829
rect 97762 593593 97846 593829
rect 98082 593593 125526 593829
rect 125762 593593 125846 593829
rect 126082 593593 153526 593829
rect 153762 593593 153846 593829
rect 154082 593593 181526 593829
rect 181762 593593 181846 593829
rect 182082 593593 209526 593829
rect 209762 593593 209846 593829
rect 210082 593593 237526 593829
rect 237762 593593 237846 593829
rect 238082 593593 265526 593829
rect 265762 593593 265846 593829
rect 266082 593593 293526 593829
rect 293762 593593 293846 593829
rect 294082 593593 321526 593829
rect 321762 593593 321846 593829
rect 322082 593593 349526 593829
rect 349762 593593 349846 593829
rect 350082 593593 377526 593829
rect 377762 593593 377846 593829
rect 378082 593593 405526 593829
rect 405762 593593 405846 593829
rect 406082 593593 433526 593829
rect 433762 593593 433846 593829
rect 434082 593593 461526 593829
rect 461762 593593 461846 593829
rect 462082 593593 489526 593829
rect 489762 593593 489846 593829
rect 490082 593593 517526 593829
rect 517762 593593 517846 593829
rect 518082 593593 545526 593829
rect 545762 593593 545846 593829
rect 546082 593593 573526 593829
rect 573762 593593 573846 593829
rect 574082 593593 585342 593829
rect 585578 593593 585662 593829
rect 585898 593593 592650 593829
rect -8726 593509 592650 593593
rect -8726 593273 -1974 593509
rect -1738 593273 -1654 593509
rect -1418 593273 41526 593509
rect 41762 593273 41846 593509
rect 42082 593273 69526 593509
rect 69762 593273 69846 593509
rect 70082 593273 97526 593509
rect 97762 593273 97846 593509
rect 98082 593273 125526 593509
rect 125762 593273 125846 593509
rect 126082 593273 153526 593509
rect 153762 593273 153846 593509
rect 154082 593273 181526 593509
rect 181762 593273 181846 593509
rect 182082 593273 209526 593509
rect 209762 593273 209846 593509
rect 210082 593273 237526 593509
rect 237762 593273 237846 593509
rect 238082 593273 265526 593509
rect 265762 593273 265846 593509
rect 266082 593273 293526 593509
rect 293762 593273 293846 593509
rect 294082 593273 321526 593509
rect 321762 593273 321846 593509
rect 322082 593273 349526 593509
rect 349762 593273 349846 593509
rect 350082 593273 377526 593509
rect 377762 593273 377846 593509
rect 378082 593273 405526 593509
rect 405762 593273 405846 593509
rect 406082 593273 433526 593509
rect 433762 593273 433846 593509
rect 434082 593273 461526 593509
rect 461762 593273 461846 593509
rect 462082 593273 489526 593509
rect 489762 593273 489846 593509
rect 490082 593273 517526 593509
rect 517762 593273 517846 593509
rect 518082 593273 545526 593509
rect 545762 593273 545846 593509
rect 546082 593273 573526 593509
rect 573762 593273 573846 593509
rect 574082 593273 585342 593509
rect 585578 593273 585662 593509
rect 585898 593273 592650 593509
rect -8726 593241 592650 593273
rect -8726 590454 592650 590486
rect -8726 590218 -2934 590454
rect -2698 590218 -2614 590454
rect -2378 590218 38026 590454
rect 38262 590218 38346 590454
rect 38582 590218 66026 590454
rect 66262 590218 66346 590454
rect 66582 590218 94026 590454
rect 94262 590218 94346 590454
rect 94582 590218 122026 590454
rect 122262 590218 122346 590454
rect 122582 590218 150026 590454
rect 150262 590218 150346 590454
rect 150582 590218 178026 590454
rect 178262 590218 178346 590454
rect 178582 590218 206026 590454
rect 206262 590218 206346 590454
rect 206582 590218 234026 590454
rect 234262 590218 234346 590454
rect 234582 590218 262026 590454
rect 262262 590218 262346 590454
rect 262582 590218 290026 590454
rect 290262 590218 290346 590454
rect 290582 590218 318026 590454
rect 318262 590218 318346 590454
rect 318582 590218 346026 590454
rect 346262 590218 346346 590454
rect 346582 590218 374026 590454
rect 374262 590218 374346 590454
rect 374582 590218 402026 590454
rect 402262 590218 402346 590454
rect 402582 590218 430026 590454
rect 430262 590218 430346 590454
rect 430582 590218 458026 590454
rect 458262 590218 458346 590454
rect 458582 590218 486026 590454
rect 486262 590218 486346 590454
rect 486582 590218 514026 590454
rect 514262 590218 514346 590454
rect 514582 590218 542026 590454
rect 542262 590218 542346 590454
rect 542582 590218 570026 590454
rect 570262 590218 570346 590454
rect 570582 590218 586302 590454
rect 586538 590218 586622 590454
rect 586858 590218 592650 590454
rect -8726 590134 592650 590218
rect -8726 589898 -2934 590134
rect -2698 589898 -2614 590134
rect -2378 589898 38026 590134
rect 38262 589898 38346 590134
rect 38582 589898 66026 590134
rect 66262 589898 66346 590134
rect 66582 589898 94026 590134
rect 94262 589898 94346 590134
rect 94582 589898 122026 590134
rect 122262 589898 122346 590134
rect 122582 589898 150026 590134
rect 150262 589898 150346 590134
rect 150582 589898 178026 590134
rect 178262 589898 178346 590134
rect 178582 589898 206026 590134
rect 206262 589898 206346 590134
rect 206582 589898 234026 590134
rect 234262 589898 234346 590134
rect 234582 589898 262026 590134
rect 262262 589898 262346 590134
rect 262582 589898 290026 590134
rect 290262 589898 290346 590134
rect 290582 589898 318026 590134
rect 318262 589898 318346 590134
rect 318582 589898 346026 590134
rect 346262 589898 346346 590134
rect 346582 589898 374026 590134
rect 374262 589898 374346 590134
rect 374582 589898 402026 590134
rect 402262 589898 402346 590134
rect 402582 589898 430026 590134
rect 430262 589898 430346 590134
rect 430582 589898 458026 590134
rect 458262 589898 458346 590134
rect 458582 589898 486026 590134
rect 486262 589898 486346 590134
rect 486582 589898 514026 590134
rect 514262 589898 514346 590134
rect 514582 589898 542026 590134
rect 542262 589898 542346 590134
rect 542582 589898 570026 590134
rect 570262 589898 570346 590134
rect 570582 589898 586302 590134
rect 586538 589898 586622 590134
rect 586858 589898 592650 590134
rect -8726 589866 592650 589898
rect -8726 566829 592650 566861
rect -8726 566593 -1974 566829
rect -1738 566593 -1654 566829
rect -1418 566593 41526 566829
rect 41762 566593 41846 566829
rect 42082 566593 69526 566829
rect 69762 566593 69846 566829
rect 70082 566593 97526 566829
rect 97762 566593 97846 566829
rect 98082 566593 125526 566829
rect 125762 566593 125846 566829
rect 126082 566593 153526 566829
rect 153762 566593 153846 566829
rect 154082 566593 181526 566829
rect 181762 566593 181846 566829
rect 182082 566593 209526 566829
rect 209762 566593 209846 566829
rect 210082 566593 237526 566829
rect 237762 566593 237846 566829
rect 238082 566593 265526 566829
rect 265762 566593 265846 566829
rect 266082 566593 293526 566829
rect 293762 566593 293846 566829
rect 294082 566593 321526 566829
rect 321762 566593 321846 566829
rect 322082 566593 349526 566829
rect 349762 566593 349846 566829
rect 350082 566593 377526 566829
rect 377762 566593 377846 566829
rect 378082 566593 405526 566829
rect 405762 566593 405846 566829
rect 406082 566593 433526 566829
rect 433762 566593 433846 566829
rect 434082 566593 461526 566829
rect 461762 566593 461846 566829
rect 462082 566593 489526 566829
rect 489762 566593 489846 566829
rect 490082 566593 517526 566829
rect 517762 566593 517846 566829
rect 518082 566593 545526 566829
rect 545762 566593 545846 566829
rect 546082 566593 573526 566829
rect 573762 566593 573846 566829
rect 574082 566593 585342 566829
rect 585578 566593 585662 566829
rect 585898 566593 592650 566829
rect -8726 566509 592650 566593
rect -8726 566273 -1974 566509
rect -1738 566273 -1654 566509
rect -1418 566273 41526 566509
rect 41762 566273 41846 566509
rect 42082 566273 69526 566509
rect 69762 566273 69846 566509
rect 70082 566273 97526 566509
rect 97762 566273 97846 566509
rect 98082 566273 125526 566509
rect 125762 566273 125846 566509
rect 126082 566273 153526 566509
rect 153762 566273 153846 566509
rect 154082 566273 181526 566509
rect 181762 566273 181846 566509
rect 182082 566273 209526 566509
rect 209762 566273 209846 566509
rect 210082 566273 237526 566509
rect 237762 566273 237846 566509
rect 238082 566273 265526 566509
rect 265762 566273 265846 566509
rect 266082 566273 293526 566509
rect 293762 566273 293846 566509
rect 294082 566273 321526 566509
rect 321762 566273 321846 566509
rect 322082 566273 349526 566509
rect 349762 566273 349846 566509
rect 350082 566273 377526 566509
rect 377762 566273 377846 566509
rect 378082 566273 405526 566509
rect 405762 566273 405846 566509
rect 406082 566273 433526 566509
rect 433762 566273 433846 566509
rect 434082 566273 461526 566509
rect 461762 566273 461846 566509
rect 462082 566273 489526 566509
rect 489762 566273 489846 566509
rect 490082 566273 517526 566509
rect 517762 566273 517846 566509
rect 518082 566273 545526 566509
rect 545762 566273 545846 566509
rect 546082 566273 573526 566509
rect 573762 566273 573846 566509
rect 574082 566273 585342 566509
rect 585578 566273 585662 566509
rect 585898 566273 592650 566509
rect -8726 566241 592650 566273
rect -8726 563454 592650 563486
rect -8726 563218 -2934 563454
rect -2698 563218 -2614 563454
rect -2378 563218 38026 563454
rect 38262 563218 38346 563454
rect 38582 563218 66026 563454
rect 66262 563218 66346 563454
rect 66582 563218 94026 563454
rect 94262 563218 94346 563454
rect 94582 563218 122026 563454
rect 122262 563218 122346 563454
rect 122582 563218 150026 563454
rect 150262 563218 150346 563454
rect 150582 563218 178026 563454
rect 178262 563218 178346 563454
rect 178582 563218 206026 563454
rect 206262 563218 206346 563454
rect 206582 563218 234026 563454
rect 234262 563218 234346 563454
rect 234582 563218 262026 563454
rect 262262 563218 262346 563454
rect 262582 563218 290026 563454
rect 290262 563218 290346 563454
rect 290582 563218 318026 563454
rect 318262 563218 318346 563454
rect 318582 563218 346026 563454
rect 346262 563218 346346 563454
rect 346582 563218 374026 563454
rect 374262 563218 374346 563454
rect 374582 563218 402026 563454
rect 402262 563218 402346 563454
rect 402582 563218 430026 563454
rect 430262 563218 430346 563454
rect 430582 563218 458026 563454
rect 458262 563218 458346 563454
rect 458582 563218 486026 563454
rect 486262 563218 486346 563454
rect 486582 563218 514026 563454
rect 514262 563218 514346 563454
rect 514582 563218 542026 563454
rect 542262 563218 542346 563454
rect 542582 563218 570026 563454
rect 570262 563218 570346 563454
rect 570582 563218 586302 563454
rect 586538 563218 586622 563454
rect 586858 563218 592650 563454
rect -8726 563134 592650 563218
rect -8726 562898 -2934 563134
rect -2698 562898 -2614 563134
rect -2378 562898 38026 563134
rect 38262 562898 38346 563134
rect 38582 562898 66026 563134
rect 66262 562898 66346 563134
rect 66582 562898 94026 563134
rect 94262 562898 94346 563134
rect 94582 562898 122026 563134
rect 122262 562898 122346 563134
rect 122582 562898 150026 563134
rect 150262 562898 150346 563134
rect 150582 562898 178026 563134
rect 178262 562898 178346 563134
rect 178582 562898 206026 563134
rect 206262 562898 206346 563134
rect 206582 562898 234026 563134
rect 234262 562898 234346 563134
rect 234582 562898 262026 563134
rect 262262 562898 262346 563134
rect 262582 562898 290026 563134
rect 290262 562898 290346 563134
rect 290582 562898 318026 563134
rect 318262 562898 318346 563134
rect 318582 562898 346026 563134
rect 346262 562898 346346 563134
rect 346582 562898 374026 563134
rect 374262 562898 374346 563134
rect 374582 562898 402026 563134
rect 402262 562898 402346 563134
rect 402582 562898 430026 563134
rect 430262 562898 430346 563134
rect 430582 562898 458026 563134
rect 458262 562898 458346 563134
rect 458582 562898 486026 563134
rect 486262 562898 486346 563134
rect 486582 562898 514026 563134
rect 514262 562898 514346 563134
rect 514582 562898 542026 563134
rect 542262 562898 542346 563134
rect 542582 562898 570026 563134
rect 570262 562898 570346 563134
rect 570582 562898 586302 563134
rect 586538 562898 586622 563134
rect 586858 562898 592650 563134
rect -8726 562866 592650 562898
rect -8726 539829 592650 539861
rect -8726 539593 -1974 539829
rect -1738 539593 -1654 539829
rect -1418 539593 41526 539829
rect 41762 539593 41846 539829
rect 42082 539593 69526 539829
rect 69762 539593 69846 539829
rect 70082 539593 97526 539829
rect 97762 539593 97846 539829
rect 98082 539593 125526 539829
rect 125762 539593 125846 539829
rect 126082 539593 153526 539829
rect 153762 539593 153846 539829
rect 154082 539593 181526 539829
rect 181762 539593 181846 539829
rect 182082 539593 209526 539829
rect 209762 539593 209846 539829
rect 210082 539593 237526 539829
rect 237762 539593 237846 539829
rect 238082 539593 265526 539829
rect 265762 539593 265846 539829
rect 266082 539593 293526 539829
rect 293762 539593 293846 539829
rect 294082 539593 321526 539829
rect 321762 539593 321846 539829
rect 322082 539593 349526 539829
rect 349762 539593 349846 539829
rect 350082 539593 377526 539829
rect 377762 539593 377846 539829
rect 378082 539593 405526 539829
rect 405762 539593 405846 539829
rect 406082 539593 433526 539829
rect 433762 539593 433846 539829
rect 434082 539593 461526 539829
rect 461762 539593 461846 539829
rect 462082 539593 489526 539829
rect 489762 539593 489846 539829
rect 490082 539593 517526 539829
rect 517762 539593 517846 539829
rect 518082 539593 545526 539829
rect 545762 539593 545846 539829
rect 546082 539593 573526 539829
rect 573762 539593 573846 539829
rect 574082 539593 585342 539829
rect 585578 539593 585662 539829
rect 585898 539593 592650 539829
rect -8726 539509 592650 539593
rect -8726 539273 -1974 539509
rect -1738 539273 -1654 539509
rect -1418 539273 41526 539509
rect 41762 539273 41846 539509
rect 42082 539273 69526 539509
rect 69762 539273 69846 539509
rect 70082 539273 97526 539509
rect 97762 539273 97846 539509
rect 98082 539273 125526 539509
rect 125762 539273 125846 539509
rect 126082 539273 153526 539509
rect 153762 539273 153846 539509
rect 154082 539273 181526 539509
rect 181762 539273 181846 539509
rect 182082 539273 209526 539509
rect 209762 539273 209846 539509
rect 210082 539273 237526 539509
rect 237762 539273 237846 539509
rect 238082 539273 265526 539509
rect 265762 539273 265846 539509
rect 266082 539273 293526 539509
rect 293762 539273 293846 539509
rect 294082 539273 321526 539509
rect 321762 539273 321846 539509
rect 322082 539273 349526 539509
rect 349762 539273 349846 539509
rect 350082 539273 377526 539509
rect 377762 539273 377846 539509
rect 378082 539273 405526 539509
rect 405762 539273 405846 539509
rect 406082 539273 433526 539509
rect 433762 539273 433846 539509
rect 434082 539273 461526 539509
rect 461762 539273 461846 539509
rect 462082 539273 489526 539509
rect 489762 539273 489846 539509
rect 490082 539273 517526 539509
rect 517762 539273 517846 539509
rect 518082 539273 545526 539509
rect 545762 539273 545846 539509
rect 546082 539273 573526 539509
rect 573762 539273 573846 539509
rect 574082 539273 585342 539509
rect 585578 539273 585662 539509
rect 585898 539273 592650 539509
rect -8726 539241 592650 539273
rect -8726 536454 592650 536486
rect -8726 536218 -2934 536454
rect -2698 536218 -2614 536454
rect -2378 536218 38026 536454
rect 38262 536218 38346 536454
rect 38582 536218 66026 536454
rect 66262 536218 66346 536454
rect 66582 536218 94026 536454
rect 94262 536218 94346 536454
rect 94582 536218 122026 536454
rect 122262 536218 122346 536454
rect 122582 536218 150026 536454
rect 150262 536218 150346 536454
rect 150582 536218 178026 536454
rect 178262 536218 178346 536454
rect 178582 536218 206026 536454
rect 206262 536218 206346 536454
rect 206582 536218 234026 536454
rect 234262 536218 234346 536454
rect 234582 536218 262026 536454
rect 262262 536218 262346 536454
rect 262582 536218 290026 536454
rect 290262 536218 290346 536454
rect 290582 536218 318026 536454
rect 318262 536218 318346 536454
rect 318582 536218 346026 536454
rect 346262 536218 346346 536454
rect 346582 536218 374026 536454
rect 374262 536218 374346 536454
rect 374582 536218 402026 536454
rect 402262 536218 402346 536454
rect 402582 536218 430026 536454
rect 430262 536218 430346 536454
rect 430582 536218 458026 536454
rect 458262 536218 458346 536454
rect 458582 536218 486026 536454
rect 486262 536218 486346 536454
rect 486582 536218 514026 536454
rect 514262 536218 514346 536454
rect 514582 536218 542026 536454
rect 542262 536218 542346 536454
rect 542582 536218 570026 536454
rect 570262 536218 570346 536454
rect 570582 536218 586302 536454
rect 586538 536218 586622 536454
rect 586858 536218 592650 536454
rect -8726 536134 592650 536218
rect -8726 535898 -2934 536134
rect -2698 535898 -2614 536134
rect -2378 535898 38026 536134
rect 38262 535898 38346 536134
rect 38582 535898 66026 536134
rect 66262 535898 66346 536134
rect 66582 535898 94026 536134
rect 94262 535898 94346 536134
rect 94582 535898 122026 536134
rect 122262 535898 122346 536134
rect 122582 535898 150026 536134
rect 150262 535898 150346 536134
rect 150582 535898 178026 536134
rect 178262 535898 178346 536134
rect 178582 535898 206026 536134
rect 206262 535898 206346 536134
rect 206582 535898 234026 536134
rect 234262 535898 234346 536134
rect 234582 535898 262026 536134
rect 262262 535898 262346 536134
rect 262582 535898 290026 536134
rect 290262 535898 290346 536134
rect 290582 535898 318026 536134
rect 318262 535898 318346 536134
rect 318582 535898 346026 536134
rect 346262 535898 346346 536134
rect 346582 535898 374026 536134
rect 374262 535898 374346 536134
rect 374582 535898 402026 536134
rect 402262 535898 402346 536134
rect 402582 535898 430026 536134
rect 430262 535898 430346 536134
rect 430582 535898 458026 536134
rect 458262 535898 458346 536134
rect 458582 535898 486026 536134
rect 486262 535898 486346 536134
rect 486582 535898 514026 536134
rect 514262 535898 514346 536134
rect 514582 535898 542026 536134
rect 542262 535898 542346 536134
rect 542582 535898 570026 536134
rect 570262 535898 570346 536134
rect 570582 535898 586302 536134
rect 586538 535898 586622 536134
rect 586858 535898 592650 536134
rect -8726 535866 592650 535898
rect -8726 512829 592650 512861
rect -8726 512593 -1974 512829
rect -1738 512593 -1654 512829
rect -1418 512593 41526 512829
rect 41762 512593 41846 512829
rect 42082 512593 69526 512829
rect 69762 512593 69846 512829
rect 70082 512593 97526 512829
rect 97762 512593 97846 512829
rect 98082 512593 125526 512829
rect 125762 512593 125846 512829
rect 126082 512593 153526 512829
rect 153762 512593 153846 512829
rect 154082 512593 181526 512829
rect 181762 512593 181846 512829
rect 182082 512593 209526 512829
rect 209762 512593 209846 512829
rect 210082 512593 237526 512829
rect 237762 512593 237846 512829
rect 238082 512593 265526 512829
rect 265762 512593 265846 512829
rect 266082 512593 293526 512829
rect 293762 512593 293846 512829
rect 294082 512593 321526 512829
rect 321762 512593 321846 512829
rect 322082 512593 349526 512829
rect 349762 512593 349846 512829
rect 350082 512593 377526 512829
rect 377762 512593 377846 512829
rect 378082 512593 405526 512829
rect 405762 512593 405846 512829
rect 406082 512593 433526 512829
rect 433762 512593 433846 512829
rect 434082 512593 461526 512829
rect 461762 512593 461846 512829
rect 462082 512593 489526 512829
rect 489762 512593 489846 512829
rect 490082 512593 517526 512829
rect 517762 512593 517846 512829
rect 518082 512593 545526 512829
rect 545762 512593 545846 512829
rect 546082 512593 573526 512829
rect 573762 512593 573846 512829
rect 574082 512593 585342 512829
rect 585578 512593 585662 512829
rect 585898 512593 592650 512829
rect -8726 512509 592650 512593
rect -8726 512273 -1974 512509
rect -1738 512273 -1654 512509
rect -1418 512273 41526 512509
rect 41762 512273 41846 512509
rect 42082 512273 69526 512509
rect 69762 512273 69846 512509
rect 70082 512273 97526 512509
rect 97762 512273 97846 512509
rect 98082 512273 125526 512509
rect 125762 512273 125846 512509
rect 126082 512273 153526 512509
rect 153762 512273 153846 512509
rect 154082 512273 181526 512509
rect 181762 512273 181846 512509
rect 182082 512273 209526 512509
rect 209762 512273 209846 512509
rect 210082 512273 237526 512509
rect 237762 512273 237846 512509
rect 238082 512273 265526 512509
rect 265762 512273 265846 512509
rect 266082 512273 293526 512509
rect 293762 512273 293846 512509
rect 294082 512273 321526 512509
rect 321762 512273 321846 512509
rect 322082 512273 349526 512509
rect 349762 512273 349846 512509
rect 350082 512273 377526 512509
rect 377762 512273 377846 512509
rect 378082 512273 405526 512509
rect 405762 512273 405846 512509
rect 406082 512273 433526 512509
rect 433762 512273 433846 512509
rect 434082 512273 461526 512509
rect 461762 512273 461846 512509
rect 462082 512273 489526 512509
rect 489762 512273 489846 512509
rect 490082 512273 517526 512509
rect 517762 512273 517846 512509
rect 518082 512273 545526 512509
rect 545762 512273 545846 512509
rect 546082 512273 573526 512509
rect 573762 512273 573846 512509
rect 574082 512273 585342 512509
rect 585578 512273 585662 512509
rect 585898 512273 592650 512509
rect -8726 512241 592650 512273
rect -8726 509454 592650 509486
rect -8726 509218 -2934 509454
rect -2698 509218 -2614 509454
rect -2378 509218 38026 509454
rect 38262 509218 38346 509454
rect 38582 509218 66026 509454
rect 66262 509218 66346 509454
rect 66582 509218 94026 509454
rect 94262 509218 94346 509454
rect 94582 509218 122026 509454
rect 122262 509218 122346 509454
rect 122582 509218 150026 509454
rect 150262 509218 150346 509454
rect 150582 509218 178026 509454
rect 178262 509218 178346 509454
rect 178582 509218 206026 509454
rect 206262 509218 206346 509454
rect 206582 509218 234026 509454
rect 234262 509218 234346 509454
rect 234582 509218 262026 509454
rect 262262 509218 262346 509454
rect 262582 509218 290026 509454
rect 290262 509218 290346 509454
rect 290582 509218 318026 509454
rect 318262 509218 318346 509454
rect 318582 509218 346026 509454
rect 346262 509218 346346 509454
rect 346582 509218 374026 509454
rect 374262 509218 374346 509454
rect 374582 509218 402026 509454
rect 402262 509218 402346 509454
rect 402582 509218 430026 509454
rect 430262 509218 430346 509454
rect 430582 509218 458026 509454
rect 458262 509218 458346 509454
rect 458582 509218 486026 509454
rect 486262 509218 486346 509454
rect 486582 509218 514026 509454
rect 514262 509218 514346 509454
rect 514582 509218 542026 509454
rect 542262 509218 542346 509454
rect 542582 509218 570026 509454
rect 570262 509218 570346 509454
rect 570582 509218 586302 509454
rect 586538 509218 586622 509454
rect 586858 509218 592650 509454
rect -8726 509134 592650 509218
rect -8726 508898 -2934 509134
rect -2698 508898 -2614 509134
rect -2378 508898 38026 509134
rect 38262 508898 38346 509134
rect 38582 508898 66026 509134
rect 66262 508898 66346 509134
rect 66582 508898 94026 509134
rect 94262 508898 94346 509134
rect 94582 508898 122026 509134
rect 122262 508898 122346 509134
rect 122582 508898 150026 509134
rect 150262 508898 150346 509134
rect 150582 508898 178026 509134
rect 178262 508898 178346 509134
rect 178582 508898 206026 509134
rect 206262 508898 206346 509134
rect 206582 508898 234026 509134
rect 234262 508898 234346 509134
rect 234582 508898 262026 509134
rect 262262 508898 262346 509134
rect 262582 508898 290026 509134
rect 290262 508898 290346 509134
rect 290582 508898 318026 509134
rect 318262 508898 318346 509134
rect 318582 508898 346026 509134
rect 346262 508898 346346 509134
rect 346582 508898 374026 509134
rect 374262 508898 374346 509134
rect 374582 508898 402026 509134
rect 402262 508898 402346 509134
rect 402582 508898 430026 509134
rect 430262 508898 430346 509134
rect 430582 508898 458026 509134
rect 458262 508898 458346 509134
rect 458582 508898 486026 509134
rect 486262 508898 486346 509134
rect 486582 508898 514026 509134
rect 514262 508898 514346 509134
rect 514582 508898 542026 509134
rect 542262 508898 542346 509134
rect 542582 508898 570026 509134
rect 570262 508898 570346 509134
rect 570582 508898 586302 509134
rect 586538 508898 586622 509134
rect 586858 508898 592650 509134
rect -8726 508866 592650 508898
rect -8726 485829 592650 485861
rect -8726 485593 -1974 485829
rect -1738 485593 -1654 485829
rect -1418 485593 41526 485829
rect 41762 485593 41846 485829
rect 42082 485593 69526 485829
rect 69762 485593 69846 485829
rect 70082 485593 97526 485829
rect 97762 485593 97846 485829
rect 98082 485593 125526 485829
rect 125762 485593 125846 485829
rect 126082 485593 153526 485829
rect 153762 485593 153846 485829
rect 154082 485593 181526 485829
rect 181762 485593 181846 485829
rect 182082 485593 209526 485829
rect 209762 485593 209846 485829
rect 210082 485593 237526 485829
rect 237762 485593 237846 485829
rect 238082 485593 265526 485829
rect 265762 485593 265846 485829
rect 266082 485593 293526 485829
rect 293762 485593 293846 485829
rect 294082 485593 321526 485829
rect 321762 485593 321846 485829
rect 322082 485593 349526 485829
rect 349762 485593 349846 485829
rect 350082 485593 377526 485829
rect 377762 485593 377846 485829
rect 378082 485593 405526 485829
rect 405762 485593 405846 485829
rect 406082 485593 433526 485829
rect 433762 485593 433846 485829
rect 434082 485593 461526 485829
rect 461762 485593 461846 485829
rect 462082 485593 489526 485829
rect 489762 485593 489846 485829
rect 490082 485593 517526 485829
rect 517762 485593 517846 485829
rect 518082 485593 545526 485829
rect 545762 485593 545846 485829
rect 546082 485593 573526 485829
rect 573762 485593 573846 485829
rect 574082 485593 585342 485829
rect 585578 485593 585662 485829
rect 585898 485593 592650 485829
rect -8726 485509 592650 485593
rect -8726 485273 -1974 485509
rect -1738 485273 -1654 485509
rect -1418 485273 41526 485509
rect 41762 485273 41846 485509
rect 42082 485273 69526 485509
rect 69762 485273 69846 485509
rect 70082 485273 97526 485509
rect 97762 485273 97846 485509
rect 98082 485273 125526 485509
rect 125762 485273 125846 485509
rect 126082 485273 153526 485509
rect 153762 485273 153846 485509
rect 154082 485273 181526 485509
rect 181762 485273 181846 485509
rect 182082 485273 209526 485509
rect 209762 485273 209846 485509
rect 210082 485273 237526 485509
rect 237762 485273 237846 485509
rect 238082 485273 265526 485509
rect 265762 485273 265846 485509
rect 266082 485273 293526 485509
rect 293762 485273 293846 485509
rect 294082 485273 321526 485509
rect 321762 485273 321846 485509
rect 322082 485273 349526 485509
rect 349762 485273 349846 485509
rect 350082 485273 377526 485509
rect 377762 485273 377846 485509
rect 378082 485273 405526 485509
rect 405762 485273 405846 485509
rect 406082 485273 433526 485509
rect 433762 485273 433846 485509
rect 434082 485273 461526 485509
rect 461762 485273 461846 485509
rect 462082 485273 489526 485509
rect 489762 485273 489846 485509
rect 490082 485273 517526 485509
rect 517762 485273 517846 485509
rect 518082 485273 545526 485509
rect 545762 485273 545846 485509
rect 546082 485273 573526 485509
rect 573762 485273 573846 485509
rect 574082 485273 585342 485509
rect 585578 485273 585662 485509
rect 585898 485273 592650 485509
rect -8726 485241 592650 485273
rect -8726 482454 592650 482486
rect -8726 482218 -2934 482454
rect -2698 482218 -2614 482454
rect -2378 482218 38026 482454
rect 38262 482218 38346 482454
rect 38582 482218 66026 482454
rect 66262 482218 66346 482454
rect 66582 482218 94026 482454
rect 94262 482218 94346 482454
rect 94582 482218 122026 482454
rect 122262 482218 122346 482454
rect 122582 482218 150026 482454
rect 150262 482218 150346 482454
rect 150582 482218 178026 482454
rect 178262 482218 178346 482454
rect 178582 482218 206026 482454
rect 206262 482218 206346 482454
rect 206582 482218 234026 482454
rect 234262 482218 234346 482454
rect 234582 482218 262026 482454
rect 262262 482218 262346 482454
rect 262582 482218 290026 482454
rect 290262 482218 290346 482454
rect 290582 482218 318026 482454
rect 318262 482218 318346 482454
rect 318582 482218 346026 482454
rect 346262 482218 346346 482454
rect 346582 482218 374026 482454
rect 374262 482218 374346 482454
rect 374582 482218 402026 482454
rect 402262 482218 402346 482454
rect 402582 482218 430026 482454
rect 430262 482218 430346 482454
rect 430582 482218 458026 482454
rect 458262 482218 458346 482454
rect 458582 482218 486026 482454
rect 486262 482218 486346 482454
rect 486582 482218 514026 482454
rect 514262 482218 514346 482454
rect 514582 482218 542026 482454
rect 542262 482218 542346 482454
rect 542582 482218 570026 482454
rect 570262 482218 570346 482454
rect 570582 482218 586302 482454
rect 586538 482218 586622 482454
rect 586858 482218 592650 482454
rect -8726 482134 592650 482218
rect -8726 481898 -2934 482134
rect -2698 481898 -2614 482134
rect -2378 481898 38026 482134
rect 38262 481898 38346 482134
rect 38582 481898 66026 482134
rect 66262 481898 66346 482134
rect 66582 481898 94026 482134
rect 94262 481898 94346 482134
rect 94582 481898 122026 482134
rect 122262 481898 122346 482134
rect 122582 481898 150026 482134
rect 150262 481898 150346 482134
rect 150582 481898 178026 482134
rect 178262 481898 178346 482134
rect 178582 481898 206026 482134
rect 206262 481898 206346 482134
rect 206582 481898 234026 482134
rect 234262 481898 234346 482134
rect 234582 481898 262026 482134
rect 262262 481898 262346 482134
rect 262582 481898 290026 482134
rect 290262 481898 290346 482134
rect 290582 481898 318026 482134
rect 318262 481898 318346 482134
rect 318582 481898 346026 482134
rect 346262 481898 346346 482134
rect 346582 481898 374026 482134
rect 374262 481898 374346 482134
rect 374582 481898 402026 482134
rect 402262 481898 402346 482134
rect 402582 481898 430026 482134
rect 430262 481898 430346 482134
rect 430582 481898 458026 482134
rect 458262 481898 458346 482134
rect 458582 481898 486026 482134
rect 486262 481898 486346 482134
rect 486582 481898 514026 482134
rect 514262 481898 514346 482134
rect 514582 481898 542026 482134
rect 542262 481898 542346 482134
rect 542582 481898 570026 482134
rect 570262 481898 570346 482134
rect 570582 481898 586302 482134
rect 586538 481898 586622 482134
rect 586858 481898 592650 482134
rect -8726 481866 592650 481898
rect -8726 458829 592650 458861
rect -8726 458593 -1974 458829
rect -1738 458593 -1654 458829
rect -1418 458593 41526 458829
rect 41762 458593 41846 458829
rect 42082 458593 69526 458829
rect 69762 458593 69846 458829
rect 70082 458593 97526 458829
rect 97762 458593 97846 458829
rect 98082 458593 125526 458829
rect 125762 458593 125846 458829
rect 126082 458593 153526 458829
rect 153762 458593 153846 458829
rect 154082 458593 181526 458829
rect 181762 458593 181846 458829
rect 182082 458593 209526 458829
rect 209762 458593 209846 458829
rect 210082 458593 237526 458829
rect 237762 458593 237846 458829
rect 238082 458593 265526 458829
rect 265762 458593 265846 458829
rect 266082 458593 293526 458829
rect 293762 458593 293846 458829
rect 294082 458593 321526 458829
rect 321762 458593 321846 458829
rect 322082 458593 349526 458829
rect 349762 458593 349846 458829
rect 350082 458593 377526 458829
rect 377762 458593 377846 458829
rect 378082 458593 405526 458829
rect 405762 458593 405846 458829
rect 406082 458593 433526 458829
rect 433762 458593 433846 458829
rect 434082 458593 461526 458829
rect 461762 458593 461846 458829
rect 462082 458593 489526 458829
rect 489762 458593 489846 458829
rect 490082 458593 517526 458829
rect 517762 458593 517846 458829
rect 518082 458593 545526 458829
rect 545762 458593 545846 458829
rect 546082 458593 573526 458829
rect 573762 458593 573846 458829
rect 574082 458593 585342 458829
rect 585578 458593 585662 458829
rect 585898 458593 592650 458829
rect -8726 458509 592650 458593
rect -8726 458273 -1974 458509
rect -1738 458273 -1654 458509
rect -1418 458273 41526 458509
rect 41762 458273 41846 458509
rect 42082 458273 69526 458509
rect 69762 458273 69846 458509
rect 70082 458273 97526 458509
rect 97762 458273 97846 458509
rect 98082 458273 125526 458509
rect 125762 458273 125846 458509
rect 126082 458273 153526 458509
rect 153762 458273 153846 458509
rect 154082 458273 181526 458509
rect 181762 458273 181846 458509
rect 182082 458273 209526 458509
rect 209762 458273 209846 458509
rect 210082 458273 237526 458509
rect 237762 458273 237846 458509
rect 238082 458273 265526 458509
rect 265762 458273 265846 458509
rect 266082 458273 293526 458509
rect 293762 458273 293846 458509
rect 294082 458273 321526 458509
rect 321762 458273 321846 458509
rect 322082 458273 349526 458509
rect 349762 458273 349846 458509
rect 350082 458273 377526 458509
rect 377762 458273 377846 458509
rect 378082 458273 405526 458509
rect 405762 458273 405846 458509
rect 406082 458273 433526 458509
rect 433762 458273 433846 458509
rect 434082 458273 461526 458509
rect 461762 458273 461846 458509
rect 462082 458273 489526 458509
rect 489762 458273 489846 458509
rect 490082 458273 517526 458509
rect 517762 458273 517846 458509
rect 518082 458273 545526 458509
rect 545762 458273 545846 458509
rect 546082 458273 573526 458509
rect 573762 458273 573846 458509
rect 574082 458273 585342 458509
rect 585578 458273 585662 458509
rect 585898 458273 592650 458509
rect -8726 458241 592650 458273
rect -8726 455454 592650 455486
rect -8726 455218 -2934 455454
rect -2698 455218 -2614 455454
rect -2378 455218 38026 455454
rect 38262 455218 38346 455454
rect 38582 455218 66026 455454
rect 66262 455218 66346 455454
rect 66582 455218 94026 455454
rect 94262 455218 94346 455454
rect 94582 455218 122026 455454
rect 122262 455218 122346 455454
rect 122582 455218 150026 455454
rect 150262 455218 150346 455454
rect 150582 455218 178026 455454
rect 178262 455218 178346 455454
rect 178582 455218 206026 455454
rect 206262 455218 206346 455454
rect 206582 455218 234026 455454
rect 234262 455218 234346 455454
rect 234582 455218 262026 455454
rect 262262 455218 262346 455454
rect 262582 455218 290026 455454
rect 290262 455218 290346 455454
rect 290582 455218 318026 455454
rect 318262 455218 318346 455454
rect 318582 455218 346026 455454
rect 346262 455218 346346 455454
rect 346582 455218 374026 455454
rect 374262 455218 374346 455454
rect 374582 455218 402026 455454
rect 402262 455218 402346 455454
rect 402582 455218 430026 455454
rect 430262 455218 430346 455454
rect 430582 455218 458026 455454
rect 458262 455218 458346 455454
rect 458582 455218 486026 455454
rect 486262 455218 486346 455454
rect 486582 455218 514026 455454
rect 514262 455218 514346 455454
rect 514582 455218 542026 455454
rect 542262 455218 542346 455454
rect 542582 455218 570026 455454
rect 570262 455218 570346 455454
rect 570582 455218 586302 455454
rect 586538 455218 586622 455454
rect 586858 455218 592650 455454
rect -8726 455134 592650 455218
rect -8726 454898 -2934 455134
rect -2698 454898 -2614 455134
rect -2378 454898 38026 455134
rect 38262 454898 38346 455134
rect 38582 454898 66026 455134
rect 66262 454898 66346 455134
rect 66582 454898 94026 455134
rect 94262 454898 94346 455134
rect 94582 454898 122026 455134
rect 122262 454898 122346 455134
rect 122582 454898 150026 455134
rect 150262 454898 150346 455134
rect 150582 454898 178026 455134
rect 178262 454898 178346 455134
rect 178582 454898 206026 455134
rect 206262 454898 206346 455134
rect 206582 454898 234026 455134
rect 234262 454898 234346 455134
rect 234582 454898 262026 455134
rect 262262 454898 262346 455134
rect 262582 454898 290026 455134
rect 290262 454898 290346 455134
rect 290582 454898 318026 455134
rect 318262 454898 318346 455134
rect 318582 454898 346026 455134
rect 346262 454898 346346 455134
rect 346582 454898 374026 455134
rect 374262 454898 374346 455134
rect 374582 454898 402026 455134
rect 402262 454898 402346 455134
rect 402582 454898 430026 455134
rect 430262 454898 430346 455134
rect 430582 454898 458026 455134
rect 458262 454898 458346 455134
rect 458582 454898 486026 455134
rect 486262 454898 486346 455134
rect 486582 454898 514026 455134
rect 514262 454898 514346 455134
rect 514582 454898 542026 455134
rect 542262 454898 542346 455134
rect 542582 454898 570026 455134
rect 570262 454898 570346 455134
rect 570582 454898 586302 455134
rect 586538 454898 586622 455134
rect 586858 454898 592650 455134
rect -8726 454866 592650 454898
rect -8726 431829 592650 431861
rect -8726 431593 -1974 431829
rect -1738 431593 -1654 431829
rect -1418 431593 41526 431829
rect 41762 431593 41846 431829
rect 42082 431593 69526 431829
rect 69762 431593 69846 431829
rect 70082 431593 97526 431829
rect 97762 431593 97846 431829
rect 98082 431593 125526 431829
rect 125762 431593 125846 431829
rect 126082 431593 153526 431829
rect 153762 431593 153846 431829
rect 154082 431593 181526 431829
rect 181762 431593 181846 431829
rect 182082 431593 209526 431829
rect 209762 431593 209846 431829
rect 210082 431593 237526 431829
rect 237762 431593 237846 431829
rect 238082 431593 265526 431829
rect 265762 431593 265846 431829
rect 266082 431593 293526 431829
rect 293762 431593 293846 431829
rect 294082 431593 321526 431829
rect 321762 431593 321846 431829
rect 322082 431593 349526 431829
rect 349762 431593 349846 431829
rect 350082 431593 377526 431829
rect 377762 431593 377846 431829
rect 378082 431593 405526 431829
rect 405762 431593 405846 431829
rect 406082 431593 433526 431829
rect 433762 431593 433846 431829
rect 434082 431593 461526 431829
rect 461762 431593 461846 431829
rect 462082 431593 489526 431829
rect 489762 431593 489846 431829
rect 490082 431593 517526 431829
rect 517762 431593 517846 431829
rect 518082 431593 545526 431829
rect 545762 431593 545846 431829
rect 546082 431593 573526 431829
rect 573762 431593 573846 431829
rect 574082 431593 585342 431829
rect 585578 431593 585662 431829
rect 585898 431593 592650 431829
rect -8726 431509 592650 431593
rect -8726 431273 -1974 431509
rect -1738 431273 -1654 431509
rect -1418 431273 41526 431509
rect 41762 431273 41846 431509
rect 42082 431273 69526 431509
rect 69762 431273 69846 431509
rect 70082 431273 97526 431509
rect 97762 431273 97846 431509
rect 98082 431273 125526 431509
rect 125762 431273 125846 431509
rect 126082 431273 153526 431509
rect 153762 431273 153846 431509
rect 154082 431273 181526 431509
rect 181762 431273 181846 431509
rect 182082 431273 209526 431509
rect 209762 431273 209846 431509
rect 210082 431273 237526 431509
rect 237762 431273 237846 431509
rect 238082 431273 265526 431509
rect 265762 431273 265846 431509
rect 266082 431273 293526 431509
rect 293762 431273 293846 431509
rect 294082 431273 321526 431509
rect 321762 431273 321846 431509
rect 322082 431273 349526 431509
rect 349762 431273 349846 431509
rect 350082 431273 377526 431509
rect 377762 431273 377846 431509
rect 378082 431273 405526 431509
rect 405762 431273 405846 431509
rect 406082 431273 433526 431509
rect 433762 431273 433846 431509
rect 434082 431273 461526 431509
rect 461762 431273 461846 431509
rect 462082 431273 489526 431509
rect 489762 431273 489846 431509
rect 490082 431273 517526 431509
rect 517762 431273 517846 431509
rect 518082 431273 545526 431509
rect 545762 431273 545846 431509
rect 546082 431273 573526 431509
rect 573762 431273 573846 431509
rect 574082 431273 585342 431509
rect 585578 431273 585662 431509
rect 585898 431273 592650 431509
rect -8726 431241 592650 431273
rect -8726 428454 592650 428486
rect -8726 428218 -2934 428454
rect -2698 428218 -2614 428454
rect -2378 428218 38026 428454
rect 38262 428218 38346 428454
rect 38582 428218 66026 428454
rect 66262 428218 66346 428454
rect 66582 428218 94026 428454
rect 94262 428218 94346 428454
rect 94582 428218 122026 428454
rect 122262 428218 122346 428454
rect 122582 428218 150026 428454
rect 150262 428218 150346 428454
rect 150582 428218 178026 428454
rect 178262 428218 178346 428454
rect 178582 428218 206026 428454
rect 206262 428218 206346 428454
rect 206582 428218 234026 428454
rect 234262 428218 234346 428454
rect 234582 428218 262026 428454
rect 262262 428218 262346 428454
rect 262582 428218 290026 428454
rect 290262 428218 290346 428454
rect 290582 428218 318026 428454
rect 318262 428218 318346 428454
rect 318582 428218 346026 428454
rect 346262 428218 346346 428454
rect 346582 428218 374026 428454
rect 374262 428218 374346 428454
rect 374582 428218 402026 428454
rect 402262 428218 402346 428454
rect 402582 428218 430026 428454
rect 430262 428218 430346 428454
rect 430582 428218 458026 428454
rect 458262 428218 458346 428454
rect 458582 428218 486026 428454
rect 486262 428218 486346 428454
rect 486582 428218 514026 428454
rect 514262 428218 514346 428454
rect 514582 428218 542026 428454
rect 542262 428218 542346 428454
rect 542582 428218 570026 428454
rect 570262 428218 570346 428454
rect 570582 428218 586302 428454
rect 586538 428218 586622 428454
rect 586858 428218 592650 428454
rect -8726 428134 592650 428218
rect -8726 427898 -2934 428134
rect -2698 427898 -2614 428134
rect -2378 427898 38026 428134
rect 38262 427898 38346 428134
rect 38582 427898 66026 428134
rect 66262 427898 66346 428134
rect 66582 427898 94026 428134
rect 94262 427898 94346 428134
rect 94582 427898 122026 428134
rect 122262 427898 122346 428134
rect 122582 427898 150026 428134
rect 150262 427898 150346 428134
rect 150582 427898 178026 428134
rect 178262 427898 178346 428134
rect 178582 427898 206026 428134
rect 206262 427898 206346 428134
rect 206582 427898 234026 428134
rect 234262 427898 234346 428134
rect 234582 427898 262026 428134
rect 262262 427898 262346 428134
rect 262582 427898 290026 428134
rect 290262 427898 290346 428134
rect 290582 427898 318026 428134
rect 318262 427898 318346 428134
rect 318582 427898 346026 428134
rect 346262 427898 346346 428134
rect 346582 427898 374026 428134
rect 374262 427898 374346 428134
rect 374582 427898 402026 428134
rect 402262 427898 402346 428134
rect 402582 427898 430026 428134
rect 430262 427898 430346 428134
rect 430582 427898 458026 428134
rect 458262 427898 458346 428134
rect 458582 427898 486026 428134
rect 486262 427898 486346 428134
rect 486582 427898 514026 428134
rect 514262 427898 514346 428134
rect 514582 427898 542026 428134
rect 542262 427898 542346 428134
rect 542582 427898 570026 428134
rect 570262 427898 570346 428134
rect 570582 427898 586302 428134
rect 586538 427898 586622 428134
rect 586858 427898 592650 428134
rect -8726 427866 592650 427898
rect -8726 404829 592650 404861
rect -8726 404593 -1974 404829
rect -1738 404593 -1654 404829
rect -1418 404593 41526 404829
rect 41762 404593 41846 404829
rect 42082 404593 69526 404829
rect 69762 404593 69846 404829
rect 70082 404593 97526 404829
rect 97762 404593 97846 404829
rect 98082 404593 125526 404829
rect 125762 404593 125846 404829
rect 126082 404593 153526 404829
rect 153762 404593 153846 404829
rect 154082 404593 181526 404829
rect 181762 404593 181846 404829
rect 182082 404593 209526 404829
rect 209762 404593 209846 404829
rect 210082 404593 237526 404829
rect 237762 404593 237846 404829
rect 238082 404593 265526 404829
rect 265762 404593 265846 404829
rect 266082 404593 293526 404829
rect 293762 404593 293846 404829
rect 294082 404593 321526 404829
rect 321762 404593 321846 404829
rect 322082 404593 349526 404829
rect 349762 404593 349846 404829
rect 350082 404593 377526 404829
rect 377762 404593 377846 404829
rect 378082 404593 405526 404829
rect 405762 404593 405846 404829
rect 406082 404593 433526 404829
rect 433762 404593 433846 404829
rect 434082 404593 461526 404829
rect 461762 404593 461846 404829
rect 462082 404593 489526 404829
rect 489762 404593 489846 404829
rect 490082 404593 517526 404829
rect 517762 404593 517846 404829
rect 518082 404593 545526 404829
rect 545762 404593 545846 404829
rect 546082 404593 573526 404829
rect 573762 404593 573846 404829
rect 574082 404593 585342 404829
rect 585578 404593 585662 404829
rect 585898 404593 592650 404829
rect -8726 404509 592650 404593
rect -8726 404273 -1974 404509
rect -1738 404273 -1654 404509
rect -1418 404273 41526 404509
rect 41762 404273 41846 404509
rect 42082 404273 69526 404509
rect 69762 404273 69846 404509
rect 70082 404273 97526 404509
rect 97762 404273 97846 404509
rect 98082 404273 125526 404509
rect 125762 404273 125846 404509
rect 126082 404273 153526 404509
rect 153762 404273 153846 404509
rect 154082 404273 181526 404509
rect 181762 404273 181846 404509
rect 182082 404273 209526 404509
rect 209762 404273 209846 404509
rect 210082 404273 237526 404509
rect 237762 404273 237846 404509
rect 238082 404273 265526 404509
rect 265762 404273 265846 404509
rect 266082 404273 293526 404509
rect 293762 404273 293846 404509
rect 294082 404273 321526 404509
rect 321762 404273 321846 404509
rect 322082 404273 349526 404509
rect 349762 404273 349846 404509
rect 350082 404273 377526 404509
rect 377762 404273 377846 404509
rect 378082 404273 405526 404509
rect 405762 404273 405846 404509
rect 406082 404273 433526 404509
rect 433762 404273 433846 404509
rect 434082 404273 461526 404509
rect 461762 404273 461846 404509
rect 462082 404273 489526 404509
rect 489762 404273 489846 404509
rect 490082 404273 517526 404509
rect 517762 404273 517846 404509
rect 518082 404273 545526 404509
rect 545762 404273 545846 404509
rect 546082 404273 573526 404509
rect 573762 404273 573846 404509
rect 574082 404273 585342 404509
rect 585578 404273 585662 404509
rect 585898 404273 592650 404509
rect -8726 404241 592650 404273
rect -8726 401454 592650 401486
rect -8726 401218 -2934 401454
rect -2698 401218 -2614 401454
rect -2378 401218 38026 401454
rect 38262 401218 38346 401454
rect 38582 401218 66026 401454
rect 66262 401218 66346 401454
rect 66582 401218 94026 401454
rect 94262 401218 94346 401454
rect 94582 401218 122026 401454
rect 122262 401218 122346 401454
rect 122582 401218 150026 401454
rect 150262 401218 150346 401454
rect 150582 401218 178026 401454
rect 178262 401218 178346 401454
rect 178582 401218 206026 401454
rect 206262 401218 206346 401454
rect 206582 401218 234026 401454
rect 234262 401218 234346 401454
rect 234582 401218 262026 401454
rect 262262 401218 262346 401454
rect 262582 401218 290026 401454
rect 290262 401218 290346 401454
rect 290582 401218 318026 401454
rect 318262 401218 318346 401454
rect 318582 401218 346026 401454
rect 346262 401218 346346 401454
rect 346582 401218 374026 401454
rect 374262 401218 374346 401454
rect 374582 401218 402026 401454
rect 402262 401218 402346 401454
rect 402582 401218 430026 401454
rect 430262 401218 430346 401454
rect 430582 401218 458026 401454
rect 458262 401218 458346 401454
rect 458582 401218 486026 401454
rect 486262 401218 486346 401454
rect 486582 401218 514026 401454
rect 514262 401218 514346 401454
rect 514582 401218 542026 401454
rect 542262 401218 542346 401454
rect 542582 401218 570026 401454
rect 570262 401218 570346 401454
rect 570582 401218 586302 401454
rect 586538 401218 586622 401454
rect 586858 401218 592650 401454
rect -8726 401134 592650 401218
rect -8726 400898 -2934 401134
rect -2698 400898 -2614 401134
rect -2378 400898 38026 401134
rect 38262 400898 38346 401134
rect 38582 400898 66026 401134
rect 66262 400898 66346 401134
rect 66582 400898 94026 401134
rect 94262 400898 94346 401134
rect 94582 400898 122026 401134
rect 122262 400898 122346 401134
rect 122582 400898 150026 401134
rect 150262 400898 150346 401134
rect 150582 400898 178026 401134
rect 178262 400898 178346 401134
rect 178582 400898 206026 401134
rect 206262 400898 206346 401134
rect 206582 400898 234026 401134
rect 234262 400898 234346 401134
rect 234582 400898 262026 401134
rect 262262 400898 262346 401134
rect 262582 400898 290026 401134
rect 290262 400898 290346 401134
rect 290582 400898 318026 401134
rect 318262 400898 318346 401134
rect 318582 400898 346026 401134
rect 346262 400898 346346 401134
rect 346582 400898 374026 401134
rect 374262 400898 374346 401134
rect 374582 400898 402026 401134
rect 402262 400898 402346 401134
rect 402582 400898 430026 401134
rect 430262 400898 430346 401134
rect 430582 400898 458026 401134
rect 458262 400898 458346 401134
rect 458582 400898 486026 401134
rect 486262 400898 486346 401134
rect 486582 400898 514026 401134
rect 514262 400898 514346 401134
rect 514582 400898 542026 401134
rect 542262 400898 542346 401134
rect 542582 400898 570026 401134
rect 570262 400898 570346 401134
rect 570582 400898 586302 401134
rect 586538 400898 586622 401134
rect 586858 400898 592650 401134
rect -8726 400866 592650 400898
rect -8726 377829 592650 377861
rect -8726 377593 -1974 377829
rect -1738 377593 -1654 377829
rect -1418 377593 41526 377829
rect 41762 377593 41846 377829
rect 42082 377593 69526 377829
rect 69762 377593 69846 377829
rect 70082 377593 97526 377829
rect 97762 377593 97846 377829
rect 98082 377593 125526 377829
rect 125762 377593 125846 377829
rect 126082 377593 153526 377829
rect 153762 377593 153846 377829
rect 154082 377593 181526 377829
rect 181762 377593 181846 377829
rect 182082 377593 209526 377829
rect 209762 377593 209846 377829
rect 210082 377593 237526 377829
rect 237762 377593 237846 377829
rect 238082 377593 265526 377829
rect 265762 377593 265846 377829
rect 266082 377593 293526 377829
rect 293762 377593 293846 377829
rect 294082 377593 321526 377829
rect 321762 377593 321846 377829
rect 322082 377593 349526 377829
rect 349762 377593 349846 377829
rect 350082 377593 377526 377829
rect 377762 377593 377846 377829
rect 378082 377593 405526 377829
rect 405762 377593 405846 377829
rect 406082 377593 433526 377829
rect 433762 377593 433846 377829
rect 434082 377593 461526 377829
rect 461762 377593 461846 377829
rect 462082 377593 489526 377829
rect 489762 377593 489846 377829
rect 490082 377593 517526 377829
rect 517762 377593 517846 377829
rect 518082 377593 545526 377829
rect 545762 377593 545846 377829
rect 546082 377593 573526 377829
rect 573762 377593 573846 377829
rect 574082 377593 585342 377829
rect 585578 377593 585662 377829
rect 585898 377593 592650 377829
rect -8726 377509 592650 377593
rect -8726 377273 -1974 377509
rect -1738 377273 -1654 377509
rect -1418 377273 41526 377509
rect 41762 377273 41846 377509
rect 42082 377273 69526 377509
rect 69762 377273 69846 377509
rect 70082 377273 97526 377509
rect 97762 377273 97846 377509
rect 98082 377273 125526 377509
rect 125762 377273 125846 377509
rect 126082 377273 153526 377509
rect 153762 377273 153846 377509
rect 154082 377273 181526 377509
rect 181762 377273 181846 377509
rect 182082 377273 209526 377509
rect 209762 377273 209846 377509
rect 210082 377273 237526 377509
rect 237762 377273 237846 377509
rect 238082 377273 265526 377509
rect 265762 377273 265846 377509
rect 266082 377273 293526 377509
rect 293762 377273 293846 377509
rect 294082 377273 321526 377509
rect 321762 377273 321846 377509
rect 322082 377273 349526 377509
rect 349762 377273 349846 377509
rect 350082 377273 377526 377509
rect 377762 377273 377846 377509
rect 378082 377273 405526 377509
rect 405762 377273 405846 377509
rect 406082 377273 433526 377509
rect 433762 377273 433846 377509
rect 434082 377273 461526 377509
rect 461762 377273 461846 377509
rect 462082 377273 489526 377509
rect 489762 377273 489846 377509
rect 490082 377273 517526 377509
rect 517762 377273 517846 377509
rect 518082 377273 545526 377509
rect 545762 377273 545846 377509
rect 546082 377273 573526 377509
rect 573762 377273 573846 377509
rect 574082 377273 585342 377509
rect 585578 377273 585662 377509
rect 585898 377273 592650 377509
rect -8726 377241 592650 377273
rect -8726 374454 592650 374486
rect -8726 374218 -2934 374454
rect -2698 374218 -2614 374454
rect -2378 374218 38026 374454
rect 38262 374218 38346 374454
rect 38582 374218 66026 374454
rect 66262 374218 66346 374454
rect 66582 374218 94026 374454
rect 94262 374218 94346 374454
rect 94582 374218 122026 374454
rect 122262 374218 122346 374454
rect 122582 374218 150026 374454
rect 150262 374218 150346 374454
rect 150582 374218 178026 374454
rect 178262 374218 178346 374454
rect 178582 374218 206026 374454
rect 206262 374218 206346 374454
rect 206582 374218 234026 374454
rect 234262 374218 234346 374454
rect 234582 374218 262026 374454
rect 262262 374218 262346 374454
rect 262582 374218 290026 374454
rect 290262 374218 290346 374454
rect 290582 374218 318026 374454
rect 318262 374218 318346 374454
rect 318582 374218 346026 374454
rect 346262 374218 346346 374454
rect 346582 374218 374026 374454
rect 374262 374218 374346 374454
rect 374582 374218 402026 374454
rect 402262 374218 402346 374454
rect 402582 374218 430026 374454
rect 430262 374218 430346 374454
rect 430582 374218 458026 374454
rect 458262 374218 458346 374454
rect 458582 374218 486026 374454
rect 486262 374218 486346 374454
rect 486582 374218 514026 374454
rect 514262 374218 514346 374454
rect 514582 374218 542026 374454
rect 542262 374218 542346 374454
rect 542582 374218 570026 374454
rect 570262 374218 570346 374454
rect 570582 374218 586302 374454
rect 586538 374218 586622 374454
rect 586858 374218 592650 374454
rect -8726 374134 592650 374218
rect -8726 373898 -2934 374134
rect -2698 373898 -2614 374134
rect -2378 373898 38026 374134
rect 38262 373898 38346 374134
rect 38582 373898 66026 374134
rect 66262 373898 66346 374134
rect 66582 373898 94026 374134
rect 94262 373898 94346 374134
rect 94582 373898 122026 374134
rect 122262 373898 122346 374134
rect 122582 373898 150026 374134
rect 150262 373898 150346 374134
rect 150582 373898 178026 374134
rect 178262 373898 178346 374134
rect 178582 373898 206026 374134
rect 206262 373898 206346 374134
rect 206582 373898 234026 374134
rect 234262 373898 234346 374134
rect 234582 373898 262026 374134
rect 262262 373898 262346 374134
rect 262582 373898 290026 374134
rect 290262 373898 290346 374134
rect 290582 373898 318026 374134
rect 318262 373898 318346 374134
rect 318582 373898 346026 374134
rect 346262 373898 346346 374134
rect 346582 373898 374026 374134
rect 374262 373898 374346 374134
rect 374582 373898 402026 374134
rect 402262 373898 402346 374134
rect 402582 373898 430026 374134
rect 430262 373898 430346 374134
rect 430582 373898 458026 374134
rect 458262 373898 458346 374134
rect 458582 373898 486026 374134
rect 486262 373898 486346 374134
rect 486582 373898 514026 374134
rect 514262 373898 514346 374134
rect 514582 373898 542026 374134
rect 542262 373898 542346 374134
rect 542582 373898 570026 374134
rect 570262 373898 570346 374134
rect 570582 373898 586302 374134
rect 586538 373898 586622 374134
rect 586858 373898 592650 374134
rect -8726 373866 592650 373898
rect -8726 350829 592650 350861
rect -8726 350593 -1974 350829
rect -1738 350593 -1654 350829
rect -1418 350593 41526 350829
rect 41762 350593 41846 350829
rect 42082 350593 69526 350829
rect 69762 350593 69846 350829
rect 70082 350593 97526 350829
rect 97762 350593 97846 350829
rect 98082 350593 125526 350829
rect 125762 350593 125846 350829
rect 126082 350593 153526 350829
rect 153762 350593 153846 350829
rect 154082 350593 181526 350829
rect 181762 350593 181846 350829
rect 182082 350593 209526 350829
rect 209762 350593 209846 350829
rect 210082 350593 237526 350829
rect 237762 350593 237846 350829
rect 238082 350593 265526 350829
rect 265762 350593 265846 350829
rect 266082 350593 293526 350829
rect 293762 350593 293846 350829
rect 294082 350593 321526 350829
rect 321762 350593 321846 350829
rect 322082 350593 349526 350829
rect 349762 350593 349846 350829
rect 350082 350593 377526 350829
rect 377762 350593 377846 350829
rect 378082 350593 405526 350829
rect 405762 350593 405846 350829
rect 406082 350593 433526 350829
rect 433762 350593 433846 350829
rect 434082 350593 461526 350829
rect 461762 350593 461846 350829
rect 462082 350593 489526 350829
rect 489762 350593 489846 350829
rect 490082 350593 517526 350829
rect 517762 350593 517846 350829
rect 518082 350593 545526 350829
rect 545762 350593 545846 350829
rect 546082 350593 573526 350829
rect 573762 350593 573846 350829
rect 574082 350593 585342 350829
rect 585578 350593 585662 350829
rect 585898 350593 592650 350829
rect -8726 350509 592650 350593
rect -8726 350273 -1974 350509
rect -1738 350273 -1654 350509
rect -1418 350273 41526 350509
rect 41762 350273 41846 350509
rect 42082 350273 69526 350509
rect 69762 350273 69846 350509
rect 70082 350273 97526 350509
rect 97762 350273 97846 350509
rect 98082 350273 125526 350509
rect 125762 350273 125846 350509
rect 126082 350273 153526 350509
rect 153762 350273 153846 350509
rect 154082 350273 181526 350509
rect 181762 350273 181846 350509
rect 182082 350273 209526 350509
rect 209762 350273 209846 350509
rect 210082 350273 237526 350509
rect 237762 350273 237846 350509
rect 238082 350273 265526 350509
rect 265762 350273 265846 350509
rect 266082 350273 293526 350509
rect 293762 350273 293846 350509
rect 294082 350273 321526 350509
rect 321762 350273 321846 350509
rect 322082 350273 349526 350509
rect 349762 350273 349846 350509
rect 350082 350273 377526 350509
rect 377762 350273 377846 350509
rect 378082 350273 405526 350509
rect 405762 350273 405846 350509
rect 406082 350273 433526 350509
rect 433762 350273 433846 350509
rect 434082 350273 461526 350509
rect 461762 350273 461846 350509
rect 462082 350273 489526 350509
rect 489762 350273 489846 350509
rect 490082 350273 517526 350509
rect 517762 350273 517846 350509
rect 518082 350273 545526 350509
rect 545762 350273 545846 350509
rect 546082 350273 573526 350509
rect 573762 350273 573846 350509
rect 574082 350273 585342 350509
rect 585578 350273 585662 350509
rect 585898 350273 592650 350509
rect -8726 350241 592650 350273
rect -8726 347454 592650 347486
rect -8726 347218 -2934 347454
rect -2698 347218 -2614 347454
rect -2378 347218 38026 347454
rect 38262 347218 38346 347454
rect 38582 347218 66026 347454
rect 66262 347218 66346 347454
rect 66582 347218 94026 347454
rect 94262 347218 94346 347454
rect 94582 347218 122026 347454
rect 122262 347218 122346 347454
rect 122582 347218 150026 347454
rect 150262 347218 150346 347454
rect 150582 347218 178026 347454
rect 178262 347218 178346 347454
rect 178582 347218 206026 347454
rect 206262 347218 206346 347454
rect 206582 347218 234026 347454
rect 234262 347218 234346 347454
rect 234582 347218 262026 347454
rect 262262 347218 262346 347454
rect 262582 347218 290026 347454
rect 290262 347218 290346 347454
rect 290582 347218 318026 347454
rect 318262 347218 318346 347454
rect 318582 347218 346026 347454
rect 346262 347218 346346 347454
rect 346582 347218 374026 347454
rect 374262 347218 374346 347454
rect 374582 347218 402026 347454
rect 402262 347218 402346 347454
rect 402582 347218 430026 347454
rect 430262 347218 430346 347454
rect 430582 347218 458026 347454
rect 458262 347218 458346 347454
rect 458582 347218 486026 347454
rect 486262 347218 486346 347454
rect 486582 347218 514026 347454
rect 514262 347218 514346 347454
rect 514582 347218 542026 347454
rect 542262 347218 542346 347454
rect 542582 347218 570026 347454
rect 570262 347218 570346 347454
rect 570582 347218 586302 347454
rect 586538 347218 586622 347454
rect 586858 347218 592650 347454
rect -8726 347134 592650 347218
rect -8726 346898 -2934 347134
rect -2698 346898 -2614 347134
rect -2378 346898 38026 347134
rect 38262 346898 38346 347134
rect 38582 346898 66026 347134
rect 66262 346898 66346 347134
rect 66582 346898 94026 347134
rect 94262 346898 94346 347134
rect 94582 346898 122026 347134
rect 122262 346898 122346 347134
rect 122582 346898 150026 347134
rect 150262 346898 150346 347134
rect 150582 346898 178026 347134
rect 178262 346898 178346 347134
rect 178582 346898 206026 347134
rect 206262 346898 206346 347134
rect 206582 346898 234026 347134
rect 234262 346898 234346 347134
rect 234582 346898 262026 347134
rect 262262 346898 262346 347134
rect 262582 346898 290026 347134
rect 290262 346898 290346 347134
rect 290582 346898 318026 347134
rect 318262 346898 318346 347134
rect 318582 346898 346026 347134
rect 346262 346898 346346 347134
rect 346582 346898 374026 347134
rect 374262 346898 374346 347134
rect 374582 346898 402026 347134
rect 402262 346898 402346 347134
rect 402582 346898 430026 347134
rect 430262 346898 430346 347134
rect 430582 346898 458026 347134
rect 458262 346898 458346 347134
rect 458582 346898 486026 347134
rect 486262 346898 486346 347134
rect 486582 346898 514026 347134
rect 514262 346898 514346 347134
rect 514582 346898 542026 347134
rect 542262 346898 542346 347134
rect 542582 346898 570026 347134
rect 570262 346898 570346 347134
rect 570582 346898 586302 347134
rect 586538 346898 586622 347134
rect 586858 346898 592650 347134
rect -8726 346866 592650 346898
rect -8726 323829 592650 323861
rect -8726 323593 -1974 323829
rect -1738 323593 -1654 323829
rect -1418 323593 41526 323829
rect 41762 323593 41846 323829
rect 42082 323593 69526 323829
rect 69762 323593 69846 323829
rect 70082 323593 97526 323829
rect 97762 323593 97846 323829
rect 98082 323593 125526 323829
rect 125762 323593 125846 323829
rect 126082 323593 153526 323829
rect 153762 323593 153846 323829
rect 154082 323593 181526 323829
rect 181762 323593 181846 323829
rect 182082 323593 209526 323829
rect 209762 323593 209846 323829
rect 210082 323593 237526 323829
rect 237762 323593 237846 323829
rect 238082 323593 265526 323829
rect 265762 323593 265846 323829
rect 266082 323593 293526 323829
rect 293762 323593 293846 323829
rect 294082 323593 321526 323829
rect 321762 323593 321846 323829
rect 322082 323593 349526 323829
rect 349762 323593 349846 323829
rect 350082 323593 377526 323829
rect 377762 323593 377846 323829
rect 378082 323593 405526 323829
rect 405762 323593 405846 323829
rect 406082 323593 433526 323829
rect 433762 323593 433846 323829
rect 434082 323593 461526 323829
rect 461762 323593 461846 323829
rect 462082 323593 489526 323829
rect 489762 323593 489846 323829
rect 490082 323593 517526 323829
rect 517762 323593 517846 323829
rect 518082 323593 545526 323829
rect 545762 323593 545846 323829
rect 546082 323593 573526 323829
rect 573762 323593 573846 323829
rect 574082 323593 585342 323829
rect 585578 323593 585662 323829
rect 585898 323593 592650 323829
rect -8726 323509 592650 323593
rect -8726 323273 -1974 323509
rect -1738 323273 -1654 323509
rect -1418 323273 41526 323509
rect 41762 323273 41846 323509
rect 42082 323273 69526 323509
rect 69762 323273 69846 323509
rect 70082 323273 97526 323509
rect 97762 323273 97846 323509
rect 98082 323273 125526 323509
rect 125762 323273 125846 323509
rect 126082 323273 153526 323509
rect 153762 323273 153846 323509
rect 154082 323273 181526 323509
rect 181762 323273 181846 323509
rect 182082 323273 209526 323509
rect 209762 323273 209846 323509
rect 210082 323273 237526 323509
rect 237762 323273 237846 323509
rect 238082 323273 265526 323509
rect 265762 323273 265846 323509
rect 266082 323273 293526 323509
rect 293762 323273 293846 323509
rect 294082 323273 321526 323509
rect 321762 323273 321846 323509
rect 322082 323273 349526 323509
rect 349762 323273 349846 323509
rect 350082 323273 377526 323509
rect 377762 323273 377846 323509
rect 378082 323273 405526 323509
rect 405762 323273 405846 323509
rect 406082 323273 433526 323509
rect 433762 323273 433846 323509
rect 434082 323273 461526 323509
rect 461762 323273 461846 323509
rect 462082 323273 489526 323509
rect 489762 323273 489846 323509
rect 490082 323273 517526 323509
rect 517762 323273 517846 323509
rect 518082 323273 545526 323509
rect 545762 323273 545846 323509
rect 546082 323273 573526 323509
rect 573762 323273 573846 323509
rect 574082 323273 585342 323509
rect 585578 323273 585662 323509
rect 585898 323273 592650 323509
rect -8726 323241 592650 323273
rect -8726 320454 592650 320486
rect -8726 320218 -2934 320454
rect -2698 320218 -2614 320454
rect -2378 320218 38026 320454
rect 38262 320218 38346 320454
rect 38582 320218 66026 320454
rect 66262 320218 66346 320454
rect 66582 320218 94026 320454
rect 94262 320218 94346 320454
rect 94582 320218 122026 320454
rect 122262 320218 122346 320454
rect 122582 320218 150026 320454
rect 150262 320218 150346 320454
rect 150582 320218 178026 320454
rect 178262 320218 178346 320454
rect 178582 320218 206026 320454
rect 206262 320218 206346 320454
rect 206582 320218 234026 320454
rect 234262 320218 234346 320454
rect 234582 320218 262026 320454
rect 262262 320218 262346 320454
rect 262582 320218 290026 320454
rect 290262 320218 290346 320454
rect 290582 320218 318026 320454
rect 318262 320218 318346 320454
rect 318582 320218 346026 320454
rect 346262 320218 346346 320454
rect 346582 320218 374026 320454
rect 374262 320218 374346 320454
rect 374582 320218 402026 320454
rect 402262 320218 402346 320454
rect 402582 320218 430026 320454
rect 430262 320218 430346 320454
rect 430582 320218 458026 320454
rect 458262 320218 458346 320454
rect 458582 320218 486026 320454
rect 486262 320218 486346 320454
rect 486582 320218 514026 320454
rect 514262 320218 514346 320454
rect 514582 320218 542026 320454
rect 542262 320218 542346 320454
rect 542582 320218 570026 320454
rect 570262 320218 570346 320454
rect 570582 320218 586302 320454
rect 586538 320218 586622 320454
rect 586858 320218 592650 320454
rect -8726 320134 592650 320218
rect -8726 319898 -2934 320134
rect -2698 319898 -2614 320134
rect -2378 319898 38026 320134
rect 38262 319898 38346 320134
rect 38582 319898 66026 320134
rect 66262 319898 66346 320134
rect 66582 319898 94026 320134
rect 94262 319898 94346 320134
rect 94582 319898 122026 320134
rect 122262 319898 122346 320134
rect 122582 319898 150026 320134
rect 150262 319898 150346 320134
rect 150582 319898 178026 320134
rect 178262 319898 178346 320134
rect 178582 319898 206026 320134
rect 206262 319898 206346 320134
rect 206582 319898 234026 320134
rect 234262 319898 234346 320134
rect 234582 319898 262026 320134
rect 262262 319898 262346 320134
rect 262582 319898 290026 320134
rect 290262 319898 290346 320134
rect 290582 319898 318026 320134
rect 318262 319898 318346 320134
rect 318582 319898 346026 320134
rect 346262 319898 346346 320134
rect 346582 319898 374026 320134
rect 374262 319898 374346 320134
rect 374582 319898 402026 320134
rect 402262 319898 402346 320134
rect 402582 319898 430026 320134
rect 430262 319898 430346 320134
rect 430582 319898 458026 320134
rect 458262 319898 458346 320134
rect 458582 319898 486026 320134
rect 486262 319898 486346 320134
rect 486582 319898 514026 320134
rect 514262 319898 514346 320134
rect 514582 319898 542026 320134
rect 542262 319898 542346 320134
rect 542582 319898 570026 320134
rect 570262 319898 570346 320134
rect 570582 319898 586302 320134
rect 586538 319898 586622 320134
rect 586858 319898 592650 320134
rect -8726 319866 592650 319898
rect -8726 296829 592650 296861
rect -8726 296593 -1974 296829
rect -1738 296593 -1654 296829
rect -1418 296593 41526 296829
rect 41762 296593 41846 296829
rect 42082 296593 69526 296829
rect 69762 296593 69846 296829
rect 70082 296593 97526 296829
rect 97762 296593 97846 296829
rect 98082 296593 125526 296829
rect 125762 296593 125846 296829
rect 126082 296593 153526 296829
rect 153762 296593 153846 296829
rect 154082 296593 181526 296829
rect 181762 296593 181846 296829
rect 182082 296593 209526 296829
rect 209762 296593 209846 296829
rect 210082 296593 237526 296829
rect 237762 296593 237846 296829
rect 238082 296593 265526 296829
rect 265762 296593 265846 296829
rect 266082 296593 293526 296829
rect 293762 296593 293846 296829
rect 294082 296593 321526 296829
rect 321762 296593 321846 296829
rect 322082 296593 349526 296829
rect 349762 296593 349846 296829
rect 350082 296593 377526 296829
rect 377762 296593 377846 296829
rect 378082 296593 405526 296829
rect 405762 296593 405846 296829
rect 406082 296593 433526 296829
rect 433762 296593 433846 296829
rect 434082 296593 461526 296829
rect 461762 296593 461846 296829
rect 462082 296593 489526 296829
rect 489762 296593 489846 296829
rect 490082 296593 517526 296829
rect 517762 296593 517846 296829
rect 518082 296593 545526 296829
rect 545762 296593 545846 296829
rect 546082 296593 573526 296829
rect 573762 296593 573846 296829
rect 574082 296593 585342 296829
rect 585578 296593 585662 296829
rect 585898 296593 592650 296829
rect -8726 296509 592650 296593
rect -8726 296273 -1974 296509
rect -1738 296273 -1654 296509
rect -1418 296273 41526 296509
rect 41762 296273 41846 296509
rect 42082 296273 69526 296509
rect 69762 296273 69846 296509
rect 70082 296273 97526 296509
rect 97762 296273 97846 296509
rect 98082 296273 125526 296509
rect 125762 296273 125846 296509
rect 126082 296273 153526 296509
rect 153762 296273 153846 296509
rect 154082 296273 181526 296509
rect 181762 296273 181846 296509
rect 182082 296273 209526 296509
rect 209762 296273 209846 296509
rect 210082 296273 237526 296509
rect 237762 296273 237846 296509
rect 238082 296273 265526 296509
rect 265762 296273 265846 296509
rect 266082 296273 293526 296509
rect 293762 296273 293846 296509
rect 294082 296273 321526 296509
rect 321762 296273 321846 296509
rect 322082 296273 349526 296509
rect 349762 296273 349846 296509
rect 350082 296273 377526 296509
rect 377762 296273 377846 296509
rect 378082 296273 405526 296509
rect 405762 296273 405846 296509
rect 406082 296273 433526 296509
rect 433762 296273 433846 296509
rect 434082 296273 461526 296509
rect 461762 296273 461846 296509
rect 462082 296273 489526 296509
rect 489762 296273 489846 296509
rect 490082 296273 517526 296509
rect 517762 296273 517846 296509
rect 518082 296273 545526 296509
rect 545762 296273 545846 296509
rect 546082 296273 573526 296509
rect 573762 296273 573846 296509
rect 574082 296273 585342 296509
rect 585578 296273 585662 296509
rect 585898 296273 592650 296509
rect -8726 296241 592650 296273
rect -8726 293454 592650 293486
rect -8726 293218 -2934 293454
rect -2698 293218 -2614 293454
rect -2378 293218 38026 293454
rect 38262 293218 38346 293454
rect 38582 293218 66026 293454
rect 66262 293218 66346 293454
rect 66582 293218 94026 293454
rect 94262 293218 94346 293454
rect 94582 293218 122026 293454
rect 122262 293218 122346 293454
rect 122582 293218 150026 293454
rect 150262 293218 150346 293454
rect 150582 293218 178026 293454
rect 178262 293218 178346 293454
rect 178582 293218 206026 293454
rect 206262 293218 206346 293454
rect 206582 293218 234026 293454
rect 234262 293218 234346 293454
rect 234582 293218 262026 293454
rect 262262 293218 262346 293454
rect 262582 293218 290026 293454
rect 290262 293218 290346 293454
rect 290582 293218 318026 293454
rect 318262 293218 318346 293454
rect 318582 293218 346026 293454
rect 346262 293218 346346 293454
rect 346582 293218 374026 293454
rect 374262 293218 374346 293454
rect 374582 293218 402026 293454
rect 402262 293218 402346 293454
rect 402582 293218 430026 293454
rect 430262 293218 430346 293454
rect 430582 293218 458026 293454
rect 458262 293218 458346 293454
rect 458582 293218 486026 293454
rect 486262 293218 486346 293454
rect 486582 293218 514026 293454
rect 514262 293218 514346 293454
rect 514582 293218 542026 293454
rect 542262 293218 542346 293454
rect 542582 293218 570026 293454
rect 570262 293218 570346 293454
rect 570582 293218 586302 293454
rect 586538 293218 586622 293454
rect 586858 293218 592650 293454
rect -8726 293134 592650 293218
rect -8726 292898 -2934 293134
rect -2698 292898 -2614 293134
rect -2378 292898 38026 293134
rect 38262 292898 38346 293134
rect 38582 292898 66026 293134
rect 66262 292898 66346 293134
rect 66582 292898 94026 293134
rect 94262 292898 94346 293134
rect 94582 292898 122026 293134
rect 122262 292898 122346 293134
rect 122582 292898 150026 293134
rect 150262 292898 150346 293134
rect 150582 292898 178026 293134
rect 178262 292898 178346 293134
rect 178582 292898 206026 293134
rect 206262 292898 206346 293134
rect 206582 292898 234026 293134
rect 234262 292898 234346 293134
rect 234582 292898 262026 293134
rect 262262 292898 262346 293134
rect 262582 292898 290026 293134
rect 290262 292898 290346 293134
rect 290582 292898 318026 293134
rect 318262 292898 318346 293134
rect 318582 292898 346026 293134
rect 346262 292898 346346 293134
rect 346582 292898 374026 293134
rect 374262 292898 374346 293134
rect 374582 292898 402026 293134
rect 402262 292898 402346 293134
rect 402582 292898 430026 293134
rect 430262 292898 430346 293134
rect 430582 292898 458026 293134
rect 458262 292898 458346 293134
rect 458582 292898 486026 293134
rect 486262 292898 486346 293134
rect 486582 292898 514026 293134
rect 514262 292898 514346 293134
rect 514582 292898 542026 293134
rect 542262 292898 542346 293134
rect 542582 292898 570026 293134
rect 570262 292898 570346 293134
rect 570582 292898 586302 293134
rect 586538 292898 586622 293134
rect 586858 292898 592650 293134
rect -8726 292866 592650 292898
rect -8726 269829 592650 269861
rect -8726 269593 -1974 269829
rect -1738 269593 -1654 269829
rect -1418 269593 41526 269829
rect 41762 269593 41846 269829
rect 42082 269593 69526 269829
rect 69762 269593 69846 269829
rect 70082 269593 97526 269829
rect 97762 269593 97846 269829
rect 98082 269593 125526 269829
rect 125762 269593 125846 269829
rect 126082 269593 153526 269829
rect 153762 269593 153846 269829
rect 154082 269593 181526 269829
rect 181762 269593 181846 269829
rect 182082 269593 209526 269829
rect 209762 269593 209846 269829
rect 210082 269593 237526 269829
rect 237762 269593 237846 269829
rect 238082 269593 265526 269829
rect 265762 269593 265846 269829
rect 266082 269593 293526 269829
rect 293762 269593 293846 269829
rect 294082 269593 321526 269829
rect 321762 269593 321846 269829
rect 322082 269593 349526 269829
rect 349762 269593 349846 269829
rect 350082 269593 377526 269829
rect 377762 269593 377846 269829
rect 378082 269593 405526 269829
rect 405762 269593 405846 269829
rect 406082 269593 433526 269829
rect 433762 269593 433846 269829
rect 434082 269593 461526 269829
rect 461762 269593 461846 269829
rect 462082 269593 489526 269829
rect 489762 269593 489846 269829
rect 490082 269593 517526 269829
rect 517762 269593 517846 269829
rect 518082 269593 545526 269829
rect 545762 269593 545846 269829
rect 546082 269593 573526 269829
rect 573762 269593 573846 269829
rect 574082 269593 585342 269829
rect 585578 269593 585662 269829
rect 585898 269593 592650 269829
rect -8726 269509 592650 269593
rect -8726 269273 -1974 269509
rect -1738 269273 -1654 269509
rect -1418 269273 41526 269509
rect 41762 269273 41846 269509
rect 42082 269273 69526 269509
rect 69762 269273 69846 269509
rect 70082 269273 97526 269509
rect 97762 269273 97846 269509
rect 98082 269273 125526 269509
rect 125762 269273 125846 269509
rect 126082 269273 153526 269509
rect 153762 269273 153846 269509
rect 154082 269273 181526 269509
rect 181762 269273 181846 269509
rect 182082 269273 209526 269509
rect 209762 269273 209846 269509
rect 210082 269273 237526 269509
rect 237762 269273 237846 269509
rect 238082 269273 265526 269509
rect 265762 269273 265846 269509
rect 266082 269273 293526 269509
rect 293762 269273 293846 269509
rect 294082 269273 321526 269509
rect 321762 269273 321846 269509
rect 322082 269273 349526 269509
rect 349762 269273 349846 269509
rect 350082 269273 377526 269509
rect 377762 269273 377846 269509
rect 378082 269273 405526 269509
rect 405762 269273 405846 269509
rect 406082 269273 433526 269509
rect 433762 269273 433846 269509
rect 434082 269273 461526 269509
rect 461762 269273 461846 269509
rect 462082 269273 489526 269509
rect 489762 269273 489846 269509
rect 490082 269273 517526 269509
rect 517762 269273 517846 269509
rect 518082 269273 545526 269509
rect 545762 269273 545846 269509
rect 546082 269273 573526 269509
rect 573762 269273 573846 269509
rect 574082 269273 585342 269509
rect 585578 269273 585662 269509
rect 585898 269273 592650 269509
rect -8726 269241 592650 269273
rect -8726 266454 592650 266486
rect -8726 266218 -2934 266454
rect -2698 266218 -2614 266454
rect -2378 266218 38026 266454
rect 38262 266218 38346 266454
rect 38582 266218 66026 266454
rect 66262 266218 66346 266454
rect 66582 266218 94026 266454
rect 94262 266218 94346 266454
rect 94582 266218 122026 266454
rect 122262 266218 122346 266454
rect 122582 266218 150026 266454
rect 150262 266218 150346 266454
rect 150582 266218 178026 266454
rect 178262 266218 178346 266454
rect 178582 266218 206026 266454
rect 206262 266218 206346 266454
rect 206582 266218 234026 266454
rect 234262 266218 234346 266454
rect 234582 266218 262026 266454
rect 262262 266218 262346 266454
rect 262582 266218 290026 266454
rect 290262 266218 290346 266454
rect 290582 266218 318026 266454
rect 318262 266218 318346 266454
rect 318582 266218 346026 266454
rect 346262 266218 346346 266454
rect 346582 266218 374026 266454
rect 374262 266218 374346 266454
rect 374582 266218 402026 266454
rect 402262 266218 402346 266454
rect 402582 266218 430026 266454
rect 430262 266218 430346 266454
rect 430582 266218 458026 266454
rect 458262 266218 458346 266454
rect 458582 266218 486026 266454
rect 486262 266218 486346 266454
rect 486582 266218 514026 266454
rect 514262 266218 514346 266454
rect 514582 266218 542026 266454
rect 542262 266218 542346 266454
rect 542582 266218 570026 266454
rect 570262 266218 570346 266454
rect 570582 266218 586302 266454
rect 586538 266218 586622 266454
rect 586858 266218 592650 266454
rect -8726 266134 592650 266218
rect -8726 265898 -2934 266134
rect -2698 265898 -2614 266134
rect -2378 265898 38026 266134
rect 38262 265898 38346 266134
rect 38582 265898 66026 266134
rect 66262 265898 66346 266134
rect 66582 265898 94026 266134
rect 94262 265898 94346 266134
rect 94582 265898 122026 266134
rect 122262 265898 122346 266134
rect 122582 265898 150026 266134
rect 150262 265898 150346 266134
rect 150582 265898 178026 266134
rect 178262 265898 178346 266134
rect 178582 265898 206026 266134
rect 206262 265898 206346 266134
rect 206582 265898 234026 266134
rect 234262 265898 234346 266134
rect 234582 265898 262026 266134
rect 262262 265898 262346 266134
rect 262582 265898 290026 266134
rect 290262 265898 290346 266134
rect 290582 265898 318026 266134
rect 318262 265898 318346 266134
rect 318582 265898 346026 266134
rect 346262 265898 346346 266134
rect 346582 265898 374026 266134
rect 374262 265898 374346 266134
rect 374582 265898 402026 266134
rect 402262 265898 402346 266134
rect 402582 265898 430026 266134
rect 430262 265898 430346 266134
rect 430582 265898 458026 266134
rect 458262 265898 458346 266134
rect 458582 265898 486026 266134
rect 486262 265898 486346 266134
rect 486582 265898 514026 266134
rect 514262 265898 514346 266134
rect 514582 265898 542026 266134
rect 542262 265898 542346 266134
rect 542582 265898 570026 266134
rect 570262 265898 570346 266134
rect 570582 265898 586302 266134
rect 586538 265898 586622 266134
rect 586858 265898 592650 266134
rect -8726 265866 592650 265898
rect -8726 242829 592650 242861
rect -8726 242593 -1974 242829
rect -1738 242593 -1654 242829
rect -1418 242593 41526 242829
rect 41762 242593 41846 242829
rect 42082 242593 69526 242829
rect 69762 242593 69846 242829
rect 70082 242593 97526 242829
rect 97762 242593 97846 242829
rect 98082 242593 125526 242829
rect 125762 242593 125846 242829
rect 126082 242593 153526 242829
rect 153762 242593 153846 242829
rect 154082 242593 181526 242829
rect 181762 242593 181846 242829
rect 182082 242593 209526 242829
rect 209762 242593 209846 242829
rect 210082 242593 237526 242829
rect 237762 242593 237846 242829
rect 238082 242593 265526 242829
rect 265762 242593 265846 242829
rect 266082 242593 293526 242829
rect 293762 242593 293846 242829
rect 294082 242593 321526 242829
rect 321762 242593 321846 242829
rect 322082 242593 349526 242829
rect 349762 242593 349846 242829
rect 350082 242593 377526 242829
rect 377762 242593 377846 242829
rect 378082 242593 405526 242829
rect 405762 242593 405846 242829
rect 406082 242593 433526 242829
rect 433762 242593 433846 242829
rect 434082 242593 461526 242829
rect 461762 242593 461846 242829
rect 462082 242593 489526 242829
rect 489762 242593 489846 242829
rect 490082 242593 517526 242829
rect 517762 242593 517846 242829
rect 518082 242593 545526 242829
rect 545762 242593 545846 242829
rect 546082 242593 573526 242829
rect 573762 242593 573846 242829
rect 574082 242593 585342 242829
rect 585578 242593 585662 242829
rect 585898 242593 592650 242829
rect -8726 242509 592650 242593
rect -8726 242273 -1974 242509
rect -1738 242273 -1654 242509
rect -1418 242273 41526 242509
rect 41762 242273 41846 242509
rect 42082 242273 69526 242509
rect 69762 242273 69846 242509
rect 70082 242273 97526 242509
rect 97762 242273 97846 242509
rect 98082 242273 125526 242509
rect 125762 242273 125846 242509
rect 126082 242273 153526 242509
rect 153762 242273 153846 242509
rect 154082 242273 181526 242509
rect 181762 242273 181846 242509
rect 182082 242273 209526 242509
rect 209762 242273 209846 242509
rect 210082 242273 237526 242509
rect 237762 242273 237846 242509
rect 238082 242273 265526 242509
rect 265762 242273 265846 242509
rect 266082 242273 293526 242509
rect 293762 242273 293846 242509
rect 294082 242273 321526 242509
rect 321762 242273 321846 242509
rect 322082 242273 349526 242509
rect 349762 242273 349846 242509
rect 350082 242273 377526 242509
rect 377762 242273 377846 242509
rect 378082 242273 405526 242509
rect 405762 242273 405846 242509
rect 406082 242273 433526 242509
rect 433762 242273 433846 242509
rect 434082 242273 461526 242509
rect 461762 242273 461846 242509
rect 462082 242273 489526 242509
rect 489762 242273 489846 242509
rect 490082 242273 517526 242509
rect 517762 242273 517846 242509
rect 518082 242273 545526 242509
rect 545762 242273 545846 242509
rect 546082 242273 573526 242509
rect 573762 242273 573846 242509
rect 574082 242273 585342 242509
rect 585578 242273 585662 242509
rect 585898 242273 592650 242509
rect -8726 242241 592650 242273
rect -8726 239454 592650 239486
rect -8726 239218 -2934 239454
rect -2698 239218 -2614 239454
rect -2378 239218 38026 239454
rect 38262 239218 38346 239454
rect 38582 239218 66026 239454
rect 66262 239218 66346 239454
rect 66582 239218 94026 239454
rect 94262 239218 94346 239454
rect 94582 239218 122026 239454
rect 122262 239218 122346 239454
rect 122582 239218 150026 239454
rect 150262 239218 150346 239454
rect 150582 239218 178026 239454
rect 178262 239218 178346 239454
rect 178582 239218 206026 239454
rect 206262 239218 206346 239454
rect 206582 239218 234026 239454
rect 234262 239218 234346 239454
rect 234582 239218 262026 239454
rect 262262 239218 262346 239454
rect 262582 239218 290026 239454
rect 290262 239218 290346 239454
rect 290582 239218 318026 239454
rect 318262 239218 318346 239454
rect 318582 239218 346026 239454
rect 346262 239218 346346 239454
rect 346582 239218 374026 239454
rect 374262 239218 374346 239454
rect 374582 239218 402026 239454
rect 402262 239218 402346 239454
rect 402582 239218 430026 239454
rect 430262 239218 430346 239454
rect 430582 239218 458026 239454
rect 458262 239218 458346 239454
rect 458582 239218 486026 239454
rect 486262 239218 486346 239454
rect 486582 239218 514026 239454
rect 514262 239218 514346 239454
rect 514582 239218 542026 239454
rect 542262 239218 542346 239454
rect 542582 239218 570026 239454
rect 570262 239218 570346 239454
rect 570582 239218 586302 239454
rect 586538 239218 586622 239454
rect 586858 239218 592650 239454
rect -8726 239134 592650 239218
rect -8726 238898 -2934 239134
rect -2698 238898 -2614 239134
rect -2378 238898 38026 239134
rect 38262 238898 38346 239134
rect 38582 238898 66026 239134
rect 66262 238898 66346 239134
rect 66582 238898 94026 239134
rect 94262 238898 94346 239134
rect 94582 238898 122026 239134
rect 122262 238898 122346 239134
rect 122582 238898 150026 239134
rect 150262 238898 150346 239134
rect 150582 238898 178026 239134
rect 178262 238898 178346 239134
rect 178582 238898 206026 239134
rect 206262 238898 206346 239134
rect 206582 238898 234026 239134
rect 234262 238898 234346 239134
rect 234582 238898 262026 239134
rect 262262 238898 262346 239134
rect 262582 238898 290026 239134
rect 290262 238898 290346 239134
rect 290582 238898 318026 239134
rect 318262 238898 318346 239134
rect 318582 238898 346026 239134
rect 346262 238898 346346 239134
rect 346582 238898 374026 239134
rect 374262 238898 374346 239134
rect 374582 238898 402026 239134
rect 402262 238898 402346 239134
rect 402582 238898 430026 239134
rect 430262 238898 430346 239134
rect 430582 238898 458026 239134
rect 458262 238898 458346 239134
rect 458582 238898 486026 239134
rect 486262 238898 486346 239134
rect 486582 238898 514026 239134
rect 514262 238898 514346 239134
rect 514582 238898 542026 239134
rect 542262 238898 542346 239134
rect 542582 238898 570026 239134
rect 570262 238898 570346 239134
rect 570582 238898 586302 239134
rect 586538 238898 586622 239134
rect 586858 238898 592650 239134
rect -8726 238866 592650 238898
rect -8726 215829 592650 215861
rect -8726 215593 -1974 215829
rect -1738 215593 -1654 215829
rect -1418 215593 41526 215829
rect 41762 215593 41846 215829
rect 42082 215593 69526 215829
rect 69762 215593 69846 215829
rect 70082 215593 97526 215829
rect 97762 215593 97846 215829
rect 98082 215593 125526 215829
rect 125762 215593 125846 215829
rect 126082 215593 153526 215829
rect 153762 215593 153846 215829
rect 154082 215593 181526 215829
rect 181762 215593 181846 215829
rect 182082 215593 209526 215829
rect 209762 215593 209846 215829
rect 210082 215593 237526 215829
rect 237762 215593 237846 215829
rect 238082 215593 265526 215829
rect 265762 215593 265846 215829
rect 266082 215593 293526 215829
rect 293762 215593 293846 215829
rect 294082 215593 321526 215829
rect 321762 215593 321846 215829
rect 322082 215593 349526 215829
rect 349762 215593 349846 215829
rect 350082 215593 377526 215829
rect 377762 215593 377846 215829
rect 378082 215593 405526 215829
rect 405762 215593 405846 215829
rect 406082 215593 433526 215829
rect 433762 215593 433846 215829
rect 434082 215593 461526 215829
rect 461762 215593 461846 215829
rect 462082 215593 489526 215829
rect 489762 215593 489846 215829
rect 490082 215593 517526 215829
rect 517762 215593 517846 215829
rect 518082 215593 545526 215829
rect 545762 215593 545846 215829
rect 546082 215593 573526 215829
rect 573762 215593 573846 215829
rect 574082 215593 585342 215829
rect 585578 215593 585662 215829
rect 585898 215593 592650 215829
rect -8726 215509 592650 215593
rect -8726 215273 -1974 215509
rect -1738 215273 -1654 215509
rect -1418 215273 41526 215509
rect 41762 215273 41846 215509
rect 42082 215273 69526 215509
rect 69762 215273 69846 215509
rect 70082 215273 97526 215509
rect 97762 215273 97846 215509
rect 98082 215273 125526 215509
rect 125762 215273 125846 215509
rect 126082 215273 153526 215509
rect 153762 215273 153846 215509
rect 154082 215273 181526 215509
rect 181762 215273 181846 215509
rect 182082 215273 209526 215509
rect 209762 215273 209846 215509
rect 210082 215273 237526 215509
rect 237762 215273 237846 215509
rect 238082 215273 265526 215509
rect 265762 215273 265846 215509
rect 266082 215273 293526 215509
rect 293762 215273 293846 215509
rect 294082 215273 321526 215509
rect 321762 215273 321846 215509
rect 322082 215273 349526 215509
rect 349762 215273 349846 215509
rect 350082 215273 377526 215509
rect 377762 215273 377846 215509
rect 378082 215273 405526 215509
rect 405762 215273 405846 215509
rect 406082 215273 433526 215509
rect 433762 215273 433846 215509
rect 434082 215273 461526 215509
rect 461762 215273 461846 215509
rect 462082 215273 489526 215509
rect 489762 215273 489846 215509
rect 490082 215273 517526 215509
rect 517762 215273 517846 215509
rect 518082 215273 545526 215509
rect 545762 215273 545846 215509
rect 546082 215273 573526 215509
rect 573762 215273 573846 215509
rect 574082 215273 585342 215509
rect 585578 215273 585662 215509
rect 585898 215273 592650 215509
rect -8726 215241 592650 215273
rect -8726 212454 592650 212486
rect -8726 212218 -2934 212454
rect -2698 212218 -2614 212454
rect -2378 212218 38026 212454
rect 38262 212218 38346 212454
rect 38582 212218 66026 212454
rect 66262 212218 66346 212454
rect 66582 212218 94026 212454
rect 94262 212218 94346 212454
rect 94582 212218 122026 212454
rect 122262 212218 122346 212454
rect 122582 212218 150026 212454
rect 150262 212218 150346 212454
rect 150582 212218 178026 212454
rect 178262 212218 178346 212454
rect 178582 212218 206026 212454
rect 206262 212218 206346 212454
rect 206582 212218 234026 212454
rect 234262 212218 234346 212454
rect 234582 212218 262026 212454
rect 262262 212218 262346 212454
rect 262582 212218 290026 212454
rect 290262 212218 290346 212454
rect 290582 212218 318026 212454
rect 318262 212218 318346 212454
rect 318582 212218 346026 212454
rect 346262 212218 346346 212454
rect 346582 212218 374026 212454
rect 374262 212218 374346 212454
rect 374582 212218 402026 212454
rect 402262 212218 402346 212454
rect 402582 212218 430026 212454
rect 430262 212218 430346 212454
rect 430582 212218 458026 212454
rect 458262 212218 458346 212454
rect 458582 212218 486026 212454
rect 486262 212218 486346 212454
rect 486582 212218 514026 212454
rect 514262 212218 514346 212454
rect 514582 212218 542026 212454
rect 542262 212218 542346 212454
rect 542582 212218 570026 212454
rect 570262 212218 570346 212454
rect 570582 212218 586302 212454
rect 586538 212218 586622 212454
rect 586858 212218 592650 212454
rect -8726 212134 592650 212218
rect -8726 211898 -2934 212134
rect -2698 211898 -2614 212134
rect -2378 211898 38026 212134
rect 38262 211898 38346 212134
rect 38582 211898 66026 212134
rect 66262 211898 66346 212134
rect 66582 211898 94026 212134
rect 94262 211898 94346 212134
rect 94582 211898 122026 212134
rect 122262 211898 122346 212134
rect 122582 211898 150026 212134
rect 150262 211898 150346 212134
rect 150582 211898 178026 212134
rect 178262 211898 178346 212134
rect 178582 211898 206026 212134
rect 206262 211898 206346 212134
rect 206582 211898 234026 212134
rect 234262 211898 234346 212134
rect 234582 211898 262026 212134
rect 262262 211898 262346 212134
rect 262582 211898 290026 212134
rect 290262 211898 290346 212134
rect 290582 211898 318026 212134
rect 318262 211898 318346 212134
rect 318582 211898 346026 212134
rect 346262 211898 346346 212134
rect 346582 211898 374026 212134
rect 374262 211898 374346 212134
rect 374582 211898 402026 212134
rect 402262 211898 402346 212134
rect 402582 211898 430026 212134
rect 430262 211898 430346 212134
rect 430582 211898 458026 212134
rect 458262 211898 458346 212134
rect 458582 211898 486026 212134
rect 486262 211898 486346 212134
rect 486582 211898 514026 212134
rect 514262 211898 514346 212134
rect 514582 211898 542026 212134
rect 542262 211898 542346 212134
rect 542582 211898 570026 212134
rect 570262 211898 570346 212134
rect 570582 211898 586302 212134
rect 586538 211898 586622 212134
rect 586858 211898 592650 212134
rect -8726 211866 592650 211898
rect -8726 188829 592650 188861
rect -8726 188593 -1974 188829
rect -1738 188593 -1654 188829
rect -1418 188593 41526 188829
rect 41762 188593 41846 188829
rect 42082 188593 69526 188829
rect 69762 188593 69846 188829
rect 70082 188593 97526 188829
rect 97762 188593 97846 188829
rect 98082 188593 125526 188829
rect 125762 188593 125846 188829
rect 126082 188593 153526 188829
rect 153762 188593 153846 188829
rect 154082 188593 181526 188829
rect 181762 188593 181846 188829
rect 182082 188593 209526 188829
rect 209762 188593 209846 188829
rect 210082 188593 237526 188829
rect 237762 188593 237846 188829
rect 238082 188593 265526 188829
rect 265762 188593 265846 188829
rect 266082 188593 293526 188829
rect 293762 188593 293846 188829
rect 294082 188593 321526 188829
rect 321762 188593 321846 188829
rect 322082 188593 349526 188829
rect 349762 188593 349846 188829
rect 350082 188593 377526 188829
rect 377762 188593 377846 188829
rect 378082 188593 405526 188829
rect 405762 188593 405846 188829
rect 406082 188593 433526 188829
rect 433762 188593 433846 188829
rect 434082 188593 461526 188829
rect 461762 188593 461846 188829
rect 462082 188593 489526 188829
rect 489762 188593 489846 188829
rect 490082 188593 517526 188829
rect 517762 188593 517846 188829
rect 518082 188593 545526 188829
rect 545762 188593 545846 188829
rect 546082 188593 573526 188829
rect 573762 188593 573846 188829
rect 574082 188593 585342 188829
rect 585578 188593 585662 188829
rect 585898 188593 592650 188829
rect -8726 188509 592650 188593
rect -8726 188273 -1974 188509
rect -1738 188273 -1654 188509
rect -1418 188273 41526 188509
rect 41762 188273 41846 188509
rect 42082 188273 69526 188509
rect 69762 188273 69846 188509
rect 70082 188273 97526 188509
rect 97762 188273 97846 188509
rect 98082 188273 125526 188509
rect 125762 188273 125846 188509
rect 126082 188273 153526 188509
rect 153762 188273 153846 188509
rect 154082 188273 181526 188509
rect 181762 188273 181846 188509
rect 182082 188273 209526 188509
rect 209762 188273 209846 188509
rect 210082 188273 237526 188509
rect 237762 188273 237846 188509
rect 238082 188273 265526 188509
rect 265762 188273 265846 188509
rect 266082 188273 293526 188509
rect 293762 188273 293846 188509
rect 294082 188273 321526 188509
rect 321762 188273 321846 188509
rect 322082 188273 349526 188509
rect 349762 188273 349846 188509
rect 350082 188273 377526 188509
rect 377762 188273 377846 188509
rect 378082 188273 405526 188509
rect 405762 188273 405846 188509
rect 406082 188273 433526 188509
rect 433762 188273 433846 188509
rect 434082 188273 461526 188509
rect 461762 188273 461846 188509
rect 462082 188273 489526 188509
rect 489762 188273 489846 188509
rect 490082 188273 517526 188509
rect 517762 188273 517846 188509
rect 518082 188273 545526 188509
rect 545762 188273 545846 188509
rect 546082 188273 573526 188509
rect 573762 188273 573846 188509
rect 574082 188273 585342 188509
rect 585578 188273 585662 188509
rect 585898 188273 592650 188509
rect -8726 188241 592650 188273
rect -8726 185454 592650 185486
rect -8726 185218 -2934 185454
rect -2698 185218 -2614 185454
rect -2378 185218 38026 185454
rect 38262 185218 38346 185454
rect 38582 185218 66026 185454
rect 66262 185218 66346 185454
rect 66582 185218 94026 185454
rect 94262 185218 94346 185454
rect 94582 185218 122026 185454
rect 122262 185218 122346 185454
rect 122582 185218 150026 185454
rect 150262 185218 150346 185454
rect 150582 185218 178026 185454
rect 178262 185218 178346 185454
rect 178582 185218 206026 185454
rect 206262 185218 206346 185454
rect 206582 185218 234026 185454
rect 234262 185218 234346 185454
rect 234582 185218 262026 185454
rect 262262 185218 262346 185454
rect 262582 185218 290026 185454
rect 290262 185218 290346 185454
rect 290582 185218 318026 185454
rect 318262 185218 318346 185454
rect 318582 185218 346026 185454
rect 346262 185218 346346 185454
rect 346582 185218 374026 185454
rect 374262 185218 374346 185454
rect 374582 185218 402026 185454
rect 402262 185218 402346 185454
rect 402582 185218 430026 185454
rect 430262 185218 430346 185454
rect 430582 185218 458026 185454
rect 458262 185218 458346 185454
rect 458582 185218 486026 185454
rect 486262 185218 486346 185454
rect 486582 185218 514026 185454
rect 514262 185218 514346 185454
rect 514582 185218 542026 185454
rect 542262 185218 542346 185454
rect 542582 185218 570026 185454
rect 570262 185218 570346 185454
rect 570582 185218 586302 185454
rect 586538 185218 586622 185454
rect 586858 185218 592650 185454
rect -8726 185134 592650 185218
rect -8726 184898 -2934 185134
rect -2698 184898 -2614 185134
rect -2378 184898 38026 185134
rect 38262 184898 38346 185134
rect 38582 184898 66026 185134
rect 66262 184898 66346 185134
rect 66582 184898 94026 185134
rect 94262 184898 94346 185134
rect 94582 184898 122026 185134
rect 122262 184898 122346 185134
rect 122582 184898 150026 185134
rect 150262 184898 150346 185134
rect 150582 184898 178026 185134
rect 178262 184898 178346 185134
rect 178582 184898 206026 185134
rect 206262 184898 206346 185134
rect 206582 184898 234026 185134
rect 234262 184898 234346 185134
rect 234582 184898 262026 185134
rect 262262 184898 262346 185134
rect 262582 184898 290026 185134
rect 290262 184898 290346 185134
rect 290582 184898 318026 185134
rect 318262 184898 318346 185134
rect 318582 184898 346026 185134
rect 346262 184898 346346 185134
rect 346582 184898 374026 185134
rect 374262 184898 374346 185134
rect 374582 184898 402026 185134
rect 402262 184898 402346 185134
rect 402582 184898 430026 185134
rect 430262 184898 430346 185134
rect 430582 184898 458026 185134
rect 458262 184898 458346 185134
rect 458582 184898 486026 185134
rect 486262 184898 486346 185134
rect 486582 184898 514026 185134
rect 514262 184898 514346 185134
rect 514582 184898 542026 185134
rect 542262 184898 542346 185134
rect 542582 184898 570026 185134
rect 570262 184898 570346 185134
rect 570582 184898 586302 185134
rect 586538 184898 586622 185134
rect 586858 184898 592650 185134
rect -8726 184866 592650 184898
rect -8726 161829 592650 161861
rect -8726 161593 -1974 161829
rect -1738 161593 -1654 161829
rect -1418 161593 41526 161829
rect 41762 161593 41846 161829
rect 42082 161593 69526 161829
rect 69762 161593 69846 161829
rect 70082 161593 97526 161829
rect 97762 161593 97846 161829
rect 98082 161593 125526 161829
rect 125762 161593 125846 161829
rect 126082 161593 153526 161829
rect 153762 161593 153846 161829
rect 154082 161593 181526 161829
rect 181762 161593 181846 161829
rect 182082 161593 209526 161829
rect 209762 161593 209846 161829
rect 210082 161593 237526 161829
rect 237762 161593 237846 161829
rect 238082 161593 265526 161829
rect 265762 161593 265846 161829
rect 266082 161593 293526 161829
rect 293762 161593 293846 161829
rect 294082 161593 321526 161829
rect 321762 161593 321846 161829
rect 322082 161593 349526 161829
rect 349762 161593 349846 161829
rect 350082 161593 377526 161829
rect 377762 161593 377846 161829
rect 378082 161593 405526 161829
rect 405762 161593 405846 161829
rect 406082 161593 433526 161829
rect 433762 161593 433846 161829
rect 434082 161593 461526 161829
rect 461762 161593 461846 161829
rect 462082 161593 489526 161829
rect 489762 161593 489846 161829
rect 490082 161593 517526 161829
rect 517762 161593 517846 161829
rect 518082 161593 545526 161829
rect 545762 161593 545846 161829
rect 546082 161593 573526 161829
rect 573762 161593 573846 161829
rect 574082 161593 585342 161829
rect 585578 161593 585662 161829
rect 585898 161593 592650 161829
rect -8726 161509 592650 161593
rect -8726 161273 -1974 161509
rect -1738 161273 -1654 161509
rect -1418 161273 41526 161509
rect 41762 161273 41846 161509
rect 42082 161273 69526 161509
rect 69762 161273 69846 161509
rect 70082 161273 97526 161509
rect 97762 161273 97846 161509
rect 98082 161273 125526 161509
rect 125762 161273 125846 161509
rect 126082 161273 153526 161509
rect 153762 161273 153846 161509
rect 154082 161273 181526 161509
rect 181762 161273 181846 161509
rect 182082 161273 209526 161509
rect 209762 161273 209846 161509
rect 210082 161273 237526 161509
rect 237762 161273 237846 161509
rect 238082 161273 265526 161509
rect 265762 161273 265846 161509
rect 266082 161273 293526 161509
rect 293762 161273 293846 161509
rect 294082 161273 321526 161509
rect 321762 161273 321846 161509
rect 322082 161273 349526 161509
rect 349762 161273 349846 161509
rect 350082 161273 377526 161509
rect 377762 161273 377846 161509
rect 378082 161273 405526 161509
rect 405762 161273 405846 161509
rect 406082 161273 433526 161509
rect 433762 161273 433846 161509
rect 434082 161273 461526 161509
rect 461762 161273 461846 161509
rect 462082 161273 489526 161509
rect 489762 161273 489846 161509
rect 490082 161273 517526 161509
rect 517762 161273 517846 161509
rect 518082 161273 545526 161509
rect 545762 161273 545846 161509
rect 546082 161273 573526 161509
rect 573762 161273 573846 161509
rect 574082 161273 585342 161509
rect 585578 161273 585662 161509
rect 585898 161273 592650 161509
rect -8726 161241 592650 161273
rect -8726 158454 592650 158486
rect -8726 158218 -2934 158454
rect -2698 158218 -2614 158454
rect -2378 158218 38026 158454
rect 38262 158218 38346 158454
rect 38582 158218 66026 158454
rect 66262 158218 66346 158454
rect 66582 158218 94026 158454
rect 94262 158218 94346 158454
rect 94582 158218 122026 158454
rect 122262 158218 122346 158454
rect 122582 158218 150026 158454
rect 150262 158218 150346 158454
rect 150582 158218 178026 158454
rect 178262 158218 178346 158454
rect 178582 158218 206026 158454
rect 206262 158218 206346 158454
rect 206582 158218 234026 158454
rect 234262 158218 234346 158454
rect 234582 158218 262026 158454
rect 262262 158218 262346 158454
rect 262582 158218 290026 158454
rect 290262 158218 290346 158454
rect 290582 158218 318026 158454
rect 318262 158218 318346 158454
rect 318582 158218 346026 158454
rect 346262 158218 346346 158454
rect 346582 158218 374026 158454
rect 374262 158218 374346 158454
rect 374582 158218 402026 158454
rect 402262 158218 402346 158454
rect 402582 158218 430026 158454
rect 430262 158218 430346 158454
rect 430582 158218 458026 158454
rect 458262 158218 458346 158454
rect 458582 158218 486026 158454
rect 486262 158218 486346 158454
rect 486582 158218 514026 158454
rect 514262 158218 514346 158454
rect 514582 158218 542026 158454
rect 542262 158218 542346 158454
rect 542582 158218 570026 158454
rect 570262 158218 570346 158454
rect 570582 158218 586302 158454
rect 586538 158218 586622 158454
rect 586858 158218 592650 158454
rect -8726 158134 592650 158218
rect -8726 157898 -2934 158134
rect -2698 157898 -2614 158134
rect -2378 157898 38026 158134
rect 38262 157898 38346 158134
rect 38582 157898 66026 158134
rect 66262 157898 66346 158134
rect 66582 157898 94026 158134
rect 94262 157898 94346 158134
rect 94582 157898 122026 158134
rect 122262 157898 122346 158134
rect 122582 157898 150026 158134
rect 150262 157898 150346 158134
rect 150582 157898 178026 158134
rect 178262 157898 178346 158134
rect 178582 157898 206026 158134
rect 206262 157898 206346 158134
rect 206582 157898 234026 158134
rect 234262 157898 234346 158134
rect 234582 157898 262026 158134
rect 262262 157898 262346 158134
rect 262582 157898 290026 158134
rect 290262 157898 290346 158134
rect 290582 157898 318026 158134
rect 318262 157898 318346 158134
rect 318582 157898 346026 158134
rect 346262 157898 346346 158134
rect 346582 157898 374026 158134
rect 374262 157898 374346 158134
rect 374582 157898 402026 158134
rect 402262 157898 402346 158134
rect 402582 157898 430026 158134
rect 430262 157898 430346 158134
rect 430582 157898 458026 158134
rect 458262 157898 458346 158134
rect 458582 157898 486026 158134
rect 486262 157898 486346 158134
rect 486582 157898 514026 158134
rect 514262 157898 514346 158134
rect 514582 157898 542026 158134
rect 542262 157898 542346 158134
rect 542582 157898 570026 158134
rect 570262 157898 570346 158134
rect 570582 157898 586302 158134
rect 586538 157898 586622 158134
rect 586858 157898 592650 158134
rect -8726 157866 592650 157898
rect -8726 134829 592650 134861
rect -8726 134593 -1974 134829
rect -1738 134593 -1654 134829
rect -1418 134593 41526 134829
rect 41762 134593 41846 134829
rect 42082 134593 69526 134829
rect 69762 134593 69846 134829
rect 70082 134593 97526 134829
rect 97762 134593 97846 134829
rect 98082 134593 125526 134829
rect 125762 134593 125846 134829
rect 126082 134593 153526 134829
rect 153762 134593 153846 134829
rect 154082 134593 181526 134829
rect 181762 134593 181846 134829
rect 182082 134593 209526 134829
rect 209762 134593 209846 134829
rect 210082 134593 237526 134829
rect 237762 134593 237846 134829
rect 238082 134593 265526 134829
rect 265762 134593 265846 134829
rect 266082 134593 293526 134829
rect 293762 134593 293846 134829
rect 294082 134593 321526 134829
rect 321762 134593 321846 134829
rect 322082 134593 349526 134829
rect 349762 134593 349846 134829
rect 350082 134593 377526 134829
rect 377762 134593 377846 134829
rect 378082 134593 405526 134829
rect 405762 134593 405846 134829
rect 406082 134593 433526 134829
rect 433762 134593 433846 134829
rect 434082 134593 461526 134829
rect 461762 134593 461846 134829
rect 462082 134593 489526 134829
rect 489762 134593 489846 134829
rect 490082 134593 517526 134829
rect 517762 134593 517846 134829
rect 518082 134593 545526 134829
rect 545762 134593 545846 134829
rect 546082 134593 573526 134829
rect 573762 134593 573846 134829
rect 574082 134593 585342 134829
rect 585578 134593 585662 134829
rect 585898 134593 592650 134829
rect -8726 134509 592650 134593
rect -8726 134273 -1974 134509
rect -1738 134273 -1654 134509
rect -1418 134273 41526 134509
rect 41762 134273 41846 134509
rect 42082 134273 69526 134509
rect 69762 134273 69846 134509
rect 70082 134273 97526 134509
rect 97762 134273 97846 134509
rect 98082 134273 125526 134509
rect 125762 134273 125846 134509
rect 126082 134273 153526 134509
rect 153762 134273 153846 134509
rect 154082 134273 181526 134509
rect 181762 134273 181846 134509
rect 182082 134273 209526 134509
rect 209762 134273 209846 134509
rect 210082 134273 237526 134509
rect 237762 134273 237846 134509
rect 238082 134273 265526 134509
rect 265762 134273 265846 134509
rect 266082 134273 293526 134509
rect 293762 134273 293846 134509
rect 294082 134273 321526 134509
rect 321762 134273 321846 134509
rect 322082 134273 349526 134509
rect 349762 134273 349846 134509
rect 350082 134273 377526 134509
rect 377762 134273 377846 134509
rect 378082 134273 405526 134509
rect 405762 134273 405846 134509
rect 406082 134273 433526 134509
rect 433762 134273 433846 134509
rect 434082 134273 461526 134509
rect 461762 134273 461846 134509
rect 462082 134273 489526 134509
rect 489762 134273 489846 134509
rect 490082 134273 517526 134509
rect 517762 134273 517846 134509
rect 518082 134273 545526 134509
rect 545762 134273 545846 134509
rect 546082 134273 573526 134509
rect 573762 134273 573846 134509
rect 574082 134273 585342 134509
rect 585578 134273 585662 134509
rect 585898 134273 592650 134509
rect -8726 134241 592650 134273
rect -8726 131454 592650 131486
rect -8726 131218 -2934 131454
rect -2698 131218 -2614 131454
rect -2378 131218 38026 131454
rect 38262 131218 38346 131454
rect 38582 131218 66026 131454
rect 66262 131218 66346 131454
rect 66582 131218 94026 131454
rect 94262 131218 94346 131454
rect 94582 131218 122026 131454
rect 122262 131218 122346 131454
rect 122582 131218 150026 131454
rect 150262 131218 150346 131454
rect 150582 131218 178026 131454
rect 178262 131218 178346 131454
rect 178582 131218 206026 131454
rect 206262 131218 206346 131454
rect 206582 131218 234026 131454
rect 234262 131218 234346 131454
rect 234582 131218 262026 131454
rect 262262 131218 262346 131454
rect 262582 131218 290026 131454
rect 290262 131218 290346 131454
rect 290582 131218 318026 131454
rect 318262 131218 318346 131454
rect 318582 131218 346026 131454
rect 346262 131218 346346 131454
rect 346582 131218 374026 131454
rect 374262 131218 374346 131454
rect 374582 131218 402026 131454
rect 402262 131218 402346 131454
rect 402582 131218 430026 131454
rect 430262 131218 430346 131454
rect 430582 131218 458026 131454
rect 458262 131218 458346 131454
rect 458582 131218 486026 131454
rect 486262 131218 486346 131454
rect 486582 131218 514026 131454
rect 514262 131218 514346 131454
rect 514582 131218 542026 131454
rect 542262 131218 542346 131454
rect 542582 131218 570026 131454
rect 570262 131218 570346 131454
rect 570582 131218 586302 131454
rect 586538 131218 586622 131454
rect 586858 131218 592650 131454
rect -8726 131134 592650 131218
rect -8726 130898 -2934 131134
rect -2698 130898 -2614 131134
rect -2378 130898 38026 131134
rect 38262 130898 38346 131134
rect 38582 130898 66026 131134
rect 66262 130898 66346 131134
rect 66582 130898 94026 131134
rect 94262 130898 94346 131134
rect 94582 130898 122026 131134
rect 122262 130898 122346 131134
rect 122582 130898 150026 131134
rect 150262 130898 150346 131134
rect 150582 130898 178026 131134
rect 178262 130898 178346 131134
rect 178582 130898 206026 131134
rect 206262 130898 206346 131134
rect 206582 130898 234026 131134
rect 234262 130898 234346 131134
rect 234582 130898 262026 131134
rect 262262 130898 262346 131134
rect 262582 130898 290026 131134
rect 290262 130898 290346 131134
rect 290582 130898 318026 131134
rect 318262 130898 318346 131134
rect 318582 130898 346026 131134
rect 346262 130898 346346 131134
rect 346582 130898 374026 131134
rect 374262 130898 374346 131134
rect 374582 130898 402026 131134
rect 402262 130898 402346 131134
rect 402582 130898 430026 131134
rect 430262 130898 430346 131134
rect 430582 130898 458026 131134
rect 458262 130898 458346 131134
rect 458582 130898 486026 131134
rect 486262 130898 486346 131134
rect 486582 130898 514026 131134
rect 514262 130898 514346 131134
rect 514582 130898 542026 131134
rect 542262 130898 542346 131134
rect 542582 130898 570026 131134
rect 570262 130898 570346 131134
rect 570582 130898 586302 131134
rect 586538 130898 586622 131134
rect 586858 130898 592650 131134
rect -8726 130866 592650 130898
rect -8726 107829 592650 107861
rect -8726 107593 -1974 107829
rect -1738 107593 -1654 107829
rect -1418 107593 41526 107829
rect 41762 107593 41846 107829
rect 42082 107593 69526 107829
rect 69762 107593 69846 107829
rect 70082 107593 97526 107829
rect 97762 107593 97846 107829
rect 98082 107593 125526 107829
rect 125762 107593 125846 107829
rect 126082 107593 153526 107829
rect 153762 107593 153846 107829
rect 154082 107593 181526 107829
rect 181762 107593 181846 107829
rect 182082 107593 209526 107829
rect 209762 107593 209846 107829
rect 210082 107593 237526 107829
rect 237762 107593 237846 107829
rect 238082 107593 265526 107829
rect 265762 107593 265846 107829
rect 266082 107593 293526 107829
rect 293762 107593 293846 107829
rect 294082 107593 321526 107829
rect 321762 107593 321846 107829
rect 322082 107593 349526 107829
rect 349762 107593 349846 107829
rect 350082 107593 377526 107829
rect 377762 107593 377846 107829
rect 378082 107593 405526 107829
rect 405762 107593 405846 107829
rect 406082 107593 433526 107829
rect 433762 107593 433846 107829
rect 434082 107593 461526 107829
rect 461762 107593 461846 107829
rect 462082 107593 489526 107829
rect 489762 107593 489846 107829
rect 490082 107593 517526 107829
rect 517762 107593 517846 107829
rect 518082 107593 545526 107829
rect 545762 107593 545846 107829
rect 546082 107593 573526 107829
rect 573762 107593 573846 107829
rect 574082 107593 585342 107829
rect 585578 107593 585662 107829
rect 585898 107593 592650 107829
rect -8726 107509 592650 107593
rect -8726 107273 -1974 107509
rect -1738 107273 -1654 107509
rect -1418 107273 41526 107509
rect 41762 107273 41846 107509
rect 42082 107273 69526 107509
rect 69762 107273 69846 107509
rect 70082 107273 97526 107509
rect 97762 107273 97846 107509
rect 98082 107273 125526 107509
rect 125762 107273 125846 107509
rect 126082 107273 153526 107509
rect 153762 107273 153846 107509
rect 154082 107273 181526 107509
rect 181762 107273 181846 107509
rect 182082 107273 209526 107509
rect 209762 107273 209846 107509
rect 210082 107273 237526 107509
rect 237762 107273 237846 107509
rect 238082 107273 265526 107509
rect 265762 107273 265846 107509
rect 266082 107273 293526 107509
rect 293762 107273 293846 107509
rect 294082 107273 321526 107509
rect 321762 107273 321846 107509
rect 322082 107273 349526 107509
rect 349762 107273 349846 107509
rect 350082 107273 377526 107509
rect 377762 107273 377846 107509
rect 378082 107273 405526 107509
rect 405762 107273 405846 107509
rect 406082 107273 433526 107509
rect 433762 107273 433846 107509
rect 434082 107273 461526 107509
rect 461762 107273 461846 107509
rect 462082 107273 489526 107509
rect 489762 107273 489846 107509
rect 490082 107273 517526 107509
rect 517762 107273 517846 107509
rect 518082 107273 545526 107509
rect 545762 107273 545846 107509
rect 546082 107273 573526 107509
rect 573762 107273 573846 107509
rect 574082 107273 585342 107509
rect 585578 107273 585662 107509
rect 585898 107273 592650 107509
rect -8726 107241 592650 107273
rect -8726 104454 592650 104486
rect -8726 104218 -2934 104454
rect -2698 104218 -2614 104454
rect -2378 104218 38026 104454
rect 38262 104218 38346 104454
rect 38582 104218 66026 104454
rect 66262 104218 66346 104454
rect 66582 104218 94026 104454
rect 94262 104218 94346 104454
rect 94582 104218 122026 104454
rect 122262 104218 122346 104454
rect 122582 104218 150026 104454
rect 150262 104218 150346 104454
rect 150582 104218 178026 104454
rect 178262 104218 178346 104454
rect 178582 104218 206026 104454
rect 206262 104218 206346 104454
rect 206582 104218 234026 104454
rect 234262 104218 234346 104454
rect 234582 104218 262026 104454
rect 262262 104218 262346 104454
rect 262582 104218 290026 104454
rect 290262 104218 290346 104454
rect 290582 104218 318026 104454
rect 318262 104218 318346 104454
rect 318582 104218 346026 104454
rect 346262 104218 346346 104454
rect 346582 104218 374026 104454
rect 374262 104218 374346 104454
rect 374582 104218 402026 104454
rect 402262 104218 402346 104454
rect 402582 104218 430026 104454
rect 430262 104218 430346 104454
rect 430582 104218 458026 104454
rect 458262 104218 458346 104454
rect 458582 104218 486026 104454
rect 486262 104218 486346 104454
rect 486582 104218 514026 104454
rect 514262 104218 514346 104454
rect 514582 104218 542026 104454
rect 542262 104218 542346 104454
rect 542582 104218 570026 104454
rect 570262 104218 570346 104454
rect 570582 104218 586302 104454
rect 586538 104218 586622 104454
rect 586858 104218 592650 104454
rect -8726 104134 592650 104218
rect -8726 103898 -2934 104134
rect -2698 103898 -2614 104134
rect -2378 103898 38026 104134
rect 38262 103898 38346 104134
rect 38582 103898 66026 104134
rect 66262 103898 66346 104134
rect 66582 103898 94026 104134
rect 94262 103898 94346 104134
rect 94582 103898 122026 104134
rect 122262 103898 122346 104134
rect 122582 103898 150026 104134
rect 150262 103898 150346 104134
rect 150582 103898 178026 104134
rect 178262 103898 178346 104134
rect 178582 103898 206026 104134
rect 206262 103898 206346 104134
rect 206582 103898 234026 104134
rect 234262 103898 234346 104134
rect 234582 103898 262026 104134
rect 262262 103898 262346 104134
rect 262582 103898 290026 104134
rect 290262 103898 290346 104134
rect 290582 103898 318026 104134
rect 318262 103898 318346 104134
rect 318582 103898 346026 104134
rect 346262 103898 346346 104134
rect 346582 103898 374026 104134
rect 374262 103898 374346 104134
rect 374582 103898 402026 104134
rect 402262 103898 402346 104134
rect 402582 103898 430026 104134
rect 430262 103898 430346 104134
rect 430582 103898 458026 104134
rect 458262 103898 458346 104134
rect 458582 103898 486026 104134
rect 486262 103898 486346 104134
rect 486582 103898 514026 104134
rect 514262 103898 514346 104134
rect 514582 103898 542026 104134
rect 542262 103898 542346 104134
rect 542582 103898 570026 104134
rect 570262 103898 570346 104134
rect 570582 103898 586302 104134
rect 586538 103898 586622 104134
rect 586858 103898 592650 104134
rect -8726 103866 592650 103898
rect -8726 80829 592650 80861
rect -8726 80593 -1974 80829
rect -1738 80593 -1654 80829
rect -1418 80593 41526 80829
rect 41762 80593 41846 80829
rect 42082 80593 69526 80829
rect 69762 80593 69846 80829
rect 70082 80593 97526 80829
rect 97762 80593 97846 80829
rect 98082 80593 125526 80829
rect 125762 80593 125846 80829
rect 126082 80593 153526 80829
rect 153762 80593 153846 80829
rect 154082 80593 181526 80829
rect 181762 80593 181846 80829
rect 182082 80593 209526 80829
rect 209762 80593 209846 80829
rect 210082 80593 237526 80829
rect 237762 80593 237846 80829
rect 238082 80593 265526 80829
rect 265762 80593 265846 80829
rect 266082 80593 293526 80829
rect 293762 80593 293846 80829
rect 294082 80593 321526 80829
rect 321762 80593 321846 80829
rect 322082 80593 349526 80829
rect 349762 80593 349846 80829
rect 350082 80593 377526 80829
rect 377762 80593 377846 80829
rect 378082 80593 405526 80829
rect 405762 80593 405846 80829
rect 406082 80593 433526 80829
rect 433762 80593 433846 80829
rect 434082 80593 461526 80829
rect 461762 80593 461846 80829
rect 462082 80593 489526 80829
rect 489762 80593 489846 80829
rect 490082 80593 517526 80829
rect 517762 80593 517846 80829
rect 518082 80593 545526 80829
rect 545762 80593 545846 80829
rect 546082 80593 573526 80829
rect 573762 80593 573846 80829
rect 574082 80593 585342 80829
rect 585578 80593 585662 80829
rect 585898 80593 592650 80829
rect -8726 80509 592650 80593
rect -8726 80273 -1974 80509
rect -1738 80273 -1654 80509
rect -1418 80273 41526 80509
rect 41762 80273 41846 80509
rect 42082 80273 69526 80509
rect 69762 80273 69846 80509
rect 70082 80273 97526 80509
rect 97762 80273 97846 80509
rect 98082 80273 125526 80509
rect 125762 80273 125846 80509
rect 126082 80273 153526 80509
rect 153762 80273 153846 80509
rect 154082 80273 181526 80509
rect 181762 80273 181846 80509
rect 182082 80273 209526 80509
rect 209762 80273 209846 80509
rect 210082 80273 237526 80509
rect 237762 80273 237846 80509
rect 238082 80273 265526 80509
rect 265762 80273 265846 80509
rect 266082 80273 293526 80509
rect 293762 80273 293846 80509
rect 294082 80273 321526 80509
rect 321762 80273 321846 80509
rect 322082 80273 349526 80509
rect 349762 80273 349846 80509
rect 350082 80273 377526 80509
rect 377762 80273 377846 80509
rect 378082 80273 405526 80509
rect 405762 80273 405846 80509
rect 406082 80273 433526 80509
rect 433762 80273 433846 80509
rect 434082 80273 461526 80509
rect 461762 80273 461846 80509
rect 462082 80273 489526 80509
rect 489762 80273 489846 80509
rect 490082 80273 517526 80509
rect 517762 80273 517846 80509
rect 518082 80273 545526 80509
rect 545762 80273 545846 80509
rect 546082 80273 573526 80509
rect 573762 80273 573846 80509
rect 574082 80273 585342 80509
rect 585578 80273 585662 80509
rect 585898 80273 592650 80509
rect -8726 80241 592650 80273
rect -8726 77454 592650 77486
rect -8726 77218 -2934 77454
rect -2698 77218 -2614 77454
rect -2378 77218 38026 77454
rect 38262 77218 38346 77454
rect 38582 77218 66026 77454
rect 66262 77218 66346 77454
rect 66582 77218 94026 77454
rect 94262 77218 94346 77454
rect 94582 77218 122026 77454
rect 122262 77218 122346 77454
rect 122582 77218 150026 77454
rect 150262 77218 150346 77454
rect 150582 77218 178026 77454
rect 178262 77218 178346 77454
rect 178582 77218 206026 77454
rect 206262 77218 206346 77454
rect 206582 77218 234026 77454
rect 234262 77218 234346 77454
rect 234582 77218 262026 77454
rect 262262 77218 262346 77454
rect 262582 77218 290026 77454
rect 290262 77218 290346 77454
rect 290582 77218 318026 77454
rect 318262 77218 318346 77454
rect 318582 77218 346026 77454
rect 346262 77218 346346 77454
rect 346582 77218 374026 77454
rect 374262 77218 374346 77454
rect 374582 77218 402026 77454
rect 402262 77218 402346 77454
rect 402582 77218 430026 77454
rect 430262 77218 430346 77454
rect 430582 77218 458026 77454
rect 458262 77218 458346 77454
rect 458582 77218 486026 77454
rect 486262 77218 486346 77454
rect 486582 77218 514026 77454
rect 514262 77218 514346 77454
rect 514582 77218 542026 77454
rect 542262 77218 542346 77454
rect 542582 77218 570026 77454
rect 570262 77218 570346 77454
rect 570582 77218 586302 77454
rect 586538 77218 586622 77454
rect 586858 77218 592650 77454
rect -8726 77134 592650 77218
rect -8726 76898 -2934 77134
rect -2698 76898 -2614 77134
rect -2378 76898 38026 77134
rect 38262 76898 38346 77134
rect 38582 76898 66026 77134
rect 66262 76898 66346 77134
rect 66582 76898 94026 77134
rect 94262 76898 94346 77134
rect 94582 76898 122026 77134
rect 122262 76898 122346 77134
rect 122582 76898 150026 77134
rect 150262 76898 150346 77134
rect 150582 76898 178026 77134
rect 178262 76898 178346 77134
rect 178582 76898 206026 77134
rect 206262 76898 206346 77134
rect 206582 76898 234026 77134
rect 234262 76898 234346 77134
rect 234582 76898 262026 77134
rect 262262 76898 262346 77134
rect 262582 76898 290026 77134
rect 290262 76898 290346 77134
rect 290582 76898 318026 77134
rect 318262 76898 318346 77134
rect 318582 76898 346026 77134
rect 346262 76898 346346 77134
rect 346582 76898 374026 77134
rect 374262 76898 374346 77134
rect 374582 76898 402026 77134
rect 402262 76898 402346 77134
rect 402582 76898 430026 77134
rect 430262 76898 430346 77134
rect 430582 76898 458026 77134
rect 458262 76898 458346 77134
rect 458582 76898 486026 77134
rect 486262 76898 486346 77134
rect 486582 76898 514026 77134
rect 514262 76898 514346 77134
rect 514582 76898 542026 77134
rect 542262 76898 542346 77134
rect 542582 76898 570026 77134
rect 570262 76898 570346 77134
rect 570582 76898 586302 77134
rect 586538 76898 586622 77134
rect 586858 76898 592650 77134
rect -8726 76866 592650 76898
rect -8726 53829 592650 53861
rect -8726 53593 -1974 53829
rect -1738 53593 -1654 53829
rect -1418 53593 41526 53829
rect 41762 53593 41846 53829
rect 42082 53593 69526 53829
rect 69762 53593 69846 53829
rect 70082 53593 97526 53829
rect 97762 53593 97846 53829
rect 98082 53593 125526 53829
rect 125762 53593 125846 53829
rect 126082 53593 153526 53829
rect 153762 53593 153846 53829
rect 154082 53593 181526 53829
rect 181762 53593 181846 53829
rect 182082 53593 192960 53829
rect 193196 53593 196908 53829
rect 197144 53593 200856 53829
rect 201092 53593 204804 53829
rect 205040 53593 213260 53829
rect 213496 53593 214208 53829
rect 214444 53593 215156 53829
rect 215392 53593 216104 53829
rect 216340 53593 221960 53829
rect 222196 53593 225908 53829
rect 226144 53593 229856 53829
rect 230092 53593 233804 53829
rect 234040 53593 242260 53829
rect 242496 53593 243208 53829
rect 243444 53593 244156 53829
rect 244392 53593 245104 53829
rect 245340 53593 250960 53829
rect 251196 53593 254908 53829
rect 255144 53593 258856 53829
rect 259092 53593 262804 53829
rect 263040 53593 271260 53829
rect 271496 53593 272208 53829
rect 272444 53593 273156 53829
rect 273392 53593 274104 53829
rect 274340 53593 279960 53829
rect 280196 53593 283908 53829
rect 284144 53593 287856 53829
rect 288092 53593 291804 53829
rect 292040 53593 300260 53829
rect 300496 53593 301208 53829
rect 301444 53593 302156 53829
rect 302392 53593 303104 53829
rect 303340 53593 308960 53829
rect 309196 53593 312908 53829
rect 313144 53593 316856 53829
rect 317092 53593 320804 53829
rect 321040 53593 329260 53829
rect 329496 53593 330208 53829
rect 330444 53593 331156 53829
rect 331392 53593 332104 53829
rect 332340 53593 337960 53829
rect 338196 53593 341908 53829
rect 342144 53593 345856 53829
rect 346092 53593 349804 53829
rect 350040 53593 358260 53829
rect 358496 53593 359208 53829
rect 359444 53593 360156 53829
rect 360392 53593 361104 53829
rect 361340 53593 366960 53829
rect 367196 53593 370908 53829
rect 371144 53593 374856 53829
rect 375092 53593 378804 53829
rect 379040 53593 387260 53829
rect 387496 53593 388208 53829
rect 388444 53593 389156 53829
rect 389392 53593 390104 53829
rect 390340 53593 395960 53829
rect 396196 53593 399908 53829
rect 400144 53593 403856 53829
rect 404092 53593 407804 53829
rect 408040 53593 416260 53829
rect 416496 53593 417208 53829
rect 417444 53593 418156 53829
rect 418392 53593 419104 53829
rect 419340 53593 424960 53829
rect 425196 53593 428908 53829
rect 429144 53593 432856 53829
rect 433092 53593 436804 53829
rect 437040 53593 445260 53829
rect 445496 53593 446208 53829
rect 446444 53593 447156 53829
rect 447392 53593 448104 53829
rect 448340 53593 453960 53829
rect 454196 53593 457908 53829
rect 458144 53593 461856 53829
rect 462092 53593 465804 53829
rect 466040 53593 474260 53829
rect 474496 53593 475208 53829
rect 475444 53593 476156 53829
rect 476392 53593 477104 53829
rect 477340 53593 482960 53829
rect 483196 53593 486908 53829
rect 487144 53593 490856 53829
rect 491092 53593 494804 53829
rect 495040 53593 503260 53829
rect 503496 53593 504208 53829
rect 504444 53593 505156 53829
rect 505392 53593 506104 53829
rect 506340 53593 511960 53829
rect 512196 53593 515908 53829
rect 516144 53593 519856 53829
rect 520092 53593 523804 53829
rect 524040 53593 532260 53829
rect 532496 53593 533208 53829
rect 533444 53593 534156 53829
rect 534392 53593 535104 53829
rect 535340 53593 540960 53829
rect 541196 53593 544908 53829
rect 545144 53593 548856 53829
rect 549092 53593 552804 53829
rect 553040 53593 561260 53829
rect 561496 53593 562208 53829
rect 562444 53593 563156 53829
rect 563392 53593 564104 53829
rect 564340 53593 573526 53829
rect 573762 53593 573846 53829
rect 574082 53593 585342 53829
rect 585578 53593 585662 53829
rect 585898 53593 592650 53829
rect -8726 53509 592650 53593
rect -8726 53273 -1974 53509
rect -1738 53273 -1654 53509
rect -1418 53273 41526 53509
rect 41762 53273 41846 53509
rect 42082 53273 69526 53509
rect 69762 53273 69846 53509
rect 70082 53273 97526 53509
rect 97762 53273 97846 53509
rect 98082 53273 125526 53509
rect 125762 53273 125846 53509
rect 126082 53273 153526 53509
rect 153762 53273 153846 53509
rect 154082 53273 181526 53509
rect 181762 53273 181846 53509
rect 182082 53273 192960 53509
rect 193196 53273 196908 53509
rect 197144 53273 200856 53509
rect 201092 53273 204804 53509
rect 205040 53273 213260 53509
rect 213496 53273 214208 53509
rect 214444 53273 215156 53509
rect 215392 53273 216104 53509
rect 216340 53273 221960 53509
rect 222196 53273 225908 53509
rect 226144 53273 229856 53509
rect 230092 53273 233804 53509
rect 234040 53273 242260 53509
rect 242496 53273 243208 53509
rect 243444 53273 244156 53509
rect 244392 53273 245104 53509
rect 245340 53273 250960 53509
rect 251196 53273 254908 53509
rect 255144 53273 258856 53509
rect 259092 53273 262804 53509
rect 263040 53273 271260 53509
rect 271496 53273 272208 53509
rect 272444 53273 273156 53509
rect 273392 53273 274104 53509
rect 274340 53273 279960 53509
rect 280196 53273 283908 53509
rect 284144 53273 287856 53509
rect 288092 53273 291804 53509
rect 292040 53273 300260 53509
rect 300496 53273 301208 53509
rect 301444 53273 302156 53509
rect 302392 53273 303104 53509
rect 303340 53273 308960 53509
rect 309196 53273 312908 53509
rect 313144 53273 316856 53509
rect 317092 53273 320804 53509
rect 321040 53273 329260 53509
rect 329496 53273 330208 53509
rect 330444 53273 331156 53509
rect 331392 53273 332104 53509
rect 332340 53273 337960 53509
rect 338196 53273 341908 53509
rect 342144 53273 345856 53509
rect 346092 53273 349804 53509
rect 350040 53273 358260 53509
rect 358496 53273 359208 53509
rect 359444 53273 360156 53509
rect 360392 53273 361104 53509
rect 361340 53273 366960 53509
rect 367196 53273 370908 53509
rect 371144 53273 374856 53509
rect 375092 53273 378804 53509
rect 379040 53273 387260 53509
rect 387496 53273 388208 53509
rect 388444 53273 389156 53509
rect 389392 53273 390104 53509
rect 390340 53273 395960 53509
rect 396196 53273 399908 53509
rect 400144 53273 403856 53509
rect 404092 53273 407804 53509
rect 408040 53273 416260 53509
rect 416496 53273 417208 53509
rect 417444 53273 418156 53509
rect 418392 53273 419104 53509
rect 419340 53273 424960 53509
rect 425196 53273 428908 53509
rect 429144 53273 432856 53509
rect 433092 53273 436804 53509
rect 437040 53273 445260 53509
rect 445496 53273 446208 53509
rect 446444 53273 447156 53509
rect 447392 53273 448104 53509
rect 448340 53273 453960 53509
rect 454196 53273 457908 53509
rect 458144 53273 461856 53509
rect 462092 53273 465804 53509
rect 466040 53273 474260 53509
rect 474496 53273 475208 53509
rect 475444 53273 476156 53509
rect 476392 53273 477104 53509
rect 477340 53273 482960 53509
rect 483196 53273 486908 53509
rect 487144 53273 490856 53509
rect 491092 53273 494804 53509
rect 495040 53273 503260 53509
rect 503496 53273 504208 53509
rect 504444 53273 505156 53509
rect 505392 53273 506104 53509
rect 506340 53273 511960 53509
rect 512196 53273 515908 53509
rect 516144 53273 519856 53509
rect 520092 53273 523804 53509
rect 524040 53273 532260 53509
rect 532496 53273 533208 53509
rect 533444 53273 534156 53509
rect 534392 53273 535104 53509
rect 535340 53273 540960 53509
rect 541196 53273 544908 53509
rect 545144 53273 548856 53509
rect 549092 53273 552804 53509
rect 553040 53273 561260 53509
rect 561496 53273 562208 53509
rect 562444 53273 563156 53509
rect 563392 53273 564104 53509
rect 564340 53273 573526 53509
rect 573762 53273 573846 53509
rect 574082 53273 585342 53509
rect 585578 53273 585662 53509
rect 585898 53273 592650 53509
rect -8726 53241 592650 53273
rect -8726 50454 592650 50486
rect -8726 50218 -2934 50454
rect -2698 50218 -2614 50454
rect -2378 50218 38026 50454
rect 38262 50218 38346 50454
rect 38582 50218 66026 50454
rect 66262 50218 66346 50454
rect 66582 50218 94026 50454
rect 94262 50218 94346 50454
rect 94582 50218 122026 50454
rect 122262 50218 122346 50454
rect 122582 50218 150026 50454
rect 150262 50218 150346 50454
rect 150582 50218 178026 50454
rect 178262 50218 178346 50454
rect 178582 50218 194934 50454
rect 195170 50218 198882 50454
rect 199118 50218 202830 50454
rect 203066 50218 213734 50454
rect 213970 50218 214682 50454
rect 214918 50218 215630 50454
rect 215866 50218 223934 50454
rect 224170 50218 227882 50454
rect 228118 50218 231830 50454
rect 232066 50218 242734 50454
rect 242970 50218 243682 50454
rect 243918 50218 244630 50454
rect 244866 50218 252934 50454
rect 253170 50218 256882 50454
rect 257118 50218 260830 50454
rect 261066 50218 271734 50454
rect 271970 50218 272682 50454
rect 272918 50218 273630 50454
rect 273866 50218 281934 50454
rect 282170 50218 285882 50454
rect 286118 50218 289830 50454
rect 290066 50218 300734 50454
rect 300970 50218 301682 50454
rect 301918 50218 302630 50454
rect 302866 50218 310934 50454
rect 311170 50218 314882 50454
rect 315118 50218 318830 50454
rect 319066 50218 329734 50454
rect 329970 50218 330682 50454
rect 330918 50218 331630 50454
rect 331866 50218 339934 50454
rect 340170 50218 343882 50454
rect 344118 50218 347830 50454
rect 348066 50218 358734 50454
rect 358970 50218 359682 50454
rect 359918 50218 360630 50454
rect 360866 50218 368934 50454
rect 369170 50218 372882 50454
rect 373118 50218 376830 50454
rect 377066 50218 387734 50454
rect 387970 50218 388682 50454
rect 388918 50218 389630 50454
rect 389866 50218 397934 50454
rect 398170 50218 401882 50454
rect 402118 50218 405830 50454
rect 406066 50218 416734 50454
rect 416970 50218 417682 50454
rect 417918 50218 418630 50454
rect 418866 50218 426934 50454
rect 427170 50218 430882 50454
rect 431118 50218 434830 50454
rect 435066 50218 445734 50454
rect 445970 50218 446682 50454
rect 446918 50218 447630 50454
rect 447866 50218 455934 50454
rect 456170 50218 459882 50454
rect 460118 50218 463830 50454
rect 464066 50218 474734 50454
rect 474970 50218 475682 50454
rect 475918 50218 476630 50454
rect 476866 50218 484934 50454
rect 485170 50218 488882 50454
rect 489118 50218 492830 50454
rect 493066 50218 503734 50454
rect 503970 50218 504682 50454
rect 504918 50218 505630 50454
rect 505866 50218 513934 50454
rect 514170 50218 517882 50454
rect 518118 50218 521830 50454
rect 522066 50218 532734 50454
rect 532970 50218 533682 50454
rect 533918 50218 534630 50454
rect 534866 50218 542934 50454
rect 543170 50218 546882 50454
rect 547118 50218 550830 50454
rect 551066 50218 561734 50454
rect 561970 50218 562682 50454
rect 562918 50218 563630 50454
rect 563866 50218 570026 50454
rect 570262 50218 570346 50454
rect 570582 50218 586302 50454
rect 586538 50218 586622 50454
rect 586858 50218 592650 50454
rect -8726 50134 592650 50218
rect -8726 49898 -2934 50134
rect -2698 49898 -2614 50134
rect -2378 49898 38026 50134
rect 38262 49898 38346 50134
rect 38582 49898 66026 50134
rect 66262 49898 66346 50134
rect 66582 49898 94026 50134
rect 94262 49898 94346 50134
rect 94582 49898 122026 50134
rect 122262 49898 122346 50134
rect 122582 49898 150026 50134
rect 150262 49898 150346 50134
rect 150582 49898 178026 50134
rect 178262 49898 178346 50134
rect 178582 49898 194934 50134
rect 195170 49898 198882 50134
rect 199118 49898 202830 50134
rect 203066 49898 213734 50134
rect 213970 49898 214682 50134
rect 214918 49898 215630 50134
rect 215866 49898 223934 50134
rect 224170 49898 227882 50134
rect 228118 49898 231830 50134
rect 232066 49898 242734 50134
rect 242970 49898 243682 50134
rect 243918 49898 244630 50134
rect 244866 49898 252934 50134
rect 253170 49898 256882 50134
rect 257118 49898 260830 50134
rect 261066 49898 271734 50134
rect 271970 49898 272682 50134
rect 272918 49898 273630 50134
rect 273866 49898 281934 50134
rect 282170 49898 285882 50134
rect 286118 49898 289830 50134
rect 290066 49898 300734 50134
rect 300970 49898 301682 50134
rect 301918 49898 302630 50134
rect 302866 49898 310934 50134
rect 311170 49898 314882 50134
rect 315118 49898 318830 50134
rect 319066 49898 329734 50134
rect 329970 49898 330682 50134
rect 330918 49898 331630 50134
rect 331866 49898 339934 50134
rect 340170 49898 343882 50134
rect 344118 49898 347830 50134
rect 348066 49898 358734 50134
rect 358970 49898 359682 50134
rect 359918 49898 360630 50134
rect 360866 49898 368934 50134
rect 369170 49898 372882 50134
rect 373118 49898 376830 50134
rect 377066 49898 387734 50134
rect 387970 49898 388682 50134
rect 388918 49898 389630 50134
rect 389866 49898 397934 50134
rect 398170 49898 401882 50134
rect 402118 49898 405830 50134
rect 406066 49898 416734 50134
rect 416970 49898 417682 50134
rect 417918 49898 418630 50134
rect 418866 49898 426934 50134
rect 427170 49898 430882 50134
rect 431118 49898 434830 50134
rect 435066 49898 445734 50134
rect 445970 49898 446682 50134
rect 446918 49898 447630 50134
rect 447866 49898 455934 50134
rect 456170 49898 459882 50134
rect 460118 49898 463830 50134
rect 464066 49898 474734 50134
rect 474970 49898 475682 50134
rect 475918 49898 476630 50134
rect 476866 49898 484934 50134
rect 485170 49898 488882 50134
rect 489118 49898 492830 50134
rect 493066 49898 503734 50134
rect 503970 49898 504682 50134
rect 504918 49898 505630 50134
rect 505866 49898 513934 50134
rect 514170 49898 517882 50134
rect 518118 49898 521830 50134
rect 522066 49898 532734 50134
rect 532970 49898 533682 50134
rect 533918 49898 534630 50134
rect 534866 49898 542934 50134
rect 543170 49898 546882 50134
rect 547118 49898 550830 50134
rect 551066 49898 561734 50134
rect 561970 49898 562682 50134
rect 562918 49898 563630 50134
rect 563866 49898 570026 50134
rect 570262 49898 570346 50134
rect 570582 49898 586302 50134
rect 586538 49898 586622 50134
rect 586858 49898 592650 50134
rect -8726 49866 592650 49898
rect -8726 26829 592650 26861
rect -8726 26593 -1974 26829
rect -1738 26593 -1654 26829
rect -1418 26593 22460 26829
rect 22696 26593 33408 26829
rect 33644 26593 44356 26829
rect 44592 26593 55304 26829
rect 55540 26593 69526 26829
rect 69762 26593 69846 26829
rect 70082 26593 75460 26829
rect 75696 26593 76408 26829
rect 76644 26593 77356 26829
rect 77592 26593 78304 26829
rect 78540 26593 84160 26829
rect 84396 26593 88108 26829
rect 88344 26593 92056 26829
rect 92292 26593 96004 26829
rect 96240 26593 104460 26829
rect 104696 26593 105408 26829
rect 105644 26593 106356 26829
rect 106592 26593 107304 26829
rect 107540 26593 113160 26829
rect 113396 26593 117108 26829
rect 117344 26593 121056 26829
rect 121292 26593 125004 26829
rect 125240 26593 133460 26829
rect 133696 26593 134408 26829
rect 134644 26593 135356 26829
rect 135592 26593 136304 26829
rect 136540 26593 142160 26829
rect 142396 26593 146108 26829
rect 146344 26593 150056 26829
rect 150292 26593 154004 26829
rect 154240 26593 162460 26829
rect 162696 26593 163408 26829
rect 163644 26593 164356 26829
rect 164592 26593 165304 26829
rect 165540 26593 171160 26829
rect 171396 26593 175108 26829
rect 175344 26593 179056 26829
rect 179292 26593 183004 26829
rect 183240 26593 191460 26829
rect 191696 26593 192408 26829
rect 192644 26593 193356 26829
rect 193592 26593 194304 26829
rect 194540 26593 200160 26829
rect 200396 26593 204108 26829
rect 204344 26593 208056 26829
rect 208292 26593 212004 26829
rect 212240 26593 220460 26829
rect 220696 26593 221408 26829
rect 221644 26593 222356 26829
rect 222592 26593 223304 26829
rect 223540 26593 229160 26829
rect 229396 26593 233108 26829
rect 233344 26593 237056 26829
rect 237292 26593 241004 26829
rect 241240 26593 249460 26829
rect 249696 26593 250408 26829
rect 250644 26593 251356 26829
rect 251592 26593 252304 26829
rect 252540 26593 258160 26829
rect 258396 26593 262108 26829
rect 262344 26593 266056 26829
rect 266292 26593 270004 26829
rect 270240 26593 278460 26829
rect 278696 26593 279408 26829
rect 279644 26593 280356 26829
rect 280592 26593 281304 26829
rect 281540 26593 287160 26829
rect 287396 26593 291108 26829
rect 291344 26593 295056 26829
rect 295292 26593 299004 26829
rect 299240 26593 307460 26829
rect 307696 26593 308408 26829
rect 308644 26593 309356 26829
rect 309592 26593 310304 26829
rect 310540 26593 316160 26829
rect 316396 26593 320108 26829
rect 320344 26593 324056 26829
rect 324292 26593 328004 26829
rect 328240 26593 336460 26829
rect 336696 26593 337408 26829
rect 337644 26593 338356 26829
rect 338592 26593 339304 26829
rect 339540 26593 345160 26829
rect 345396 26593 349108 26829
rect 349344 26593 353056 26829
rect 353292 26593 357004 26829
rect 357240 26593 365460 26829
rect 365696 26593 366408 26829
rect 366644 26593 367356 26829
rect 367592 26593 368304 26829
rect 368540 26593 374160 26829
rect 374396 26593 378108 26829
rect 378344 26593 382056 26829
rect 382292 26593 386004 26829
rect 386240 26593 394460 26829
rect 394696 26593 395408 26829
rect 395644 26593 396356 26829
rect 396592 26593 397304 26829
rect 397540 26593 403160 26829
rect 403396 26593 407108 26829
rect 407344 26593 411056 26829
rect 411292 26593 415004 26829
rect 415240 26593 423460 26829
rect 423696 26593 424408 26829
rect 424644 26593 425356 26829
rect 425592 26593 426304 26829
rect 426540 26593 432160 26829
rect 432396 26593 436108 26829
rect 436344 26593 440056 26829
rect 440292 26593 444004 26829
rect 444240 26593 452460 26829
rect 452696 26593 453408 26829
rect 453644 26593 454356 26829
rect 454592 26593 455304 26829
rect 455540 26593 461160 26829
rect 461396 26593 465108 26829
rect 465344 26593 469056 26829
rect 469292 26593 473004 26829
rect 473240 26593 481460 26829
rect 481696 26593 482408 26829
rect 482644 26593 483356 26829
rect 483592 26593 484304 26829
rect 484540 26593 490160 26829
rect 490396 26593 494108 26829
rect 494344 26593 498056 26829
rect 498292 26593 502004 26829
rect 502240 26593 510460 26829
rect 510696 26593 511408 26829
rect 511644 26593 512356 26829
rect 512592 26593 513304 26829
rect 513540 26593 519160 26829
rect 519396 26593 523108 26829
rect 523344 26593 527056 26829
rect 527292 26593 531004 26829
rect 531240 26593 539460 26829
rect 539696 26593 540408 26829
rect 540644 26593 541356 26829
rect 541592 26593 542304 26829
rect 542540 26593 548160 26829
rect 548396 26593 552108 26829
rect 552344 26593 556056 26829
rect 556292 26593 560004 26829
rect 560240 26593 573526 26829
rect 573762 26593 573846 26829
rect 574082 26593 585342 26829
rect 585578 26593 585662 26829
rect 585898 26593 592650 26829
rect -8726 26509 592650 26593
rect -8726 26273 -1974 26509
rect -1738 26273 -1654 26509
rect -1418 26273 22460 26509
rect 22696 26273 33408 26509
rect 33644 26273 44356 26509
rect 44592 26273 55304 26509
rect 55540 26273 69526 26509
rect 69762 26273 69846 26509
rect 70082 26273 75460 26509
rect 75696 26273 76408 26509
rect 76644 26273 77356 26509
rect 77592 26273 78304 26509
rect 78540 26273 84160 26509
rect 84396 26273 88108 26509
rect 88344 26273 92056 26509
rect 92292 26273 96004 26509
rect 96240 26273 104460 26509
rect 104696 26273 105408 26509
rect 105644 26273 106356 26509
rect 106592 26273 107304 26509
rect 107540 26273 113160 26509
rect 113396 26273 117108 26509
rect 117344 26273 121056 26509
rect 121292 26273 125004 26509
rect 125240 26273 133460 26509
rect 133696 26273 134408 26509
rect 134644 26273 135356 26509
rect 135592 26273 136304 26509
rect 136540 26273 142160 26509
rect 142396 26273 146108 26509
rect 146344 26273 150056 26509
rect 150292 26273 154004 26509
rect 154240 26273 162460 26509
rect 162696 26273 163408 26509
rect 163644 26273 164356 26509
rect 164592 26273 165304 26509
rect 165540 26273 171160 26509
rect 171396 26273 175108 26509
rect 175344 26273 179056 26509
rect 179292 26273 183004 26509
rect 183240 26273 191460 26509
rect 191696 26273 192408 26509
rect 192644 26273 193356 26509
rect 193592 26273 194304 26509
rect 194540 26273 200160 26509
rect 200396 26273 204108 26509
rect 204344 26273 208056 26509
rect 208292 26273 212004 26509
rect 212240 26273 220460 26509
rect 220696 26273 221408 26509
rect 221644 26273 222356 26509
rect 222592 26273 223304 26509
rect 223540 26273 229160 26509
rect 229396 26273 233108 26509
rect 233344 26273 237056 26509
rect 237292 26273 241004 26509
rect 241240 26273 249460 26509
rect 249696 26273 250408 26509
rect 250644 26273 251356 26509
rect 251592 26273 252304 26509
rect 252540 26273 258160 26509
rect 258396 26273 262108 26509
rect 262344 26273 266056 26509
rect 266292 26273 270004 26509
rect 270240 26273 278460 26509
rect 278696 26273 279408 26509
rect 279644 26273 280356 26509
rect 280592 26273 281304 26509
rect 281540 26273 287160 26509
rect 287396 26273 291108 26509
rect 291344 26273 295056 26509
rect 295292 26273 299004 26509
rect 299240 26273 307460 26509
rect 307696 26273 308408 26509
rect 308644 26273 309356 26509
rect 309592 26273 310304 26509
rect 310540 26273 316160 26509
rect 316396 26273 320108 26509
rect 320344 26273 324056 26509
rect 324292 26273 328004 26509
rect 328240 26273 336460 26509
rect 336696 26273 337408 26509
rect 337644 26273 338356 26509
rect 338592 26273 339304 26509
rect 339540 26273 345160 26509
rect 345396 26273 349108 26509
rect 349344 26273 353056 26509
rect 353292 26273 357004 26509
rect 357240 26273 365460 26509
rect 365696 26273 366408 26509
rect 366644 26273 367356 26509
rect 367592 26273 368304 26509
rect 368540 26273 374160 26509
rect 374396 26273 378108 26509
rect 378344 26273 382056 26509
rect 382292 26273 386004 26509
rect 386240 26273 394460 26509
rect 394696 26273 395408 26509
rect 395644 26273 396356 26509
rect 396592 26273 397304 26509
rect 397540 26273 403160 26509
rect 403396 26273 407108 26509
rect 407344 26273 411056 26509
rect 411292 26273 415004 26509
rect 415240 26273 423460 26509
rect 423696 26273 424408 26509
rect 424644 26273 425356 26509
rect 425592 26273 426304 26509
rect 426540 26273 432160 26509
rect 432396 26273 436108 26509
rect 436344 26273 440056 26509
rect 440292 26273 444004 26509
rect 444240 26273 452460 26509
rect 452696 26273 453408 26509
rect 453644 26273 454356 26509
rect 454592 26273 455304 26509
rect 455540 26273 461160 26509
rect 461396 26273 465108 26509
rect 465344 26273 469056 26509
rect 469292 26273 473004 26509
rect 473240 26273 481460 26509
rect 481696 26273 482408 26509
rect 482644 26273 483356 26509
rect 483592 26273 484304 26509
rect 484540 26273 490160 26509
rect 490396 26273 494108 26509
rect 494344 26273 498056 26509
rect 498292 26273 502004 26509
rect 502240 26273 510460 26509
rect 510696 26273 511408 26509
rect 511644 26273 512356 26509
rect 512592 26273 513304 26509
rect 513540 26273 519160 26509
rect 519396 26273 523108 26509
rect 523344 26273 527056 26509
rect 527292 26273 531004 26509
rect 531240 26273 539460 26509
rect 539696 26273 540408 26509
rect 540644 26273 541356 26509
rect 541592 26273 542304 26509
rect 542540 26273 548160 26509
rect 548396 26273 552108 26509
rect 552344 26273 556056 26509
rect 556292 26273 560004 26509
rect 560240 26273 573526 26509
rect 573762 26273 573846 26509
rect 574082 26273 585342 26509
rect 585578 26273 585662 26509
rect 585898 26273 592650 26509
rect -8726 26241 592650 26273
rect -8726 23454 592650 23486
rect -8726 23218 -2934 23454
rect -2698 23218 -2614 23454
rect -2378 23218 27934 23454
rect 28170 23218 38882 23454
rect 39118 23218 49830 23454
rect 50066 23218 60778 23454
rect 61014 23218 66026 23454
rect 66262 23218 66346 23454
rect 66582 23218 75934 23454
rect 76170 23218 76882 23454
rect 77118 23218 77830 23454
rect 78066 23218 86134 23454
rect 86370 23218 90082 23454
rect 90318 23218 94030 23454
rect 94266 23218 104934 23454
rect 105170 23218 105882 23454
rect 106118 23218 106830 23454
rect 107066 23218 115134 23454
rect 115370 23218 119082 23454
rect 119318 23218 123030 23454
rect 123266 23218 133934 23454
rect 134170 23218 134882 23454
rect 135118 23218 135830 23454
rect 136066 23218 144134 23454
rect 144370 23218 148082 23454
rect 148318 23218 152030 23454
rect 152266 23218 162934 23454
rect 163170 23218 163882 23454
rect 164118 23218 164830 23454
rect 165066 23218 173134 23454
rect 173370 23218 177082 23454
rect 177318 23218 181030 23454
rect 181266 23218 191934 23454
rect 192170 23218 192882 23454
rect 193118 23218 193830 23454
rect 194066 23218 202134 23454
rect 202370 23218 206082 23454
rect 206318 23218 210030 23454
rect 210266 23218 220934 23454
rect 221170 23218 221882 23454
rect 222118 23218 222830 23454
rect 223066 23218 231134 23454
rect 231370 23218 235082 23454
rect 235318 23218 239030 23454
rect 239266 23218 249934 23454
rect 250170 23218 250882 23454
rect 251118 23218 251830 23454
rect 252066 23218 260134 23454
rect 260370 23218 264082 23454
rect 264318 23218 268030 23454
rect 268266 23218 278934 23454
rect 279170 23218 279882 23454
rect 280118 23218 280830 23454
rect 281066 23218 289134 23454
rect 289370 23218 293082 23454
rect 293318 23218 297030 23454
rect 297266 23218 307934 23454
rect 308170 23218 308882 23454
rect 309118 23218 309830 23454
rect 310066 23218 318134 23454
rect 318370 23218 322082 23454
rect 322318 23218 326030 23454
rect 326266 23218 336934 23454
rect 337170 23218 337882 23454
rect 338118 23218 338830 23454
rect 339066 23218 347134 23454
rect 347370 23218 351082 23454
rect 351318 23218 355030 23454
rect 355266 23218 365934 23454
rect 366170 23218 366882 23454
rect 367118 23218 367830 23454
rect 368066 23218 376134 23454
rect 376370 23218 380082 23454
rect 380318 23218 384030 23454
rect 384266 23218 394934 23454
rect 395170 23218 395882 23454
rect 396118 23218 396830 23454
rect 397066 23218 405134 23454
rect 405370 23218 409082 23454
rect 409318 23218 413030 23454
rect 413266 23218 423934 23454
rect 424170 23218 424882 23454
rect 425118 23218 425830 23454
rect 426066 23218 434134 23454
rect 434370 23218 438082 23454
rect 438318 23218 442030 23454
rect 442266 23218 452934 23454
rect 453170 23218 453882 23454
rect 454118 23218 454830 23454
rect 455066 23218 463134 23454
rect 463370 23218 467082 23454
rect 467318 23218 471030 23454
rect 471266 23218 481934 23454
rect 482170 23218 482882 23454
rect 483118 23218 483830 23454
rect 484066 23218 492134 23454
rect 492370 23218 496082 23454
rect 496318 23218 500030 23454
rect 500266 23218 510934 23454
rect 511170 23218 511882 23454
rect 512118 23218 512830 23454
rect 513066 23218 521134 23454
rect 521370 23218 525082 23454
rect 525318 23218 529030 23454
rect 529266 23218 539934 23454
rect 540170 23218 540882 23454
rect 541118 23218 541830 23454
rect 542066 23218 550134 23454
rect 550370 23218 554082 23454
rect 554318 23218 558030 23454
rect 558266 23218 570026 23454
rect 570262 23218 570346 23454
rect 570582 23218 586302 23454
rect 586538 23218 586622 23454
rect 586858 23218 592650 23454
rect -8726 23134 592650 23218
rect -8726 22898 -2934 23134
rect -2698 22898 -2614 23134
rect -2378 22898 27934 23134
rect 28170 22898 38882 23134
rect 39118 22898 49830 23134
rect 50066 22898 60778 23134
rect 61014 22898 66026 23134
rect 66262 22898 66346 23134
rect 66582 22898 75934 23134
rect 76170 22898 76882 23134
rect 77118 22898 77830 23134
rect 78066 22898 86134 23134
rect 86370 22898 90082 23134
rect 90318 22898 94030 23134
rect 94266 22898 104934 23134
rect 105170 22898 105882 23134
rect 106118 22898 106830 23134
rect 107066 22898 115134 23134
rect 115370 22898 119082 23134
rect 119318 22898 123030 23134
rect 123266 22898 133934 23134
rect 134170 22898 134882 23134
rect 135118 22898 135830 23134
rect 136066 22898 144134 23134
rect 144370 22898 148082 23134
rect 148318 22898 152030 23134
rect 152266 22898 162934 23134
rect 163170 22898 163882 23134
rect 164118 22898 164830 23134
rect 165066 22898 173134 23134
rect 173370 22898 177082 23134
rect 177318 22898 181030 23134
rect 181266 22898 191934 23134
rect 192170 22898 192882 23134
rect 193118 22898 193830 23134
rect 194066 22898 202134 23134
rect 202370 22898 206082 23134
rect 206318 22898 210030 23134
rect 210266 22898 220934 23134
rect 221170 22898 221882 23134
rect 222118 22898 222830 23134
rect 223066 22898 231134 23134
rect 231370 22898 235082 23134
rect 235318 22898 239030 23134
rect 239266 22898 249934 23134
rect 250170 22898 250882 23134
rect 251118 22898 251830 23134
rect 252066 22898 260134 23134
rect 260370 22898 264082 23134
rect 264318 22898 268030 23134
rect 268266 22898 278934 23134
rect 279170 22898 279882 23134
rect 280118 22898 280830 23134
rect 281066 22898 289134 23134
rect 289370 22898 293082 23134
rect 293318 22898 297030 23134
rect 297266 22898 307934 23134
rect 308170 22898 308882 23134
rect 309118 22898 309830 23134
rect 310066 22898 318134 23134
rect 318370 22898 322082 23134
rect 322318 22898 326030 23134
rect 326266 22898 336934 23134
rect 337170 22898 337882 23134
rect 338118 22898 338830 23134
rect 339066 22898 347134 23134
rect 347370 22898 351082 23134
rect 351318 22898 355030 23134
rect 355266 22898 365934 23134
rect 366170 22898 366882 23134
rect 367118 22898 367830 23134
rect 368066 22898 376134 23134
rect 376370 22898 380082 23134
rect 380318 22898 384030 23134
rect 384266 22898 394934 23134
rect 395170 22898 395882 23134
rect 396118 22898 396830 23134
rect 397066 22898 405134 23134
rect 405370 22898 409082 23134
rect 409318 22898 413030 23134
rect 413266 22898 423934 23134
rect 424170 22898 424882 23134
rect 425118 22898 425830 23134
rect 426066 22898 434134 23134
rect 434370 22898 438082 23134
rect 438318 22898 442030 23134
rect 442266 22898 452934 23134
rect 453170 22898 453882 23134
rect 454118 22898 454830 23134
rect 455066 22898 463134 23134
rect 463370 22898 467082 23134
rect 467318 22898 471030 23134
rect 471266 22898 481934 23134
rect 482170 22898 482882 23134
rect 483118 22898 483830 23134
rect 484066 22898 492134 23134
rect 492370 22898 496082 23134
rect 496318 22898 500030 23134
rect 500266 22898 510934 23134
rect 511170 22898 511882 23134
rect 512118 22898 512830 23134
rect 513066 22898 521134 23134
rect 521370 22898 525082 23134
rect 525318 22898 529030 23134
rect 529266 22898 539934 23134
rect 540170 22898 540882 23134
rect 541118 22898 541830 23134
rect 542066 22898 550134 23134
rect 550370 22898 554082 23134
rect 554318 22898 558030 23134
rect 558266 22898 570026 23134
rect 570262 22898 570346 23134
rect 570582 22898 586302 23134
rect 586538 22898 586622 23134
rect 586858 22898 592650 23134
rect -8726 22866 592650 22898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 69526 -346
rect 69762 -582 69846 -346
rect 70082 -582 573526 -346
rect 573762 -582 573846 -346
rect 574082 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 69526 -666
rect 69762 -902 69846 -666
rect 70082 -902 573526 -666
rect 573762 -902 573846 -666
rect 574082 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 66026 -1306
rect 66262 -1542 66346 -1306
rect 66582 -1542 570026 -1306
rect 570262 -1542 570346 -1306
rect 570582 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 66026 -1626
rect 66262 -1862 66346 -1626
rect 66582 -1862 570026 -1626
rect 570262 -1862 570346 -1626
rect 570582 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use scan_controller  scan_controller
timestamp 0
transform 1 0 16000 0 1 16000
box -10 0 46000 20000
use scanchain  scanchain_0
timestamp 0
transform 1 0 74000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_1
timestamp 0
transform 1 0 103000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_2
timestamp 0
transform 1 0 132000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_3
timestamp 0
transform 1 0 161000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_4
timestamp 0
transform 1 0 190000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_5
timestamp 0
transform 1 0 219000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_6
timestamp 0
transform 1 0 248000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_7
timestamp 0
transform 1 0 277000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_8
timestamp 0
transform 1 0 306000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_9
timestamp 0
transform 1 0 335000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_10
timestamp 0
transform 1 0 364000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_11
timestamp 0
transform 1 0 393000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_12
timestamp 0
transform 1 0 422000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_13
timestamp 0
transform 1 0 451000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_14
timestamp 0
transform 1 0 480000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_15
timestamp 0
transform 1 0 509000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_16
timestamp 0
transform 1 0 538000 0 1 16000
box 0 688 6000 23248
use scanchain  scanchain_17
timestamp 0
transform -1 0 565800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_18
timestamp 0
transform -1 0 536800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_19
timestamp 0
transform -1 0 507800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_20
timestamp 0
transform -1 0 478800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_21
timestamp 0
transform -1 0 449800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_22
timestamp 0
transform -1 0 420800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_23
timestamp 0
transform -1 0 391800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_24
timestamp 0
transform -1 0 362800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_25
timestamp 0
transform -1 0 333800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_26
timestamp 0
transform -1 0 304800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_27
timestamp 0
transform -1 0 275800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_28
timestamp 0
transform -1 0 246800 0 -1 67000
box 0 688 6000 23248
use scanchain  scanchain_29
timestamp 0
transform -1 0 217800 0 -1 67000
box 0 688 6000 23248
use user_module_341535056611770964  user_module_341535056611770964_0
timestamp 0
transform 1 0 81200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_1
timestamp 0
transform 1 0 110200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_2
timestamp 0
transform 1 0 139200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_3
timestamp 0
transform 1 0 168200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_4
timestamp 0
transform 1 0 197200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_5
timestamp 0
transform 1 0 226200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_6
timestamp 0
transform 1 0 255200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_7
timestamp 0
transform 1 0 284200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_8
timestamp 0
transform 1 0 313200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_9
timestamp 0
transform 1 0 342200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_10
timestamp 0
transform 1 0 371200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_11
timestamp 0
transform 1 0 400200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_12
timestamp 0
transform 1 0 429200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_13
timestamp 0
transform 1 0 458200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_14
timestamp 0
transform 1 0 487200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_15
timestamp 0
transform 1 0 516200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_16
timestamp 0
transform 1 0 545200 0 1 16000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_17
timestamp 0
transform -1 0 556000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_18
timestamp 0
transform -1 0 527000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_19
timestamp 0
transform -1 0 498000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_20
timestamp 0
transform -1 0 469000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_21
timestamp 0
transform -1 0 440000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_22
timestamp 0
transform -1 0 411000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_23
timestamp 0
transform -1 0 382000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_24
timestamp 0
transform -1 0 353000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_25
timestamp 0
transform -1 0 324000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_26
timestamp 0
transform -1 0 295000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_27
timestamp 0
transform -1 0 266000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_28
timestamp 0
transform -1 0 237000 0 -1 67000
box 0 688 16836 23248
use user_module_341535056611770964  user_module_341535056611770964_29
timestamp 0
transform -1 0 208000 0 -1 67000
box 0 688 16836 23248
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 41494 38000 42114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 69494 -7654 70114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 97494 42000 98114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 125494 42000 126114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 153494 42000 154114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181494 42000 182114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 209494 69000 210114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 237494 69000 238114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 265494 69000 266114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 293494 69000 294114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 321494 69000 322114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 349494 69000 350114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 377494 69000 378114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 405494 69000 406114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433494 69000 434114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 461494 69000 462114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 489494 69000 490114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 517494 69000 518114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 545494 69000 546114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 573494 -7654 574114 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 26241 592650 26861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 53241 592650 53861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 80241 592650 80861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 107241 592650 107861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 134241 592650 134861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 161241 592650 161861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 188241 592650 188861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 215241 592650 215861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 242241 592650 242861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 269241 592650 269861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 296241 592650 296861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 323241 592650 323861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 350241 592650 350861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 377241 592650 377861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 404241 592650 404861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 431241 592650 431861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 458241 592650 458861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 485241 592650 485861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 512241 592650 512861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 539241 592650 539861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 566241 592650 566861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 593241 592650 593861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 620241 592650 620861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 647241 592650 647861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 674241 592650 674861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 701241 592650 701861 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 37994 38000 38614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 65994 -7654 66614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 93994 42000 94614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 121994 42000 122614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149994 42000 150614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 177994 42000 178614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 205994 69000 206614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 233994 69000 234614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 261994 69000 262614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 289994 69000 290614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 317994 69000 318614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 345994 69000 346614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 373994 69000 374614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401994 69000 402614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 429994 69000 430614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 457994 69000 458614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 485994 69000 486614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 513994 69000 514614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 541994 69000 542614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 569994 -7654 570614 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 22866 592650 23486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 49866 592650 50486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 76866 592650 77486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 103866 592650 104486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 130866 592650 131486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 157866 592650 158486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 184866 592650 185486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 211866 592650 212486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 238866 592650 239486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 265866 592650 266486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 292866 592650 293486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 319866 592650 320486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 346866 592650 347486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 373866 592650 374486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 400866 592650 401486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 427866 592650 428486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 454866 592650 455486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 481866 592650 482486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 508866 592650 509486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 535866 592650 536486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 562866 592650 563486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 589866 592650 590486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 616866 592650 617486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 643866 592650 644486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 670866 592650 671486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 697866 592650 698486 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
