module gatecat_fpga_top (vccd1,
    vssd1,
    io_in,
    io_out);
 input vccd1;
 input vssd1;
 input [7:0] io_in;
 output [7:0] io_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire cfg_datain;
 wire cfg_frameinc;
 wire cfg_framestrb;
 wire \frame_ctr[0] ;
 wire \frame_ctr[1] ;
 wire \frame_ctr[2] ;
 wire \frame_ctr[3] ;
 wire gated_strobe;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \y_c[0].x_c[0].lc_i.B ;
 wire \y_c[0].x_c[0].lc_i.L ;
 wire \y_c[0].x_c[0].lc_i.Q ;
 wire \y_c[0].x_c[0].lc_i.R ;
 wire \y_c[0].x_c[0].lc_i.T ;
 wire \y_c[0].x_c[0].lc_i.cfg[0] ;
 wire \y_c[0].x_c[0].lc_i.cfg[1] ;
 wire \y_c[0].x_c[0].lc_i.cfg[2] ;
 wire \y_c[0].x_c[0].lc_i.cfg[3] ;
 wire \y_c[0].x_c[0].lc_i.cfg[4] ;
 wire \y_c[0].x_c[0].lc_i.cfg[5] ;
 wire \y_c[0].x_c[0].lc_i.cfg[6] ;
 wire \y_c[0].x_c[0].lc_i.cfg[7] ;
 wire \y_c[0].x_c[0].lc_i.cfg_data[0] ;
 wire \y_c[0].x_c[0].lc_i.cfg_data[1] ;
 wire \y_c[0].x_c[0].lc_i.cfg_data[2] ;
 wire \y_c[0].x_c[0].lc_i.cfg_data[3] ;
 wire \y_c[0].x_c[0].lc_i.cfg_mode ;
 wire \y_c[0].x_c[0].lc_i.cfg_strb[0] ;
 wire \y_c[0].x_c[0].lc_i.cfg_strb[1] ;
 wire \y_c[0].x_c[0].lc_i.dff.dffo_n ;
 wire \y_c[0].x_c[0].lc_i.i0 ;
 wire \y_c[0].x_c[0].lc_i.i0a ;
 wire \y_c[0].x_c[0].lc_i.i0b ;
 wire \y_c[0].x_c[0].lc_i.i1 ;
 wire \y_c[0].x_c[0].lc_i.i1a ;
 wire \y_c[0].x_c[0].lc_i.i1b ;
 wire \y_c[0].x_c[0].lc_i.muxo_n ;
 wire \y_c[0].x_c[0].lc_i.s0 ;
 wire \y_c[0].x_c[0].lc_i.s0a ;
 wire \y_c[0].x_c[0].lc_i.s0b ;
 wire \y_c[0].x_c[0].lc_i.s0s ;
 wire \y_c[0].x_c[1].lc_i.B ;
 wire \y_c[0].x_c[1].lc_i.R ;
 wire \y_c[0].x_c[1].lc_i.cfg[0] ;
 wire \y_c[0].x_c[1].lc_i.cfg[1] ;
 wire \y_c[0].x_c[1].lc_i.cfg[2] ;
 wire \y_c[0].x_c[1].lc_i.cfg[3] ;
 wire \y_c[0].x_c[1].lc_i.cfg[4] ;
 wire \y_c[0].x_c[1].lc_i.cfg[5] ;
 wire \y_c[0].x_c[1].lc_i.cfg[6] ;
 wire \y_c[0].x_c[1].lc_i.cfg[7] ;
 wire \y_c[0].x_c[1].lc_i.cfg_data[0] ;
 wire \y_c[0].x_c[1].lc_i.cfg_data[1] ;
 wire \y_c[0].x_c[1].lc_i.cfg_data[2] ;
 wire \y_c[0].x_c[1].lc_i.cfg_data[3] ;
 wire \y_c[0].x_c[1].lc_i.dff.dffo_n ;
 wire \y_c[0].x_c[1].lc_i.i0 ;
 wire \y_c[0].x_c[1].lc_i.i0a ;
 wire \y_c[0].x_c[1].lc_i.i0b ;
 wire \y_c[0].x_c[1].lc_i.i1 ;
 wire \y_c[0].x_c[1].lc_i.i1a ;
 wire \y_c[0].x_c[1].lc_i.i1b ;
 wire \y_c[0].x_c[1].lc_i.muxo_n ;
 wire \y_c[0].x_c[1].lc_i.s0 ;
 wire \y_c[0].x_c[1].lc_i.s0a ;
 wire \y_c[0].x_c[1].lc_i.s0b ;
 wire \y_c[0].x_c[1].lc_i.s0s ;
 wire \y_c[0].x_c[2].lc_i.B ;
 wire \y_c[0].x_c[2].lc_i.R ;
 wire \y_c[0].x_c[2].lc_i.T ;
 wire \y_c[0].x_c[2].lc_i.cfg[0] ;
 wire \y_c[0].x_c[2].lc_i.cfg[1] ;
 wire \y_c[0].x_c[2].lc_i.cfg[2] ;
 wire \y_c[0].x_c[2].lc_i.cfg[3] ;
 wire \y_c[0].x_c[2].lc_i.cfg[4] ;
 wire \y_c[0].x_c[2].lc_i.cfg[5] ;
 wire \y_c[0].x_c[2].lc_i.cfg[6] ;
 wire \y_c[0].x_c[2].lc_i.cfg[7] ;
 wire \y_c[0].x_c[2].lc_i.cfg_data[0] ;
 wire \y_c[0].x_c[2].lc_i.cfg_data[1] ;
 wire \y_c[0].x_c[2].lc_i.cfg_data[2] ;
 wire \y_c[0].x_c[2].lc_i.cfg_data[3] ;
 wire \y_c[0].x_c[2].lc_i.dff.dffo_n ;
 wire \y_c[0].x_c[2].lc_i.i0 ;
 wire \y_c[0].x_c[2].lc_i.i0a ;
 wire \y_c[0].x_c[2].lc_i.i0b ;
 wire \y_c[0].x_c[2].lc_i.i1 ;
 wire \y_c[0].x_c[2].lc_i.i1a ;
 wire \y_c[0].x_c[2].lc_i.i1b ;
 wire \y_c[0].x_c[2].lc_i.muxo_n ;
 wire \y_c[0].x_c[2].lc_i.s0 ;
 wire \y_c[0].x_c[2].lc_i.s0a ;
 wire \y_c[0].x_c[2].lc_i.s0b ;
 wire \y_c[0].x_c[2].lc_i.s0s ;
 wire \y_c[0].x_c[3].lc_i.B ;
 wire \y_c[0].x_c[3].lc_i.R ;
 wire \y_c[0].x_c[3].lc_i.T ;
 wire \y_c[0].x_c[3].lc_i.cfg[0] ;
 wire \y_c[0].x_c[3].lc_i.cfg[1] ;
 wire \y_c[0].x_c[3].lc_i.cfg[2] ;
 wire \y_c[0].x_c[3].lc_i.cfg[3] ;
 wire \y_c[0].x_c[3].lc_i.cfg[4] ;
 wire \y_c[0].x_c[3].lc_i.cfg[5] ;
 wire \y_c[0].x_c[3].lc_i.cfg[6] ;
 wire \y_c[0].x_c[3].lc_i.cfg[7] ;
 wire \y_c[0].x_c[3].lc_i.cfg_data[0] ;
 wire \y_c[0].x_c[3].lc_i.cfg_data[1] ;
 wire \y_c[0].x_c[3].lc_i.cfg_data[2] ;
 wire \y_c[0].x_c[3].lc_i.cfg_data[3] ;
 wire \y_c[0].x_c[3].lc_i.dff.dffo_n ;
 wire \y_c[0].x_c[3].lc_i.i0 ;
 wire \y_c[0].x_c[3].lc_i.i0a ;
 wire \y_c[0].x_c[3].lc_i.i0b ;
 wire \y_c[0].x_c[3].lc_i.i1 ;
 wire \y_c[0].x_c[3].lc_i.i1a ;
 wire \y_c[0].x_c[3].lc_i.i1b ;
 wire \y_c[0].x_c[3].lc_i.muxo_n ;
 wire \y_c[0].x_c[3].lc_i.s0 ;
 wire \y_c[0].x_c[3].lc_i.s0a ;
 wire \y_c[0].x_c[3].lc_i.s0b ;
 wire \y_c[0].x_c[3].lc_i.s0s ;
 wire \y_c[0].x_c[4].lc_i.B ;
 wire \y_c[0].x_c[4].lc_i.T ;
 wire \y_c[0].x_c[4].lc_i.cfg[0] ;
 wire \y_c[0].x_c[4].lc_i.cfg[1] ;
 wire \y_c[0].x_c[4].lc_i.cfg[2] ;
 wire \y_c[0].x_c[4].lc_i.cfg[3] ;
 wire \y_c[0].x_c[4].lc_i.cfg[4] ;
 wire \y_c[0].x_c[4].lc_i.cfg[5] ;
 wire \y_c[0].x_c[4].lc_i.cfg[6] ;
 wire \y_c[0].x_c[4].lc_i.cfg[7] ;
 wire \y_c[0].x_c[4].lc_i.cfg_data[0] ;
 wire \y_c[0].x_c[4].lc_i.cfg_data[1] ;
 wire \y_c[0].x_c[4].lc_i.cfg_data[2] ;
 wire \y_c[0].x_c[4].lc_i.cfg_data[3] ;
 wire \y_c[0].x_c[4].lc_i.dff.dffo_n ;
 wire \y_c[0].x_c[4].lc_i.i0 ;
 wire \y_c[0].x_c[4].lc_i.i0a ;
 wire \y_c[0].x_c[4].lc_i.i0b ;
 wire \y_c[0].x_c[4].lc_i.i1 ;
 wire \y_c[0].x_c[4].lc_i.i1a ;
 wire \y_c[0].x_c[4].lc_i.i1b ;
 wire \y_c[0].x_c[4].lc_i.muxo_n ;
 wire \y_c[0].x_c[4].lc_i.s0 ;
 wire \y_c[0].x_c[4].lc_i.s0a ;
 wire \y_c[0].x_c[4].lc_i.s0b ;
 wire \y_c[0].x_c[4].lc_i.s0s ;
 wire \y_c[1].x_c[0].lc_i.B ;
 wire \y_c[1].x_c[0].lc_i.cfg[0] ;
 wire \y_c[1].x_c[0].lc_i.cfg[1] ;
 wire \y_c[1].x_c[0].lc_i.cfg[2] ;
 wire \y_c[1].x_c[0].lc_i.cfg[3] ;
 wire \y_c[1].x_c[0].lc_i.cfg[4] ;
 wire \y_c[1].x_c[0].lc_i.cfg[5] ;
 wire \y_c[1].x_c[0].lc_i.cfg[6] ;
 wire \y_c[1].x_c[0].lc_i.cfg[7] ;
 wire \y_c[1].x_c[0].lc_i.cfg_strb[0] ;
 wire \y_c[1].x_c[0].lc_i.cfg_strb[1] ;
 wire \y_c[1].x_c[0].lc_i.dff.dffo_n ;
 wire \y_c[1].x_c[0].lc_i.i0 ;
 wire \y_c[1].x_c[0].lc_i.i0a ;
 wire \y_c[1].x_c[0].lc_i.i0b ;
 wire \y_c[1].x_c[0].lc_i.i1 ;
 wire \y_c[1].x_c[0].lc_i.i1a ;
 wire \y_c[1].x_c[0].lc_i.i1b ;
 wire \y_c[1].x_c[0].lc_i.muxo_n ;
 wire \y_c[1].x_c[0].lc_i.s0 ;
 wire \y_c[1].x_c[0].lc_i.s0a ;
 wire \y_c[1].x_c[0].lc_i.s0b ;
 wire \y_c[1].x_c[0].lc_i.s0s ;
 wire \y_c[1].x_c[1].lc_i.B ;
 wire \y_c[1].x_c[1].lc_i.cfg[0] ;
 wire \y_c[1].x_c[1].lc_i.cfg[1] ;
 wire \y_c[1].x_c[1].lc_i.cfg[2] ;
 wire \y_c[1].x_c[1].lc_i.cfg[3] ;
 wire \y_c[1].x_c[1].lc_i.cfg[4] ;
 wire \y_c[1].x_c[1].lc_i.cfg[5] ;
 wire \y_c[1].x_c[1].lc_i.cfg[6] ;
 wire \y_c[1].x_c[1].lc_i.cfg[7] ;
 wire \y_c[1].x_c[1].lc_i.dff.dffo_n ;
 wire \y_c[1].x_c[1].lc_i.i0 ;
 wire \y_c[1].x_c[1].lc_i.i0a ;
 wire \y_c[1].x_c[1].lc_i.i0b ;
 wire \y_c[1].x_c[1].lc_i.i1 ;
 wire \y_c[1].x_c[1].lc_i.i1a ;
 wire \y_c[1].x_c[1].lc_i.i1b ;
 wire \y_c[1].x_c[1].lc_i.muxo_n ;
 wire \y_c[1].x_c[1].lc_i.s0 ;
 wire \y_c[1].x_c[1].lc_i.s0a ;
 wire \y_c[1].x_c[1].lc_i.s0b ;
 wire \y_c[1].x_c[1].lc_i.s0s ;
 wire \y_c[1].x_c[2].lc_i.B ;
 wire \y_c[1].x_c[2].lc_i.cfg[0] ;
 wire \y_c[1].x_c[2].lc_i.cfg[1] ;
 wire \y_c[1].x_c[2].lc_i.cfg[2] ;
 wire \y_c[1].x_c[2].lc_i.cfg[3] ;
 wire \y_c[1].x_c[2].lc_i.cfg[4] ;
 wire \y_c[1].x_c[2].lc_i.cfg[5] ;
 wire \y_c[1].x_c[2].lc_i.cfg[6] ;
 wire \y_c[1].x_c[2].lc_i.cfg[7] ;
 wire \y_c[1].x_c[2].lc_i.dff.dffo_n ;
 wire \y_c[1].x_c[2].lc_i.i0 ;
 wire \y_c[1].x_c[2].lc_i.i0a ;
 wire \y_c[1].x_c[2].lc_i.i0b ;
 wire \y_c[1].x_c[2].lc_i.i1 ;
 wire \y_c[1].x_c[2].lc_i.i1a ;
 wire \y_c[1].x_c[2].lc_i.i1b ;
 wire \y_c[1].x_c[2].lc_i.muxo_n ;
 wire \y_c[1].x_c[2].lc_i.s0 ;
 wire \y_c[1].x_c[2].lc_i.s0a ;
 wire \y_c[1].x_c[2].lc_i.s0b ;
 wire \y_c[1].x_c[2].lc_i.s0s ;
 wire \y_c[1].x_c[3].lc_i.B ;
 wire \y_c[1].x_c[3].lc_i.cfg[0] ;
 wire \y_c[1].x_c[3].lc_i.cfg[1] ;
 wire \y_c[1].x_c[3].lc_i.cfg[2] ;
 wire \y_c[1].x_c[3].lc_i.cfg[3] ;
 wire \y_c[1].x_c[3].lc_i.cfg[4] ;
 wire \y_c[1].x_c[3].lc_i.cfg[5] ;
 wire \y_c[1].x_c[3].lc_i.cfg[6] ;
 wire \y_c[1].x_c[3].lc_i.cfg[7] ;
 wire \y_c[1].x_c[3].lc_i.dff.dffo_n ;
 wire \y_c[1].x_c[3].lc_i.i0 ;
 wire \y_c[1].x_c[3].lc_i.i0a ;
 wire \y_c[1].x_c[3].lc_i.i0b ;
 wire \y_c[1].x_c[3].lc_i.i1 ;
 wire \y_c[1].x_c[3].lc_i.i1a ;
 wire \y_c[1].x_c[3].lc_i.i1b ;
 wire \y_c[1].x_c[3].lc_i.muxo_n ;
 wire \y_c[1].x_c[3].lc_i.s0 ;
 wire \y_c[1].x_c[3].lc_i.s0a ;
 wire \y_c[1].x_c[3].lc_i.s0b ;
 wire \y_c[1].x_c[3].lc_i.s0s ;
 wire \y_c[1].x_c[4].lc_i.B ;
 wire \y_c[1].x_c[4].lc_i.cfg[0] ;
 wire \y_c[1].x_c[4].lc_i.cfg[1] ;
 wire \y_c[1].x_c[4].lc_i.cfg[2] ;
 wire \y_c[1].x_c[4].lc_i.cfg[3] ;
 wire \y_c[1].x_c[4].lc_i.cfg[4] ;
 wire \y_c[1].x_c[4].lc_i.cfg[5] ;
 wire \y_c[1].x_c[4].lc_i.cfg[6] ;
 wire \y_c[1].x_c[4].lc_i.cfg[7] ;
 wire \y_c[1].x_c[4].lc_i.dff.dffo_n ;
 wire \y_c[1].x_c[4].lc_i.i0 ;
 wire \y_c[1].x_c[4].lc_i.i0a ;
 wire \y_c[1].x_c[4].lc_i.i0b ;
 wire \y_c[1].x_c[4].lc_i.i1 ;
 wire \y_c[1].x_c[4].lc_i.i1a ;
 wire \y_c[1].x_c[4].lc_i.i1b ;
 wire \y_c[1].x_c[4].lc_i.muxo_n ;
 wire \y_c[1].x_c[4].lc_i.s0 ;
 wire \y_c[1].x_c[4].lc_i.s0a ;
 wire \y_c[1].x_c[4].lc_i.s0b ;
 wire \y_c[1].x_c[4].lc_i.s0s ;
 wire \y_c[2].x_c[0].lc_i.B ;
 wire \y_c[2].x_c[0].lc_i.cfg[0] ;
 wire \y_c[2].x_c[0].lc_i.cfg[1] ;
 wire \y_c[2].x_c[0].lc_i.cfg[2] ;
 wire \y_c[2].x_c[0].lc_i.cfg[3] ;
 wire \y_c[2].x_c[0].lc_i.cfg[4] ;
 wire \y_c[2].x_c[0].lc_i.cfg[5] ;
 wire \y_c[2].x_c[0].lc_i.cfg[6] ;
 wire \y_c[2].x_c[0].lc_i.cfg[7] ;
 wire \y_c[2].x_c[0].lc_i.cfg_strb[0] ;
 wire \y_c[2].x_c[0].lc_i.cfg_strb[1] ;
 wire \y_c[2].x_c[0].lc_i.dff.dffo_n ;
 wire \y_c[2].x_c[0].lc_i.i0 ;
 wire \y_c[2].x_c[0].lc_i.i0a ;
 wire \y_c[2].x_c[0].lc_i.i0b ;
 wire \y_c[2].x_c[0].lc_i.i1 ;
 wire \y_c[2].x_c[0].lc_i.i1a ;
 wire \y_c[2].x_c[0].lc_i.i1b ;
 wire \y_c[2].x_c[0].lc_i.muxo_n ;
 wire \y_c[2].x_c[0].lc_i.s0 ;
 wire \y_c[2].x_c[0].lc_i.s0a ;
 wire \y_c[2].x_c[0].lc_i.s0b ;
 wire \y_c[2].x_c[0].lc_i.s0s ;
 wire \y_c[2].x_c[1].lc_i.B ;
 wire \y_c[2].x_c[1].lc_i.cfg[0] ;
 wire \y_c[2].x_c[1].lc_i.cfg[1] ;
 wire \y_c[2].x_c[1].lc_i.cfg[2] ;
 wire \y_c[2].x_c[1].lc_i.cfg[3] ;
 wire \y_c[2].x_c[1].lc_i.cfg[4] ;
 wire \y_c[2].x_c[1].lc_i.cfg[5] ;
 wire \y_c[2].x_c[1].lc_i.cfg[6] ;
 wire \y_c[2].x_c[1].lc_i.cfg[7] ;
 wire \y_c[2].x_c[1].lc_i.dff.dffo_n ;
 wire \y_c[2].x_c[1].lc_i.i0 ;
 wire \y_c[2].x_c[1].lc_i.i0a ;
 wire \y_c[2].x_c[1].lc_i.i0b ;
 wire \y_c[2].x_c[1].lc_i.i1 ;
 wire \y_c[2].x_c[1].lc_i.i1a ;
 wire \y_c[2].x_c[1].lc_i.i1b ;
 wire \y_c[2].x_c[1].lc_i.muxo_n ;
 wire \y_c[2].x_c[1].lc_i.s0 ;
 wire \y_c[2].x_c[1].lc_i.s0a ;
 wire \y_c[2].x_c[1].lc_i.s0b ;
 wire \y_c[2].x_c[1].lc_i.s0s ;
 wire \y_c[2].x_c[2].lc_i.B ;
 wire \y_c[2].x_c[2].lc_i.cfg[0] ;
 wire \y_c[2].x_c[2].lc_i.cfg[1] ;
 wire \y_c[2].x_c[2].lc_i.cfg[2] ;
 wire \y_c[2].x_c[2].lc_i.cfg[3] ;
 wire \y_c[2].x_c[2].lc_i.cfg[4] ;
 wire \y_c[2].x_c[2].lc_i.cfg[5] ;
 wire \y_c[2].x_c[2].lc_i.cfg[6] ;
 wire \y_c[2].x_c[2].lc_i.cfg[7] ;
 wire \y_c[2].x_c[2].lc_i.dff.dffo_n ;
 wire \y_c[2].x_c[2].lc_i.i0 ;
 wire \y_c[2].x_c[2].lc_i.i0a ;
 wire \y_c[2].x_c[2].lc_i.i0b ;
 wire \y_c[2].x_c[2].lc_i.i1 ;
 wire \y_c[2].x_c[2].lc_i.i1a ;
 wire \y_c[2].x_c[2].lc_i.i1b ;
 wire \y_c[2].x_c[2].lc_i.muxo_n ;
 wire \y_c[2].x_c[2].lc_i.s0 ;
 wire \y_c[2].x_c[2].lc_i.s0a ;
 wire \y_c[2].x_c[2].lc_i.s0b ;
 wire \y_c[2].x_c[2].lc_i.s0s ;
 wire \y_c[2].x_c[3].lc_i.B ;
 wire \y_c[2].x_c[3].lc_i.cfg[0] ;
 wire \y_c[2].x_c[3].lc_i.cfg[1] ;
 wire \y_c[2].x_c[3].lc_i.cfg[2] ;
 wire \y_c[2].x_c[3].lc_i.cfg[3] ;
 wire \y_c[2].x_c[3].lc_i.cfg[4] ;
 wire \y_c[2].x_c[3].lc_i.cfg[5] ;
 wire \y_c[2].x_c[3].lc_i.cfg[6] ;
 wire \y_c[2].x_c[3].lc_i.cfg[7] ;
 wire \y_c[2].x_c[3].lc_i.dff.dffo_n ;
 wire \y_c[2].x_c[3].lc_i.i0 ;
 wire \y_c[2].x_c[3].lc_i.i0a ;
 wire \y_c[2].x_c[3].lc_i.i0b ;
 wire \y_c[2].x_c[3].lc_i.i1 ;
 wire \y_c[2].x_c[3].lc_i.i1a ;
 wire \y_c[2].x_c[3].lc_i.i1b ;
 wire \y_c[2].x_c[3].lc_i.muxo_n ;
 wire \y_c[2].x_c[3].lc_i.s0 ;
 wire \y_c[2].x_c[3].lc_i.s0a ;
 wire \y_c[2].x_c[3].lc_i.s0b ;
 wire \y_c[2].x_c[3].lc_i.s0s ;
 wire \y_c[2].x_c[4].lc_i.B ;
 wire \y_c[2].x_c[4].lc_i.cfg[0] ;
 wire \y_c[2].x_c[4].lc_i.cfg[1] ;
 wire \y_c[2].x_c[4].lc_i.cfg[2] ;
 wire \y_c[2].x_c[4].lc_i.cfg[3] ;
 wire \y_c[2].x_c[4].lc_i.cfg[4] ;
 wire \y_c[2].x_c[4].lc_i.cfg[5] ;
 wire \y_c[2].x_c[4].lc_i.cfg[6] ;
 wire \y_c[2].x_c[4].lc_i.cfg[7] ;
 wire \y_c[2].x_c[4].lc_i.dff.dffo_n ;
 wire \y_c[2].x_c[4].lc_i.i0 ;
 wire \y_c[2].x_c[4].lc_i.i0a ;
 wire \y_c[2].x_c[4].lc_i.i0b ;
 wire \y_c[2].x_c[4].lc_i.i1 ;
 wire \y_c[2].x_c[4].lc_i.i1a ;
 wire \y_c[2].x_c[4].lc_i.i1b ;
 wire \y_c[2].x_c[4].lc_i.muxo_n ;
 wire \y_c[2].x_c[4].lc_i.s0 ;
 wire \y_c[2].x_c[4].lc_i.s0a ;
 wire \y_c[2].x_c[4].lc_i.s0b ;
 wire \y_c[2].x_c[4].lc_i.s0s ;
 wire \y_c[3].x_c[0].lc_i.B ;
 wire \y_c[3].x_c[0].lc_i.cfg[0] ;
 wire \y_c[3].x_c[0].lc_i.cfg[1] ;
 wire \y_c[3].x_c[0].lc_i.cfg[2] ;
 wire \y_c[3].x_c[0].lc_i.cfg[3] ;
 wire \y_c[3].x_c[0].lc_i.cfg[4] ;
 wire \y_c[3].x_c[0].lc_i.cfg[5] ;
 wire \y_c[3].x_c[0].lc_i.cfg[6] ;
 wire \y_c[3].x_c[0].lc_i.cfg[7] ;
 wire \y_c[3].x_c[0].lc_i.cfg_strb[0] ;
 wire \y_c[3].x_c[0].lc_i.cfg_strb[1] ;
 wire \y_c[3].x_c[0].lc_i.dff.dffo_n ;
 wire \y_c[3].x_c[0].lc_i.i0 ;
 wire \y_c[3].x_c[0].lc_i.i0a ;
 wire \y_c[3].x_c[0].lc_i.i0b ;
 wire \y_c[3].x_c[0].lc_i.i1 ;
 wire \y_c[3].x_c[0].lc_i.i1a ;
 wire \y_c[3].x_c[0].lc_i.i1b ;
 wire \y_c[3].x_c[0].lc_i.muxo_n ;
 wire \y_c[3].x_c[0].lc_i.s0 ;
 wire \y_c[3].x_c[0].lc_i.s0a ;
 wire \y_c[3].x_c[0].lc_i.s0b ;
 wire \y_c[3].x_c[0].lc_i.s0s ;
 wire \y_c[3].x_c[1].lc_i.B ;
 wire \y_c[3].x_c[1].lc_i.cfg[0] ;
 wire \y_c[3].x_c[1].lc_i.cfg[1] ;
 wire \y_c[3].x_c[1].lc_i.cfg[2] ;
 wire \y_c[3].x_c[1].lc_i.cfg[3] ;
 wire \y_c[3].x_c[1].lc_i.cfg[4] ;
 wire \y_c[3].x_c[1].lc_i.cfg[5] ;
 wire \y_c[3].x_c[1].lc_i.cfg[6] ;
 wire \y_c[3].x_c[1].lc_i.cfg[7] ;
 wire \y_c[3].x_c[1].lc_i.dff.dffo_n ;
 wire \y_c[3].x_c[1].lc_i.i0 ;
 wire \y_c[3].x_c[1].lc_i.i0a ;
 wire \y_c[3].x_c[1].lc_i.i0b ;
 wire \y_c[3].x_c[1].lc_i.i1 ;
 wire \y_c[3].x_c[1].lc_i.i1a ;
 wire \y_c[3].x_c[1].lc_i.i1b ;
 wire \y_c[3].x_c[1].lc_i.muxo_n ;
 wire \y_c[3].x_c[1].lc_i.s0 ;
 wire \y_c[3].x_c[1].lc_i.s0a ;
 wire \y_c[3].x_c[1].lc_i.s0b ;
 wire \y_c[3].x_c[1].lc_i.s0s ;
 wire \y_c[3].x_c[2].lc_i.B ;
 wire \y_c[3].x_c[2].lc_i.cfg[0] ;
 wire \y_c[3].x_c[2].lc_i.cfg[1] ;
 wire \y_c[3].x_c[2].lc_i.cfg[2] ;
 wire \y_c[3].x_c[2].lc_i.cfg[3] ;
 wire \y_c[3].x_c[2].lc_i.cfg[4] ;
 wire \y_c[3].x_c[2].lc_i.cfg[5] ;
 wire \y_c[3].x_c[2].lc_i.cfg[6] ;
 wire \y_c[3].x_c[2].lc_i.cfg[7] ;
 wire \y_c[3].x_c[2].lc_i.dff.dffo_n ;
 wire \y_c[3].x_c[2].lc_i.i0 ;
 wire \y_c[3].x_c[2].lc_i.i0a ;
 wire \y_c[3].x_c[2].lc_i.i0b ;
 wire \y_c[3].x_c[2].lc_i.i1 ;
 wire \y_c[3].x_c[2].lc_i.i1a ;
 wire \y_c[3].x_c[2].lc_i.i1b ;
 wire \y_c[3].x_c[2].lc_i.muxo_n ;
 wire \y_c[3].x_c[2].lc_i.s0 ;
 wire \y_c[3].x_c[2].lc_i.s0a ;
 wire \y_c[3].x_c[2].lc_i.s0b ;
 wire \y_c[3].x_c[2].lc_i.s0s ;
 wire \y_c[3].x_c[3].lc_i.B ;
 wire \y_c[3].x_c[3].lc_i.cfg[0] ;
 wire \y_c[3].x_c[3].lc_i.cfg[1] ;
 wire \y_c[3].x_c[3].lc_i.cfg[2] ;
 wire \y_c[3].x_c[3].lc_i.cfg[3] ;
 wire \y_c[3].x_c[3].lc_i.cfg[4] ;
 wire \y_c[3].x_c[3].lc_i.cfg[5] ;
 wire \y_c[3].x_c[3].lc_i.cfg[6] ;
 wire \y_c[3].x_c[3].lc_i.cfg[7] ;
 wire \y_c[3].x_c[3].lc_i.dff.dffo_n ;
 wire \y_c[3].x_c[3].lc_i.i0 ;
 wire \y_c[3].x_c[3].lc_i.i0a ;
 wire \y_c[3].x_c[3].lc_i.i0b ;
 wire \y_c[3].x_c[3].lc_i.i1 ;
 wire \y_c[3].x_c[3].lc_i.i1a ;
 wire \y_c[3].x_c[3].lc_i.i1b ;
 wire \y_c[3].x_c[3].lc_i.muxo_n ;
 wire \y_c[3].x_c[3].lc_i.s0 ;
 wire \y_c[3].x_c[3].lc_i.s0a ;
 wire \y_c[3].x_c[3].lc_i.s0b ;
 wire \y_c[3].x_c[3].lc_i.s0s ;
 wire \y_c[3].x_c[4].lc_i.B ;
 wire \y_c[3].x_c[4].lc_i.cfg[0] ;
 wire \y_c[3].x_c[4].lc_i.cfg[1] ;
 wire \y_c[3].x_c[4].lc_i.cfg[2] ;
 wire \y_c[3].x_c[4].lc_i.cfg[3] ;
 wire \y_c[3].x_c[4].lc_i.cfg[4] ;
 wire \y_c[3].x_c[4].lc_i.cfg[5] ;
 wire \y_c[3].x_c[4].lc_i.cfg[6] ;
 wire \y_c[3].x_c[4].lc_i.cfg[7] ;
 wire \y_c[3].x_c[4].lc_i.dff.dffo_n ;
 wire \y_c[3].x_c[4].lc_i.i0 ;
 wire \y_c[3].x_c[4].lc_i.i0a ;
 wire \y_c[3].x_c[4].lc_i.i0b ;
 wire \y_c[3].x_c[4].lc_i.i1 ;
 wire \y_c[3].x_c[4].lc_i.i1a ;
 wire \y_c[3].x_c[4].lc_i.i1b ;
 wire \y_c[3].x_c[4].lc_i.muxo_n ;
 wire \y_c[3].x_c[4].lc_i.s0 ;
 wire \y_c[3].x_c[4].lc_i.s0a ;
 wire \y_c[3].x_c[4].lc_i.s0b ;
 wire \y_c[3].x_c[4].lc_i.s0s ;
 wire \y_c[4].x_c[0].lc_i.B ;
 wire \y_c[4].x_c[0].lc_i.L ;
 wire \y_c[4].x_c[0].lc_i.cfg[0] ;
 wire \y_c[4].x_c[0].lc_i.cfg[1] ;
 wire \y_c[4].x_c[0].lc_i.cfg[2] ;
 wire \y_c[4].x_c[0].lc_i.cfg[3] ;
 wire \y_c[4].x_c[0].lc_i.cfg[4] ;
 wire \y_c[4].x_c[0].lc_i.cfg[5] ;
 wire \y_c[4].x_c[0].lc_i.cfg[6] ;
 wire \y_c[4].x_c[0].lc_i.cfg[7] ;
 wire \y_c[4].x_c[0].lc_i.cfg_strb[0] ;
 wire \y_c[4].x_c[0].lc_i.cfg_strb[1] ;
 wire \y_c[4].x_c[0].lc_i.dff.dffo_n ;
 wire \y_c[4].x_c[0].lc_i.i0 ;
 wire \y_c[4].x_c[0].lc_i.i0a ;
 wire \y_c[4].x_c[0].lc_i.i0b ;
 wire \y_c[4].x_c[0].lc_i.i1 ;
 wire \y_c[4].x_c[0].lc_i.i1a ;
 wire \y_c[4].x_c[0].lc_i.i1b ;
 wire \y_c[4].x_c[0].lc_i.muxo_n ;
 wire \y_c[4].x_c[0].lc_i.s0 ;
 wire \y_c[4].x_c[0].lc_i.s0a ;
 wire \y_c[4].x_c[0].lc_i.s0b ;
 wire \y_c[4].x_c[0].lc_i.s0s ;
 wire \y_c[4].x_c[1].lc_i.B ;
 wire \y_c[4].x_c[1].lc_i.cfg[0] ;
 wire \y_c[4].x_c[1].lc_i.cfg[1] ;
 wire \y_c[4].x_c[1].lc_i.cfg[2] ;
 wire \y_c[4].x_c[1].lc_i.cfg[3] ;
 wire \y_c[4].x_c[1].lc_i.cfg[4] ;
 wire \y_c[4].x_c[1].lc_i.cfg[5] ;
 wire \y_c[4].x_c[1].lc_i.cfg[6] ;
 wire \y_c[4].x_c[1].lc_i.cfg[7] ;
 wire \y_c[4].x_c[1].lc_i.dff.dffo_n ;
 wire \y_c[4].x_c[1].lc_i.i0 ;
 wire \y_c[4].x_c[1].lc_i.i0a ;
 wire \y_c[4].x_c[1].lc_i.i0b ;
 wire \y_c[4].x_c[1].lc_i.i1 ;
 wire \y_c[4].x_c[1].lc_i.i1a ;
 wire \y_c[4].x_c[1].lc_i.i1b ;
 wire \y_c[4].x_c[1].lc_i.muxo_n ;
 wire \y_c[4].x_c[1].lc_i.s0 ;
 wire \y_c[4].x_c[1].lc_i.s0a ;
 wire \y_c[4].x_c[1].lc_i.s0b ;
 wire \y_c[4].x_c[1].lc_i.s0s ;
 wire \y_c[4].x_c[2].lc_i.B ;
 wire \y_c[4].x_c[2].lc_i.cfg[0] ;
 wire \y_c[4].x_c[2].lc_i.cfg[1] ;
 wire \y_c[4].x_c[2].lc_i.cfg[2] ;
 wire \y_c[4].x_c[2].lc_i.cfg[3] ;
 wire \y_c[4].x_c[2].lc_i.cfg[4] ;
 wire \y_c[4].x_c[2].lc_i.cfg[5] ;
 wire \y_c[4].x_c[2].lc_i.cfg[6] ;
 wire \y_c[4].x_c[2].lc_i.cfg[7] ;
 wire \y_c[4].x_c[2].lc_i.dff.dffo_n ;
 wire \y_c[4].x_c[2].lc_i.i0 ;
 wire \y_c[4].x_c[2].lc_i.i0a ;
 wire \y_c[4].x_c[2].lc_i.i0b ;
 wire \y_c[4].x_c[2].lc_i.i1 ;
 wire \y_c[4].x_c[2].lc_i.i1a ;
 wire \y_c[4].x_c[2].lc_i.i1b ;
 wire \y_c[4].x_c[2].lc_i.muxo_n ;
 wire \y_c[4].x_c[2].lc_i.s0 ;
 wire \y_c[4].x_c[2].lc_i.s0a ;
 wire \y_c[4].x_c[2].lc_i.s0b ;
 wire \y_c[4].x_c[2].lc_i.s0s ;
 wire \y_c[4].x_c[3].lc_i.B ;
 wire \y_c[4].x_c[3].lc_i.cfg[0] ;
 wire \y_c[4].x_c[3].lc_i.cfg[1] ;
 wire \y_c[4].x_c[3].lc_i.cfg[2] ;
 wire \y_c[4].x_c[3].lc_i.cfg[3] ;
 wire \y_c[4].x_c[3].lc_i.cfg[4] ;
 wire \y_c[4].x_c[3].lc_i.cfg[5] ;
 wire \y_c[4].x_c[3].lc_i.cfg[6] ;
 wire \y_c[4].x_c[3].lc_i.cfg[7] ;
 wire \y_c[4].x_c[3].lc_i.dff.dffo_n ;
 wire \y_c[4].x_c[3].lc_i.i0 ;
 wire \y_c[4].x_c[3].lc_i.i0a ;
 wire \y_c[4].x_c[3].lc_i.i0b ;
 wire \y_c[4].x_c[3].lc_i.i1 ;
 wire \y_c[4].x_c[3].lc_i.i1a ;
 wire \y_c[4].x_c[3].lc_i.i1b ;
 wire \y_c[4].x_c[3].lc_i.muxo_n ;
 wire \y_c[4].x_c[3].lc_i.s0 ;
 wire \y_c[4].x_c[3].lc_i.s0a ;
 wire \y_c[4].x_c[3].lc_i.s0b ;
 wire \y_c[4].x_c[3].lc_i.s0s ;
 wire \y_c[4].x_c[4].lc_i.B ;
 wire \y_c[4].x_c[4].lc_i.cfg[0] ;
 wire \y_c[4].x_c[4].lc_i.cfg[1] ;
 wire \y_c[4].x_c[4].lc_i.cfg[2] ;
 wire \y_c[4].x_c[4].lc_i.cfg[3] ;
 wire \y_c[4].x_c[4].lc_i.cfg[4] ;
 wire \y_c[4].x_c[4].lc_i.cfg[5] ;
 wire \y_c[4].x_c[4].lc_i.cfg[6] ;
 wire \y_c[4].x_c[4].lc_i.cfg[7] ;
 wire \y_c[4].x_c[4].lc_i.dff.dffo_n ;
 wire \y_c[4].x_c[4].lc_i.i0 ;
 wire \y_c[4].x_c[4].lc_i.i0a ;
 wire \y_c[4].x_c[4].lc_i.i0b ;
 wire \y_c[4].x_c[4].lc_i.i1 ;
 wire \y_c[4].x_c[4].lc_i.i1a ;
 wire \y_c[4].x_c[4].lc_i.i1b ;
 wire \y_c[4].x_c[4].lc_i.muxo_n ;
 wire \y_c[4].x_c[4].lc_i.s0 ;
 wire \y_c[4].x_c[4].lc_i.s0a ;
 wire \y_c[4].x_c[4].lc_i.s0b ;
 wire \y_c[4].x_c[4].lc_i.s0s ;
 wire \y_c[5].x_c[0].lc_i.L ;
 wire \y_c[5].x_c[0].lc_i.cfg[0] ;
 wire \y_c[5].x_c[0].lc_i.cfg[1] ;
 wire \y_c[5].x_c[0].lc_i.cfg[2] ;
 wire \y_c[5].x_c[0].lc_i.cfg[3] ;
 wire \y_c[5].x_c[0].lc_i.cfg[4] ;
 wire \y_c[5].x_c[0].lc_i.cfg[5] ;
 wire \y_c[5].x_c[0].lc_i.cfg[6] ;
 wire \y_c[5].x_c[0].lc_i.cfg[7] ;
 wire \y_c[5].x_c[0].lc_i.cfg_strb[0] ;
 wire \y_c[5].x_c[0].lc_i.cfg_strb[1] ;
 wire \y_c[5].x_c[0].lc_i.dff.dffo_n ;
 wire \y_c[5].x_c[0].lc_i.i0 ;
 wire \y_c[5].x_c[0].lc_i.i0a ;
 wire \y_c[5].x_c[0].lc_i.i0b ;
 wire \y_c[5].x_c[0].lc_i.i1 ;
 wire \y_c[5].x_c[0].lc_i.i1a ;
 wire \y_c[5].x_c[0].lc_i.i1b ;
 wire \y_c[5].x_c[0].lc_i.muxo_n ;
 wire \y_c[5].x_c[0].lc_i.s0 ;
 wire \y_c[5].x_c[0].lc_i.s0a ;
 wire \y_c[5].x_c[0].lc_i.s0b ;
 wire \y_c[5].x_c[0].lc_i.s0s ;
 wire \y_c[5].x_c[1].lc_i.cfg[0] ;
 wire \y_c[5].x_c[1].lc_i.cfg[1] ;
 wire \y_c[5].x_c[1].lc_i.cfg[2] ;
 wire \y_c[5].x_c[1].lc_i.cfg[3] ;
 wire \y_c[5].x_c[1].lc_i.cfg[4] ;
 wire \y_c[5].x_c[1].lc_i.cfg[5] ;
 wire \y_c[5].x_c[1].lc_i.cfg[6] ;
 wire \y_c[5].x_c[1].lc_i.cfg[7] ;
 wire \y_c[5].x_c[1].lc_i.dff.dffo_n ;
 wire \y_c[5].x_c[1].lc_i.i0 ;
 wire \y_c[5].x_c[1].lc_i.i0a ;
 wire \y_c[5].x_c[1].lc_i.i0b ;
 wire \y_c[5].x_c[1].lc_i.i1 ;
 wire \y_c[5].x_c[1].lc_i.i1a ;
 wire \y_c[5].x_c[1].lc_i.i1b ;
 wire \y_c[5].x_c[1].lc_i.muxo_n ;
 wire \y_c[5].x_c[1].lc_i.s0 ;
 wire \y_c[5].x_c[1].lc_i.s0a ;
 wire \y_c[5].x_c[1].lc_i.s0b ;
 wire \y_c[5].x_c[1].lc_i.s0s ;
 wire \y_c[5].x_c[2].lc_i.cfg[0] ;
 wire \y_c[5].x_c[2].lc_i.cfg[1] ;
 wire \y_c[5].x_c[2].lc_i.cfg[2] ;
 wire \y_c[5].x_c[2].lc_i.cfg[3] ;
 wire \y_c[5].x_c[2].lc_i.cfg[4] ;
 wire \y_c[5].x_c[2].lc_i.cfg[5] ;
 wire \y_c[5].x_c[2].lc_i.cfg[6] ;
 wire \y_c[5].x_c[2].lc_i.cfg[7] ;
 wire \y_c[5].x_c[2].lc_i.dff.dffo_n ;
 wire \y_c[5].x_c[2].lc_i.i0 ;
 wire \y_c[5].x_c[2].lc_i.i0a ;
 wire \y_c[5].x_c[2].lc_i.i0b ;
 wire \y_c[5].x_c[2].lc_i.i1 ;
 wire \y_c[5].x_c[2].lc_i.i1a ;
 wire \y_c[5].x_c[2].lc_i.i1b ;
 wire \y_c[5].x_c[2].lc_i.muxo_n ;
 wire \y_c[5].x_c[2].lc_i.s0 ;
 wire \y_c[5].x_c[2].lc_i.s0a ;
 wire \y_c[5].x_c[2].lc_i.s0b ;
 wire \y_c[5].x_c[2].lc_i.s0s ;
 wire \y_c[5].x_c[3].lc_i.cfg[0] ;
 wire \y_c[5].x_c[3].lc_i.cfg[1] ;
 wire \y_c[5].x_c[3].lc_i.cfg[2] ;
 wire \y_c[5].x_c[3].lc_i.cfg[3] ;
 wire \y_c[5].x_c[3].lc_i.cfg[4] ;
 wire \y_c[5].x_c[3].lc_i.cfg[5] ;
 wire \y_c[5].x_c[3].lc_i.cfg[6] ;
 wire \y_c[5].x_c[3].lc_i.cfg[7] ;
 wire \y_c[5].x_c[3].lc_i.dff.dffo_n ;
 wire \y_c[5].x_c[3].lc_i.i0 ;
 wire \y_c[5].x_c[3].lc_i.i0a ;
 wire \y_c[5].x_c[3].lc_i.i0b ;
 wire \y_c[5].x_c[3].lc_i.i1 ;
 wire \y_c[5].x_c[3].lc_i.i1a ;
 wire \y_c[5].x_c[3].lc_i.i1b ;
 wire \y_c[5].x_c[3].lc_i.muxo_n ;
 wire \y_c[5].x_c[3].lc_i.s0 ;
 wire \y_c[5].x_c[3].lc_i.s0a ;
 wire \y_c[5].x_c[3].lc_i.s0b ;
 wire \y_c[5].x_c[3].lc_i.s0s ;
 wire \y_c[5].x_c[4].lc_i.cfg[0] ;
 wire \y_c[5].x_c[4].lc_i.cfg[1] ;
 wire \y_c[5].x_c[4].lc_i.cfg[2] ;
 wire \y_c[5].x_c[4].lc_i.cfg[3] ;
 wire \y_c[5].x_c[4].lc_i.cfg[4] ;
 wire \y_c[5].x_c[4].lc_i.cfg[5] ;
 wire \y_c[5].x_c[4].lc_i.cfg[6] ;
 wire \y_c[5].x_c[4].lc_i.cfg[7] ;
 wire \y_c[5].x_c[4].lc_i.dff.dffo_n ;
 wire \y_c[5].x_c[4].lc_i.i0 ;
 wire \y_c[5].x_c[4].lc_i.i0a ;
 wire \y_c[5].x_c[4].lc_i.i0b ;
 wire \y_c[5].x_c[4].lc_i.i1 ;
 wire \y_c[5].x_c[4].lc_i.i1a ;
 wire \y_c[5].x_c[4].lc_i.i1b ;
 wire \y_c[5].x_c[4].lc_i.muxo_n ;
 wire \y_c[5].x_c[4].lc_i.s0 ;
 wire \y_c[5].x_c[4].lc_i.s0a ;
 wire \y_c[5].x_c[4].lc_i.s0b ;
 wire \y_c[5].x_c[4].lc_i.s0s ;
 wire [0:0] clknet_0_io_in;
 wire [0:0] clknet_2_0__leaf_io_in;
 wire [0:0] clknet_2_1__leaf_io_in;
 wire [0:0] clknet_2_2__leaf_io_in;
 wire [0:0] clknet_2_3__leaf_io_in;

 sky130_fd_sc_hd__diode_2 ANTENNA_0 (.DIODE(io_in[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(io_in[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(cfg_datain),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(io_in[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(io_in[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_15_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_25_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_29_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\y_c[2].x_c[1].lc_i.muxo_n ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_13_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_10_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_272 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_284 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_10_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_10_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_10_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_11_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_11_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_11_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_284 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_11_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_11_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_12_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_13_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_13_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_13_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_14_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_14_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_263 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_275 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_287 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_14_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_15_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_15_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_15_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_15_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_15_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_16_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_16_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_17_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_17_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_18_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_18_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_270 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_282 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_18_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_18_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_241 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_1_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_1_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_20_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_224 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_20_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_256 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_20_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_283 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_20_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_20_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_20_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_21_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_254 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_21_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_21_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_21_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_22_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_256 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_268 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_280 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_23_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_266 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_23_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_24_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_263 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_275 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_287 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_24_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_25_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_255 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_25_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_25_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_25_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_256 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_290 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_26_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_27_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_27_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_254 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_266 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_278 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_290 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_29_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_245 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_29_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_2_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_30_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_262 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_31_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_31_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_32_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_32_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_32_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_32_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_32_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_33_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_33_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_33_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_33_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_33_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_33_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_170 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_219 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_231 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_35_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_35_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_35_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_202 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_35_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_35_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_35_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_35_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_248 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_35_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_36_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_36_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_36_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_235 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_36_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_36_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_37_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_37_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_37_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_37_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_38_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_173 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_38_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_38_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_238 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_270 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_282 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_38_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_39_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_255 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_267 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_3_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_3_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_40_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_40_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_40_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_40_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_40_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_40_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_41_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_200 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_212 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_41_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_42_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_42_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_42_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_43_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_44_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_44_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_44_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_44_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_44_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_44_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_195 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_239 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_251 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_263 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_45_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_45_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_46_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_46_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_46_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_46_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_46_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_192 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_204 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_47_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_47_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_213 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_48_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_48_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_49_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_49_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_187 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_256 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_268 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_280 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_4_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_50_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_50_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_50_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_50_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_50_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_50_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_51_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_51_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_212 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_217 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_52_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_53_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_198 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_210 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_53_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_53_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_151 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_163 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_175 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_54_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_54_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_54_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_54_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_144 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_156 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_55_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_55_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_56_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_155 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_167 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_179 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_56_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_56_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_56_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_56_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_123 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_57_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_57_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_5_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_5_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_256 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_268 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_5_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_5_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_6_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_7_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_267 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_7_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_8_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_8_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_256 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_268 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_280 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_8_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_8_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_9_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_254 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_9_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_268 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 _33_ (.A(\frame_ctr[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_17_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _34_ (.A(\frame_ctr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_18_));
 sky130_fd_sc_hd__or2_1 _35_ (.A(_17_),
    .B(_18_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_19_));
 sky130_fd_sc_hd__clkbuf_1 _36_ (.A(\frame_ctr[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_20_));
 sky130_fd_sc_hd__or2_1 _37_ (.A(\frame_ctr[3] ),
    .B(_20_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_21_));
 sky130_fd_sc_hd__nor2_1 _38_ (.A(_19_),
    .B(_21_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_00_));
 sky130_fd_sc_hd__nand2b_1 _39_ (.A_N(_17_),
    .B(\frame_ctr[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_22_));
 sky130_fd_sc_hd__nor2_1 _40_ (.A(_21_),
    .B(_22_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_01_));
 sky130_fd_sc_hd__or2b_1 _41_ (.A(\frame_ctr[0] ),
    .B_N(\frame_ctr[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_23_));
 sky130_fd_sc_hd__nor2_1 _42_ (.A(_21_),
    .B(_23_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02_));
 sky130_fd_sc_hd__clkbuf_2 _43_ (.A(\frame_ctr[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_24_));
 sky130_fd_sc_hd__and4bb_1 _44_ (.A_N(_24_),
    .B_N(_20_),
    .C(_17_),
    .D(_18_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_25_));
 sky130_fd_sc_hd__clkbuf_1 _45_ (.A(_25_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03_));
 sky130_fd_sc_hd__or2b_1 _46_ (.A(\frame_ctr[3] ),
    .B_N(_20_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_26_));
 sky130_fd_sc_hd__nor2_1 _47_ (.A(_19_),
    .B(_26_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04_));
 sky130_fd_sc_hd__nor2_1 _48_ (.A(_22_),
    .B(_26_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_05_));
 sky130_fd_sc_hd__nor2_1 _49_ (.A(_23_),
    .B(_26_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_06_));
 sky130_fd_sc_hd__and3_1 _50_ (.A(\frame_ctr[1] ),
    .B(\frame_ctr[0] ),
    .C(\frame_ctr[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_27_));
 sky130_fd_sc_hd__and2b_1 _51_ (.A_N(_24_),
    .B(_27_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_28_));
 sky130_fd_sc_hd__clkbuf_1 _52_ (.A(_28_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_07_));
 sky130_fd_sc_hd__or2b_1 _53_ (.A(\frame_ctr[2] ),
    .B_N(_24_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_29_));
 sky130_fd_sc_hd__nor2_1 _54_ (.A(_19_),
    .B(_29_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_08_));
 sky130_fd_sc_hd__nor2_1 _55_ (.A(_22_),
    .B(_29_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_09_));
 sky130_fd_sc_hd__nor2_1 _56_ (.A(_23_),
    .B(_29_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_10_));
 sky130_fd_sc_hd__and4b_1 _57_ (.A_N(_20_),
    .B(_24_),
    .C(_18_),
    .D(_17_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_30_));
 sky130_fd_sc_hd__clkbuf_1 _58_ (.A(_30_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_11_));
 sky130_fd_sc_hd__clkinv_4 _59_ (.A(\y_c[0].x_c[0].lc_i.cfg_mode ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_12_));
 sky130_fd_sc_hd__and2_1 _60_ (.A(\y_c[0].x_c[0].lc_i.cfg_mode ),
    .B(cfg_framestrb),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_31_));
 sky130_fd_sc_hd__clkbuf_1 _61_ (.A(_31_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(gated_strobe));
 sky130_fd_sc_hd__nand2_1 _62_ (.A(_22_),
    .B(_23_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_14_));
 sky130_fd_sc_hd__a21oi_1 _63_ (.A1(_17_),
    .A2(_18_),
    .B1(_20_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_32_));
 sky130_fd_sc_hd__nor2_1 _64_ (.A(_27_),
    .B(_32_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_15_));
 sky130_fd_sc_hd__xor2_1 _65_ (.A(_24_),
    .B(_27_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_16_));
 sky130_fd_sc_hd__inv_2 _66_ (.A(_18_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_13_));
 sky130_fd_sc_hd__dfrtp_1 _67_ (.CLK(cfg_frameinc),
    .D(_13_),
    .RESET_B(\y_c[0].x_c[0].lc_i.cfg_mode ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\frame_ctr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _68_ (.CLK(cfg_frameinc),
    .D(_14_),
    .RESET_B(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\frame_ctr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _69_ (.CLK(cfg_frameinc),
    .D(_15_),
    .RESET_B(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\frame_ctr[2] ));
 sky130_fd_sc_hd__dfrtp_1 _70_ (.CLK(cfg_frameinc),
    .D(_16_),
    .RESET_B(net145),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\frame_ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _71_ (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(\y_c[0].x_c[0].lc_i.cfg_data[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _72_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(\y_c[0].x_c[0].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _73_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[0].x_c[0].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _74_ (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(\y_c[0].x_c[1].lc_i.cfg_data[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _75_ (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _76_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _77_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _78_ (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(\y_c[0].x_c[2].lc_i.cfg_data[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _79_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[0].x_c[2].lc_i.cfg_data[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _80_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _81_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[0].x_c[2].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _82_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(\y_c[0].x_c[3].lc_i.cfg_data[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _83_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(net169),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _84_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[0].x_c[3].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _85_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[0].x_c[3].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _86_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[0].x_c[4].lc_i.cfg_data[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _87_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[0].x_c[4].lc_i.cfg_data[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _88_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(\y_c[0].x_c[4].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _89_ (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[0].x_c[4].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _90_ (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(cfg_datain),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg_data[3] ));
 sky130_fd_sc_hd__buf_2 _91_ (.A(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 _92_ (.A(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_2 _93_ (.A(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_2 _94_ (.A(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_2 _95_ (.A(\y_c[4].x_c[0].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 _96_ (.A(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 _97_ (.A(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_2 _98_ (.A(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[7]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_io_in[0]  (.A(io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_2_0__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_2_1__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_2_2__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_2_3__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_2 din_buf (.A(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(cfg_datain));
 sky130_fd_sc_hd__clkbuf_1 \din_buf[0]  (.A(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[0].x_c[0].lc_i.T ));
 sky130_fd_sc_hd__clkbuf_2 \din_buf[1]  (.A(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[0].x_c[0].lc_i.L ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \din_buf[2]  (.A(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[0].x_c[2].lc_i.T ));
 sky130_fd_sc_hd__clkbuf_2 \din_buf[3]  (.A(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[0].x_c[3].lc_i.T ));
 sky130_fd_sc_hd__clkbuf_2 \din_buf[4]  (.A(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[0].x_c[4].lc_i.T ));
 sky130_fd_sc_hd__clkbuf_1 \din_buf[5]  (.A(net6),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[4].x_c[0].lc_i.L ));
 sky130_fd_sc_hd__clkbuf_1 \din_buf[6]  (.A(net7),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[5].x_c[0].lc_i.L ));
 sky130_fd_sc_hd__clkbuf_2 frameinc_clkbuf (.A(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(cfg_frameinc));
 sky130_fd_sc_hd__clkbuf_1 framestrb_clkbuf (.A(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(cfg_framestrb));
 sky130_fd_sc_hd__nand2_1 \genblk1[0].cfg_nand  (.A(net133),
    .B(_00_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.cfg_strb[0] ));
 sky130_fd_sc_hd__nand2_1 \genblk1[10].cfg_nand  (.A(net134),
    .B(_10_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.cfg_strb[0] ));
 sky130_fd_sc_hd__nand2_1 \genblk1[11].cfg_nand  (.A(net134),
    .B(_11_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.cfg_strb[1] ));
 sky130_fd_sc_hd__nand2_1 \genblk1[1].cfg_nand  (.A(net133),
    .B(_01_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.cfg_strb[1] ));
 sky130_fd_sc_hd__nand2_1 \genblk1[2].cfg_nand  (.A(net135),
    .B(_02_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.cfg_strb[0] ));
 sky130_fd_sc_hd__nand2_1 \genblk1[3].cfg_nand  (.A(net133),
    .B(_03_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.cfg_strb[1] ));
 sky130_fd_sc_hd__nand2_1 \genblk1[4].cfg_nand  (.A(net135),
    .B(_04_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.cfg_strb[0] ));
 sky130_fd_sc_hd__nand2_1 \genblk1[5].cfg_nand  (.A(net133),
    .B(_05_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.cfg_strb[1] ));
 sky130_fd_sc_hd__nand2_1 \genblk1[6].cfg_nand  (.A(gated_strobe),
    .B(_06_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.cfg_strb[0] ));
 sky130_fd_sc_hd__nand2_1 \genblk1[7].cfg_nand  (.A(net135),
    .B(_07_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.cfg_strb[1] ));
 sky130_fd_sc_hd__nand2_1 \genblk1[8].cfg_nand  (.A(net134),
    .B(_08_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.cfg_strb[0] ));
 sky130_fd_sc_hd__nand2_1 \genblk1[9].cfg_nand  (.A(net134),
    .B(_09_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.cfg_strb[1] ));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\y_c[0].x_c[1].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\y_c[0].x_c[1].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(io_in[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(io_in[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 mode_clkbuf (.A(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[0].x_c[0].lc_i.cfg_mode ));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater10 (.A(\y_c[3].x_c[4].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 repeater100 (.A(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 repeater101 (.A(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 repeater102 (.A(\y_c[1].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 repeater103 (.A(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 repeater104 (.A(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 repeater105 (.A(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 repeater106 (.A(net107),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 repeater107 (.A(net108),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 repeater108 (.A(\y_c[1].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 repeater109 (.A(net110),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 repeater11 (.A(\y_c[3].x_c[4].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 repeater110 (.A(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net110));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater111 (.A(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 repeater112 (.A(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net112));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater113 (.A(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 repeater114 (.A(\y_c[0].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 repeater115 (.A(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 repeater116 (.A(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 repeater117 (.A(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 repeater118 (.A(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 repeater119 (.A(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net119));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater12 (.A(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 repeater120 (.A(\y_c[5].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 repeater121 (.A(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 repeater122 (.A(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 repeater123 (.A(net124),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 repeater124 (.A(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 repeater125 (.A(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 repeater126 (.A(\y_c[5].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 repeater127 (.A(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 repeater128 (.A(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 repeater129 (.A(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 repeater13 (.A(\y_c[3].x_c[1].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 repeater130 (.A(net132),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 repeater131 (.A(net132),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 repeater132 (.A(\y_c[0].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 repeater133 (.A(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 repeater134 (.A(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 repeater135 (.A(gated_strobe),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 repeater136 (.A(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 repeater137 (.A(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net137));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater138 (.A(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net138));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater139 (.A(net140),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 repeater14 (.A(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater140 (.A(net141),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net140));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater141 (.A(_12_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 repeater142 (.A(net143),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net142));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater143 (.A(net144),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 repeater144 (.A(_12_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 repeater145 (.A(\y_c[0].x_c[0].lc_i.cfg_mode ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 repeater146 (.A(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 repeater147 (.A(\y_c[0].x_c[4].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 repeater148 (.A(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 repeater149 (.A(\y_c[0].x_c[4].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 repeater15 (.A(\y_c[2].x_c[4].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 repeater150 (.A(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net150));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater151 (.A(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 repeater152 (.A(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net152));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater153 (.A(\y_c[0].x_c[4].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 repeater154 (.A(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 repeater155 (.A(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 repeater156 (.A(\y_c[0].x_c[4].lc_i.cfg_data[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 repeater157 (.A(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net157));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater158 (.A(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net158));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater159 (.A(\y_c[0].x_c[4].lc_i.cfg_data[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 repeater16 (.A(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 repeater160 (.A(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 repeater161 (.A(net163),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 repeater162 (.A(net163),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 repeater163 (.A(\y_c[0].x_c[3].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net163));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater164 (.A(net165),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net164));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater165 (.A(\y_c[0].x_c[3].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 repeater166 (.A(\y_c[0].x_c[3].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 repeater167 (.A(net169),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 repeater168 (.A(\y_c[0].x_c[3].lc_i.cfg_data[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 repeater169 (.A(\y_c[0].x_c[3].lc_i.cfg_data[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net169));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater17 (.A(\y_c[3].x_c[2].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 repeater170 (.A(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 repeater171 (.A(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 repeater172 (.A(\y_c[0].x_c[3].lc_i.cfg_data[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net172));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater173 (.A(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 repeater174 (.A(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net174));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater175 (.A(\y_c[0].x_c[2].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net175));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater176 (.A(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 repeater177 (.A(\y_c[0].x_c[2].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 repeater178 (.A(\y_c[0].x_c[2].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 repeater179 (.A(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net179));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater18 (.A(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater180 (.A(\y_c[0].x_c[2].lc_i.cfg_data[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 repeater181 (.A(\y_c[0].x_c[2].lc_i.cfg_data[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net181));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater182 (.A(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net182));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater183 (.A(\y_c[0].x_c[2].lc_i.cfg_data[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_2 repeater184 (.A(\y_c[0].x_c[2].lc_i.cfg_data[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 repeater185 (.A(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 repeater186 (.A(net187),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 repeater187 (.A(net188),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_2 repeater188 (.A(\y_c[0].x_c[1].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 repeater189 (.A(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net189));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater19 (.A(\y_c[2].x_c[3].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 repeater190 (.A(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 repeater191 (.A(\y_c[0].x_c[1].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 repeater192 (.A(\y_c[0].x_c[1].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_2 repeater193 (.A(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 repeater194 (.A(\y_c[0].x_c[1].lc_i.cfg_data[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 repeater195 (.A(\y_c[0].x_c[1].lc_i.cfg_data[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 repeater196 (.A(net198),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 repeater197 (.A(net198),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 repeater198 (.A(\y_c[0].x_c[1].lc_i.cfg_data[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 repeater199 (.A(net200),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 repeater20 (.A(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 repeater200 (.A(\y_c[0].x_c[0].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 repeater201 (.A(\y_c[0].x_c[0].lc_i.cfg_data[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net201));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater202 (.A(\y_c[0].x_c[0].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 repeater203 (.A(net204),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 repeater204 (.A(\y_c[0].x_c[0].lc_i.cfg_data[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net204));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater205 (.A(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 repeater206 (.A(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 repeater207 (.A(\y_c[0].x_c[0].lc_i.cfg_data[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 repeater208 (.A(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net208));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater209 (.A(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 repeater21 (.A(\y_c[3].x_c[3].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 repeater210 (.A(\y_c[0].x_c[0].lc_i.cfg_data[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net210));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater22 (.A(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 repeater23 (.A(\y_c[4].x_c[3].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 repeater24 (.A(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 repeater25 (.A(\y_c[4].x_c[2].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 repeater26 (.A(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater27 (.A(\y_c[4].x_c[1].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 repeater28 (.A(\y_c[4].x_c[0].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater29 (.A(\y_c[3].x_c[0].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 repeater30 (.A(\y_c[2].x_c[0].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater31 (.A(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 repeater32 (.A(\y_c[2].x_c[1].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater33 (.A(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 repeater34 (.A(\y_c[2].x_c[2].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 repeater35 (.A(\y_c[1].x_c[2].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 repeater36 (.A(\y_c[1].x_c[2].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 repeater37 (.A(\y_c[1].x_c[1].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 repeater38 (.A(\y_c[1].x_c[1].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 repeater39 (.A(\y_c[1].x_c[0].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 repeater40 (.A(\y_c[0].x_c[0].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 repeater41 (.A(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 repeater42 (.A(\y_c[0].x_c[1].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 repeater43 (.A(\y_c[0].x_c[2].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 repeater44 (.A(\y_c[0].x_c[2].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 repeater45 (.A(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 repeater46 (.A(\y_c[0].x_c[3].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 repeater47 (.A(\y_c[1].x_c[3].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 repeater48 (.A(\y_c[1].x_c[3].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater49 (.A(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 repeater50 (.A(\y_c[1].x_c[4].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 repeater51 (.A(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 repeater52 (.A(\y_c[0].x_c[4].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 repeater53 (.A(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 repeater54 (.A(\y_c[0].x_c[3].lc_i.R ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net54));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater55 (.A(\y_c[0].x_c[2].lc_i.R ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 repeater56 (.A(\y_c[0].x_c[2].lc_i.R ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 repeater57 (.A(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater58 (.A(\y_c[0].x_c[1].lc_i.R ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 repeater59 (.A(\y_c[0].x_c[0].lc_i.R ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 repeater60 (.A(\y_c[0].x_c[0].lc_i.R ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 repeater61 (.A(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 repeater62 (.A(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 repeater63 (.A(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 repeater64 (.A(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater65 (.A(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 repeater66 (.A(\y_c[4].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 repeater67 (.A(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 repeater68 (.A(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 repeater69 (.A(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 repeater70 (.A(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 repeater71 (.A(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 repeater72 (.A(\y_c[4].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 repeater73 (.A(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 repeater74 (.A(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 repeater75 (.A(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 repeater76 (.A(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 repeater77 (.A(\y_c[3].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 repeater78 (.A(\y_c[3].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 repeater79 (.A(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 repeater8 (.A(\y_c[4].x_c[4].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 repeater80 (.A(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 repeater81 (.A(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 repeater82 (.A(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 repeater83 (.A(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 repeater84 (.A(\y_c[3].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 repeater85 (.A(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net85));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater86 (.A(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 repeater87 (.A(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 repeater88 (.A(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 repeater89 (.A(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 repeater9 (.A(\y_c[4].x_c[4].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 repeater90 (.A(\y_c[2].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 repeater91 (.A(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 repeater92 (.A(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 repeater93 (.A(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 repeater94 (.A(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 repeater95 (.A(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 repeater96 (.A(\y_c[2].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 repeater97 (.A(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 repeater98 (.A(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 repeater99 (.A(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net99));
 sky130_fd_sc_hd__dfsbp_1 \y_c[0].x_c[0].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[0].x_c[0].lc_i.muxo_n ),
    .SET_B(net141),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[0].x_c[0].lc_i.dff.ffsel  (.A0(\y_c[0].x_c[0].lc_i.muxo_n ),
    .A1(\y_c[0].x_c[0].lc_i.dff.dffo_n ),
    .S(\y_c[0].x_c[0].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.Q ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[0].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net208),
    .GATE_N(\y_c[0].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[0].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net205),
    .GATE_N(net132),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[0].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net203),
    .GATE_N(net132),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[0].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net200),
    .GATE_N(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[0].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net208),
    .GATE_N(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[0].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net205),
    .GATE_N(\y_c[0].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[0].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net204),
    .GATE_N(net110),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[0].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net200),
    .GATE_N(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[0].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[0].x_c[0].lc_i.i0muxa0  (.A(\y_c[0].x_c[0].lc_i.T ),
    .B(\y_c[0].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_2 \y_c[0].x_c[0].lc_i.i0muxa1  (.A0(net59),
    .A1(\y_c[0].x_c[0].lc_i.L ),
    .S(\y_c[0].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_4 \y_c[0].x_c[0].lc_i.i0muxb  (.A0(\y_c[0].x_c[0].lc_i.i0a ),
    .A1(\y_c[0].x_c[0].lc_i.i0b ),
    .S(\y_c[0].x_c[0].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[0].x_c[0].lc_i.i1muxa0  (.A(\y_c[0].x_c[0].lc_i.cfg[2] ),
    .B(\y_c[0].x_c[0].lc_i.L ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[0].x_c[0].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_2 \y_c[0].x_c[0].lc_i.i1muxa1  (.A0(net40),
    .A1(net59),
    .S(\y_c[0].x_c[0].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_4 \y_c[0].x_c[0].lc_i.i1muxb  (.A0(\y_c[0].x_c[0].lc_i.i1a ),
    .A1(\y_c[0].x_c[0].lc_i.i1b ),
    .S(\y_c[0].x_c[0].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[0].x_c[0].lc_i.lmux  (.A0(\y_c[0].x_c[0].lc_i.i0 ),
    .A1(\y_c[0].x_c[0].lc_i.i1 ),
    .S(\y_c[0].x_c[0].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[0].x_c[0].lc_i.s0muxa0  (.A(\y_c[0].x_c[0].lc_i.T ),
    .B(\y_c[0].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_2 \y_c[0].x_c[0].lc_i.s0muxa1  (.A0(net59),
    .A1(\y_c[0].x_c[0].lc_i.L ),
    .S(\y_c[0].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[0].x_c[0].lc_i.s0muxb  (.A0(\y_c[0].x_c[0].lc_i.s0a ),
    .A1(\y_c[0].x_c[0].lc_i.s0b ),
    .S(\y_c[0].x_c[0].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[0].x_c[0].lc_i.sinv  (.A(\y_c[0].x_c[0].lc_i.s0s ),
    .B(\y_c[0].x_c[0].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[0].x_c[1].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[0].x_c[1].lc_i.muxo_n ),
    .SET_B(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_2 \y_c[0].x_c[1].lc_i.dff.ffsel  (.A0(\y_c[0].x_c[1].lc_i.muxo_n ),
    .A1(\y_c[0].x_c[1].lc_i.dff.dffo_n ),
    .S(\y_c[0].x_c[1].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.R ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[1].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net197),
    .GATE_N(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[1].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net194),
    .GATE_N(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[1].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net189),
    .GATE_N(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[1].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net186),
    .GATE_N(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[1].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net197),
    .GATE_N(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[1].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net194),
    .GATE_N(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[1].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net189),
    .GATE_N(net110),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[1].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net185),
    .GATE_N(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[1].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[0].x_c[1].lc_i.i0muxa0  (.A(\y_c[0].x_c[0].lc_i.L ),
    .B(\y_c[0].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[1].lc_i.i0muxa1  (.A0(net58),
    .A1(\y_c[0].x_c[0].lc_i.Q ),
    .S(\y_c[0].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[0].x_c[1].lc_i.i0muxb  (.A0(\y_c[0].x_c[1].lc_i.i0a ),
    .A1(\y_c[0].x_c[1].lc_i.i0b ),
    .S(\y_c[0].x_c[1].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[0].x_c[1].lc_i.i1muxa0  (.A(\y_c[0].x_c[1].lc_i.cfg[2] ),
    .B(\y_c[0].x_c[0].lc_i.Q ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[0].x_c[1].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[1].lc_i.i1muxa1  (.A0(net41),
    .A1(net58),
    .S(\y_c[0].x_c[1].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[1].lc_i.i1muxb  (.A0(\y_c[0].x_c[1].lc_i.i1a ),
    .A1(\y_c[0].x_c[1].lc_i.i1b ),
    .S(\y_c[0].x_c[1].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[0].x_c[1].lc_i.lmux  (.A0(\y_c[0].x_c[1].lc_i.i0 ),
    .A1(\y_c[0].x_c[1].lc_i.i1 ),
    .S(\y_c[0].x_c[1].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[0].x_c[1].lc_i.s0muxa0  (.A(\y_c[0].x_c[0].lc_i.L ),
    .B(\y_c[0].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[1].lc_i.s0muxa1  (.A0(net58),
    .A1(\y_c[0].x_c[0].lc_i.Q ),
    .S(\y_c[0].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[1].lc_i.s0muxb  (.A0(\y_c[0].x_c[1].lc_i.s0a ),
    .A1(\y_c[0].x_c[1].lc_i.s0b ),
    .S(\y_c[0].x_c[1].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[0].x_c[1].lc_i.sinv  (.A(\y_c[0].x_c[1].lc_i.s0s ),
    .B(\y_c[0].x_c[1].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[0].x_c[2].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[0].x_c[2].lc_i.muxo_n ),
    .SET_B(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_2 \y_c[0].x_c[2].lc_i.dff.ffsel  (.A0(\y_c[0].x_c[2].lc_i.muxo_n ),
    .A1(\y_c[0].x_c[2].lc_i.dff.dffo_n ),
    .S(\y_c[0].x_c[2].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.R ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[2].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net184),
    .GATE_N(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[2].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net180),
    .GATE_N(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[2].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net177),
    .GATE_N(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[2].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net173),
    .GATE_N(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[2].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net184),
    .GATE_N(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[2].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net180),
    .GATE_N(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[2].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(\y_c[0].x_c[2].lc_i.cfg_data[2] ),
    .GATE_N(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[2].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net173),
    .GATE_N(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[2].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[0].x_c[2].lc_i.i0muxa0  (.A(\y_c[0].x_c[2].lc_i.T ),
    .B(\y_c[0].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[2].lc_i.i0muxa1  (.A0(net56),
    .A1(\y_c[0].x_c[0].lc_i.R ),
    .S(\y_c[0].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[2].lc_i.i0muxb  (.A0(\y_c[0].x_c[2].lc_i.i0a ),
    .A1(\y_c[0].x_c[2].lc_i.i0b ),
    .S(\y_c[0].x_c[2].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[0].x_c[2].lc_i.i1muxa0  (.A(\y_c[0].x_c[2].lc_i.cfg[2] ),
    .B(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[0].x_c[2].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[2].lc_i.i1muxa1  (.A0(net43),
    .A1(net56),
    .S(\y_c[0].x_c[2].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_4 \y_c[0].x_c[2].lc_i.i1muxb  (.A0(\y_c[0].x_c[2].lc_i.i1a ),
    .A1(\y_c[0].x_c[2].lc_i.i1b ),
    .S(\y_c[0].x_c[2].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[0].x_c[2].lc_i.lmux  (.A0(\y_c[0].x_c[2].lc_i.i0 ),
    .A1(\y_c[0].x_c[2].lc_i.i1 ),
    .S(\y_c[0].x_c[2].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[0].x_c[2].lc_i.s0muxa0  (.A(\y_c[0].x_c[2].lc_i.T ),
    .B(\y_c[0].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[2].lc_i.s0muxa1  (.A0(net56),
    .A1(net60),
    .S(\y_c[0].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[2].lc_i.s0muxb  (.A0(\y_c[0].x_c[2].lc_i.s0a ),
    .A1(\y_c[0].x_c[2].lc_i.s0b ),
    .S(\y_c[0].x_c[2].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[0].x_c[2].lc_i.sinv  (.A(\y_c[0].x_c[2].lc_i.s0s ),
    .B(\y_c[0].x_c[2].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[0].x_c[3].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[0].x_c[3].lc_i.muxo_n ),
    .SET_B(net136),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_2 \y_c[0].x_c[3].lc_i.dff.ffsel  (.A0(\y_c[0].x_c[3].lc_i.muxo_n ),
    .A1(\y_c[0].x_c[3].lc_i.dff.dffo_n ),
    .S(\y_c[0].x_c[3].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.R ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[3].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net170),
    .GATE_N(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[3].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(\y_c[0].x_c[3].lc_i.cfg_data[1] ),
    .GATE_N(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[3].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net166),
    .GATE_N(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[3].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net162),
    .GATE_N(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[3].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net170),
    .GATE_N(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[3].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(\y_c[0].x_c[3].lc_i.cfg_data[1] ),
    .GATE_N(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[3].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net166),
    .GATE_N(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[3].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net163),
    .GATE_N(net110),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[3].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[0].x_c[3].lc_i.i0muxa0  (.A(\y_c[0].x_c[3].lc_i.T ),
    .B(\y_c[0].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[3].lc_i.i0muxa1  (.A0(net54),
    .A1(\y_c[0].x_c[1].lc_i.R ),
    .S(\y_c[0].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[0].x_c[3].lc_i.i0muxb  (.A0(\y_c[0].x_c[3].lc_i.i0a ),
    .A1(\y_c[0].x_c[3].lc_i.i0b ),
    .S(\y_c[0].x_c[3].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[0].x_c[3].lc_i.i1muxa0  (.A(\y_c[0].x_c[3].lc_i.cfg[2] ),
    .B(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[0].x_c[3].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[3].lc_i.i1muxa1  (.A0(net45),
    .A1(\y_c[0].x_c[3].lc_i.R ),
    .S(\y_c[0].x_c[3].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[3].lc_i.i1muxb  (.A0(\y_c[0].x_c[3].lc_i.i1a ),
    .A1(\y_c[0].x_c[3].lc_i.i1b ),
    .S(\y_c[0].x_c[3].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[0].x_c[3].lc_i.lmux  (.A0(\y_c[0].x_c[3].lc_i.i0 ),
    .A1(\y_c[0].x_c[3].lc_i.i1 ),
    .S(\y_c[0].x_c[3].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[0].x_c[3].lc_i.s0muxa0  (.A(\y_c[0].x_c[3].lc_i.T ),
    .B(\y_c[0].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[3].lc_i.s0muxa1  (.A0(\y_c[0].x_c[3].lc_i.R ),
    .A1(\y_c[0].x_c[1].lc_i.R ),
    .S(\y_c[0].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[3].lc_i.s0muxb  (.A0(\y_c[0].x_c[3].lc_i.s0a ),
    .A1(\y_c[0].x_c[3].lc_i.s0b ),
    .S(\y_c[0].x_c[3].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[0].x_c[3].lc_i.sinv  (.A(\y_c[0].x_c[3].lc_i.s0s ),
    .B(\y_c[0].x_c[3].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[0].x_c[4].lc_i.dff.dff  (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[0].x_c[4].lc_i.muxo_n ),
    .SET_B(net140),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_2 \y_c[0].x_c[4].lc_i.dff.ffsel  (.A0(\y_c[0].x_c[4].lc_i.muxo_n ),
    .A1(\y_c[0].x_c[4].lc_i.dff.dffo_n ),
    .S(\y_c[0].x_c[4].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.R ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[4].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net157),
    .GATE_N(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[4].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net154),
    .GATE_N(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[4].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net150),
    .GATE_N(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[4].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net147),
    .GATE_N(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[4].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net157),
    .GATE_N(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[4].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net154),
    .GATE_N(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[4].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net150),
    .GATE_N(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[0].x_c[4].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net146),
    .GATE_N(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[0].x_c[4].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[0].x_c[4].lc_i.i0muxa0  (.A(\y_c[0].x_c[4].lc_i.T ),
    .B(\y_c[0].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[4].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[4].lc_i.i0muxa1  (.A0(net54),
    .A1(\y_c[0].x_c[2].lc_i.R ),
    .S(\y_c[0].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[4].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[0].x_c[4].lc_i.i0muxb  (.A0(\y_c[0].x_c[4].lc_i.i0a ),
    .A1(\y_c[0].x_c[4].lc_i.i0b ),
    .S(\y_c[0].x_c[4].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[4].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[0].x_c[4].lc_i.i1muxa0  (.A(\y_c[0].x_c[4].lc_i.cfg[2] ),
    .B(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[0].x_c[4].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[4].lc_i.i1muxa1  (.A0(net52),
    .A1(net53),
    .S(\y_c[0].x_c[4].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[4].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[4].lc_i.i1muxb  (.A0(\y_c[0].x_c[4].lc_i.i1a ),
    .A1(\y_c[0].x_c[4].lc_i.i1b ),
    .S(\y_c[0].x_c[4].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[4].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[0].x_c[4].lc_i.lmux  (.A0(\y_c[0].x_c[4].lc_i.i0 ),
    .A1(\y_c[0].x_c[4].lc_i.i1 ),
    .S(\y_c[0].x_c[4].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[4].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[0].x_c[4].lc_i.s0muxa0  (.A(\y_c[0].x_c[4].lc_i.T ),
    .B(\y_c[0].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[4].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[4].lc_i.s0muxa1  (.A0(net53),
    .A1(net55),
    .S(\y_c[0].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[4].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[0].x_c[4].lc_i.s0muxb  (.A0(\y_c[0].x_c[4].lc_i.s0a ),
    .A1(\y_c[0].x_c[4].lc_i.s0b ),
    .S(\y_c[0].x_c[4].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[4].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[0].x_c[4].lc_i.sinv  (.A(\y_c[0].x_c[4].lc_i.s0s ),
    .B(\y_c[0].x_c[4].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[4].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[1].x_c[0].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[1].x_c[0].lc_i.muxo_n ),
    .SET_B(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[0].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_2 \y_c[1].x_c[0].lc_i.dff.ffsel  (.A0(\y_c[1].x_c[0].lc_i.muxo_n ),
    .A1(\y_c[1].x_c[0].lc_i.dff.dffo_n ),
    .S(\y_c[1].x_c[0].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[0].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[0].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net209),
    .GATE_N(net108),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[0].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[0].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net205),
    .GATE_N(net108),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[0].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[0].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net204),
    .GATE_N(net107),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[0].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[0].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net200),
    .GATE_N(\y_c[1].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[0].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[0].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net209),
    .GATE_N(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[0].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[0].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net205),
    .GATE_N(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[0].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[0].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net204),
    .GATE_N(\y_c[1].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[0].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[0].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net199),
    .GATE_N(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[0].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[1].x_c[0].lc_i.i0muxa0  (.A(\y_c[0].x_c[0].lc_i.Q ),
    .B(\y_c[1].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[0].lc_i.i0muxa1  (.A0(net41),
    .A1(\y_c[0].x_c[2].lc_i.T ),
    .S(\y_c[1].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[1].x_c[0].lc_i.i0muxb  (.A0(\y_c[1].x_c[0].lc_i.i0a ),
    .A1(\y_c[1].x_c[0].lc_i.i0b ),
    .S(\y_c[1].x_c[0].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[1].x_c[0].lc_i.i1muxa0  (.A(\y_c[1].x_c[0].lc_i.cfg[2] ),
    .B(\y_c[0].x_c[2].lc_i.T ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[1].x_c[0].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[0].lc_i.i1muxa1  (.A0(\y_c[1].x_c[0].lc_i.B ),
    .A1(net41),
    .S(\y_c[1].x_c[0].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[0].lc_i.i1muxb  (.A0(\y_c[1].x_c[0].lc_i.i1a ),
    .A1(\y_c[1].x_c[0].lc_i.i1b ),
    .S(\y_c[1].x_c[0].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[1].x_c[0].lc_i.lmux  (.A0(\y_c[1].x_c[0].lc_i.i0 ),
    .A1(\y_c[1].x_c[0].lc_i.i1 ),
    .S(\y_c[1].x_c[0].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[1].x_c[0].lc_i.s0muxa0  (.A(\y_c[0].x_c[0].lc_i.Q ),
    .B(\y_c[1].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[0].lc_i.s0muxa1  (.A0(net42),
    .A1(\y_c[0].x_c[2].lc_i.T ),
    .S(\y_c[1].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[1].x_c[0].lc_i.s0muxb  (.A0(\y_c[1].x_c[0].lc_i.s0a ),
    .A1(\y_c[1].x_c[0].lc_i.s0b ),
    .S(\y_c[1].x_c[0].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[1].x_c[0].lc_i.sinv  (.A(\y_c[1].x_c[0].lc_i.s0s ),
    .B(\y_c[1].x_c[0].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_2 \y_c[1].x_c[1].lc_i.dff.dff  (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(\y_c[1].x_c[1].lc_i.muxo_n ),
    .SET_B(net143),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[1].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[1].x_c[1].lc_i.dff.ffsel  (.A0(\y_c[1].x_c[1].lc_i.muxo_n ),
    .A1(\y_c[1].x_c[1].lc_i.dff.dffo_n ),
    .S(\y_c[1].x_c[1].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[1].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[1].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net197),
    .GATE_N(net107),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[1].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[1].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net194),
    .GATE_N(net108),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[1].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[1].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net189),
    .GATE_N(net107),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[1].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[1].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net186),
    .GATE_N(\y_c[1].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[1].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[1].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net197),
    .GATE_N(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[1].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[1].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net194),
    .GATE_N(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[1].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[1].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net189),
    .GATE_N(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[1].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[1].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net185),
    .GATE_N(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[1].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[1].x_c[1].lc_i.i0muxa0  (.A(net59),
    .B(\y_c[1].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[1].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[1].lc_i.i0muxa1  (.A0(net43),
    .A1(net40),
    .S(\y_c[1].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[1].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[1].lc_i.i0muxb  (.A0(\y_c[1].x_c[1].lc_i.i0a ),
    .A1(\y_c[1].x_c[1].lc_i.i0b ),
    .S(\y_c[1].x_c[1].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[1].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[1].x_c[1].lc_i.i1muxa0  (.A(\y_c[1].x_c[1].lc_i.cfg[2] ),
    .B(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[1].x_c[1].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[1].lc_i.i1muxa1  (.A0(net37),
    .A1(net43),
    .S(\y_c[1].x_c[1].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[1].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[1].lc_i.i1muxb  (.A0(\y_c[1].x_c[1].lc_i.i1a ),
    .A1(\y_c[1].x_c[1].lc_i.i1b ),
    .S(\y_c[1].x_c[1].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[1].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[1].x_c[1].lc_i.lmux  (.A0(\y_c[1].x_c[1].lc_i.i0 ),
    .A1(\y_c[1].x_c[1].lc_i.i1 ),
    .S(\y_c[1].x_c[1].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[1].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[1].x_c[1].lc_i.s0muxa0  (.A(net60),
    .B(\y_c[1].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[1].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_2 \y_c[1].x_c[1].lc_i.s0muxa1  (.A0(net43),
    .A1(\y_c[0].x_c[0].lc_i.B ),
    .S(\y_c[1].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[1].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[1].x_c[1].lc_i.s0muxb  (.A0(\y_c[1].x_c[1].lc_i.s0a ),
    .A1(\y_c[1].x_c[1].lc_i.s0b ),
    .S(\y_c[1].x_c[1].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[1].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[1].x_c[1].lc_i.sinv  (.A(\y_c[1].x_c[1].lc_i.s0s ),
    .B(\y_c[1].x_c[1].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[1].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[1].x_c[2].lc_i.dff.dff  (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(\y_c[1].x_c[2].lc_i.muxo_n ),
    .SET_B(net144),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[2].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_2 \y_c[1].x_c[2].lc_i.dff.ffsel  (.A0(\y_c[1].x_c[2].lc_i.muxo_n ),
    .A1(\y_c[1].x_c[2].lc_i.dff.dffo_n ),
    .S(\y_c[1].x_c[2].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[2].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[2].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net184),
    .GATE_N(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[2].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[2].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net180),
    .GATE_N(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[2].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[2].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net177),
    .GATE_N(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[2].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[2].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net173),
    .GATE_N(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[2].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[2].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net184),
    .GATE_N(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[2].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[2].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net180),
    .GATE_N(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[2].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[2].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(\y_c[0].x_c[2].lc_i.cfg_data[2] ),
    .GATE_N(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[2].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[2].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net174),
    .GATE_N(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[2].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[1].x_c[2].lc_i.i0muxa0  (.A(net57),
    .B(\y_c[1].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[2].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[2].lc_i.i0muxa1  (.A0(net45),
    .A1(\y_c[0].x_c[1].lc_i.B ),
    .S(\y_c[1].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[2].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[2].lc_i.i0muxb  (.A0(\y_c[1].x_c[2].lc_i.i0a ),
    .A1(\y_c[1].x_c[2].lc_i.i0b ),
    .S(\y_c[1].x_c[2].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[2].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[1].x_c[2].lc_i.i1muxa0  (.A(\y_c[1].x_c[2].lc_i.cfg[2] ),
    .B(\y_c[0].x_c[1].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[1].x_c[2].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[2].lc_i.i1muxa1  (.A0(net35),
    .A1(net45),
    .S(\y_c[1].x_c[2].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[2].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[2].lc_i.i1muxb  (.A0(\y_c[1].x_c[2].lc_i.i1a ),
    .A1(\y_c[1].x_c[2].lc_i.i1b ),
    .S(\y_c[1].x_c[2].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[2].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[1].x_c[2].lc_i.lmux  (.A0(\y_c[1].x_c[2].lc_i.i0 ),
    .A1(\y_c[1].x_c[2].lc_i.i1 ),
    .S(\y_c[1].x_c[2].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[2].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[1].x_c[2].lc_i.s0muxa0  (.A(net57),
    .B(\y_c[1].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[2].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[2].lc_i.s0muxa1  (.A0(net45),
    .A1(\y_c[0].x_c[1].lc_i.B ),
    .S(\y_c[1].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[2].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[1].x_c[2].lc_i.s0muxb  (.A0(\y_c[1].x_c[2].lc_i.s0a ),
    .A1(\y_c[1].x_c[2].lc_i.s0b ),
    .S(\y_c[1].x_c[2].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[2].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[1].x_c[2].lc_i.sinv  (.A(\y_c[1].x_c[2].lc_i.s0s ),
    .B(\y_c[1].x_c[2].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[2].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[1].x_c[3].lc_i.dff.dff  (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(\y_c[1].x_c[3].lc_i.muxo_n ),
    .SET_B(_12_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[3].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[3].lc_i.dff.ffsel  (.A0(\y_c[1].x_c[3].lc_i.muxo_n ),
    .A1(\y_c[1].x_c[3].lc_i.dff.dffo_n ),
    .S(\y_c[1].x_c[3].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[3].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[3].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net170),
    .GATE_N(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[3].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[3].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net168),
    .GATE_N(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[3].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[3].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net166),
    .GATE_N(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[3].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[3].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net162),
    .GATE_N(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[3].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[3].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net170),
    .GATE_N(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[3].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[3].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net168),
    .GATE_N(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[3].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[3].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net166),
    .GATE_N(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[3].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[3].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(\y_c[0].x_c[3].lc_i.cfg_data[3] ),
    .GATE_N(\y_c[1].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[3].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[1].x_c[3].lc_i.i0muxa0  (.A(net55),
    .B(\y_c[1].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[3].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[3].lc_i.i0muxa1  (.A0(\y_c[0].x_c[4].lc_i.B ),
    .A1(net44),
    .S(\y_c[1].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[3].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[3].lc_i.i0muxb  (.A0(\y_c[1].x_c[3].lc_i.i0a ),
    .A1(\y_c[1].x_c[3].lc_i.i0b ),
    .S(\y_c[1].x_c[3].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[3].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[1].x_c[3].lc_i.i1muxa0  (.A(\y_c[1].x_c[3].lc_i.cfg[2] ),
    .B(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[1].x_c[3].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_2 \y_c[1].x_c[3].lc_i.i1muxa1  (.A0(\y_c[1].x_c[3].lc_i.B ),
    .A1(\y_c[0].x_c[4].lc_i.B ),
    .S(\y_c[1].x_c[3].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[3].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_4 \y_c[1].x_c[3].lc_i.i1muxb  (.A0(\y_c[1].x_c[3].lc_i.i1a ),
    .A1(\y_c[1].x_c[3].lc_i.i1b ),
    .S(\y_c[1].x_c[3].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[3].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[1].x_c[3].lc_i.lmux  (.A0(\y_c[1].x_c[3].lc_i.i0 ),
    .A1(\y_c[1].x_c[3].lc_i.i1 ),
    .S(\y_c[1].x_c[3].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[3].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[1].x_c[3].lc_i.s0muxa0  (.A(net55),
    .B(\y_c[1].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[3].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[3].lc_i.s0muxa1  (.A0(net52),
    .A1(net44),
    .S(\y_c[1].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[3].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[3].lc_i.s0muxb  (.A0(\y_c[1].x_c[3].lc_i.s0a ),
    .A1(\y_c[1].x_c[3].lc_i.s0b ),
    .S(\y_c[1].x_c[3].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[3].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[1].x_c[3].lc_i.sinv  (.A(\y_c[1].x_c[3].lc_i.s0s ),
    .B(\y_c[1].x_c[3].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[3].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[1].x_c[4].lc_i.dff.dff  (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(\y_c[1].x_c[4].lc_i.muxo_n ),
    .SET_B(net144),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[4].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[1].x_c[4].lc_i.dff.ffsel  (.A0(\y_c[1].x_c[4].lc_i.muxo_n ),
    .A1(\y_c[1].x_c[4].lc_i.dff.dffo_n ),
    .S(\y_c[1].x_c[4].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[0].x_c[4].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[4].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net157),
    .GATE_N(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[4].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[4].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net154),
    .GATE_N(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[4].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[4].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net150),
    .GATE_N(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[4].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[4].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net148),
    .GATE_N(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[4].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[4].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net157),
    .GATE_N(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[4].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[4].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net154),
    .GATE_N(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[4].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[4].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net150),
    .GATE_N(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[4].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[1].x_c[4].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net146),
    .GATE_N(\y_c[1].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[1].x_c[4].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[1].x_c[4].lc_i.i0muxa0  (.A(net53),
    .B(\y_c[1].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[4].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[4].lc_i.i0muxa1  (.A0(net52),
    .A1(\y_c[0].x_c[3].lc_i.B ),
    .S(\y_c[1].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[4].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[4].lc_i.i0muxb  (.A0(\y_c[1].x_c[4].lc_i.i0a ),
    .A1(\y_c[1].x_c[4].lc_i.i0b ),
    .S(\y_c[1].x_c[4].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[4].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[1].x_c[4].lc_i.i1muxa0  (.A(\y_c[1].x_c[4].lc_i.cfg[2] ),
    .B(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[1].x_c[4].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[4].lc_i.i1muxa1  (.A0(\y_c[1].x_c[4].lc_i.B ),
    .A1(net51),
    .S(\y_c[1].x_c[4].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[4].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[4].lc_i.i1muxb  (.A0(\y_c[1].x_c[4].lc_i.i1a ),
    .A1(\y_c[1].x_c[4].lc_i.i1b ),
    .S(\y_c[1].x_c[4].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[4].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[1].x_c[4].lc_i.lmux  (.A0(\y_c[1].x_c[4].lc_i.i0 ),
    .A1(\y_c[1].x_c[4].lc_i.i1 ),
    .S(\y_c[1].x_c[4].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[4].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[1].x_c[4].lc_i.s0muxa0  (.A(net53),
    .B(\y_c[1].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[4].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[1].x_c[4].lc_i.s0muxa1  (.A0(net51),
    .A1(net46),
    .S(\y_c[1].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[4].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[1].x_c[4].lc_i.s0muxb  (.A0(\y_c[1].x_c[4].lc_i.s0a ),
    .A1(\y_c[1].x_c[4].lc_i.s0b ),
    .S(\y_c[1].x_c[4].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[4].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[1].x_c[4].lc_i.sinv  (.A(\y_c[1].x_c[4].lc_i.s0s ),
    .B(\y_c[1].x_c[4].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[4].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[2].x_c[0].lc_i.dff.dff  (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(\y_c[2].x_c[0].lc_i.muxo_n ),
    .SET_B(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[0].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_2 \y_c[2].x_c[0].lc_i.dff.ffsel  (.A0(\y_c[2].x_c[0].lc_i.muxo_n ),
    .A1(\y_c[2].x_c[0].lc_i.dff.dffo_n ),
    .S(\y_c[2].x_c[0].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[0].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[0].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net208),
    .GATE_N(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[0].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[0].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net206),
    .GATE_N(\y_c[2].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[0].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[0].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net203),
    .GATE_N(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[0].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[0].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(\y_c[0].x_c[0].lc_i.cfg_data[3] ),
    .GATE_N(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[0].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[0].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net209),
    .GATE_N(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[0].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[0].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net206),
    .GATE_N(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[0].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[0].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net203),
    .GATE_N(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[0].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[0].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net199),
    .GATE_N(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[0].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[2].x_c[0].lc_i.i0muxa0  (.A(net40),
    .B(\y_c[2].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[0].lc_i.i0muxa1  (.A0(net37),
    .A1(\y_c[0].x_c[3].lc_i.T ),
    .S(\y_c[2].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[2].x_c[0].lc_i.i0muxb  (.A0(\y_c[2].x_c[0].lc_i.i0a ),
    .A1(\y_c[2].x_c[0].lc_i.i0b ),
    .S(\y_c[2].x_c[0].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[2].x_c[0].lc_i.i1muxa0  (.A(\y_c[2].x_c[0].lc_i.cfg[2] ),
    .B(\y_c[0].x_c[3].lc_i.T ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[2].x_c[0].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[0].lc_i.i1muxa1  (.A0(\y_c[2].x_c[0].lc_i.B ),
    .A1(net37),
    .S(\y_c[2].x_c[0].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[0].lc_i.i1muxb  (.A0(\y_c[2].x_c[0].lc_i.i1a ),
    .A1(\y_c[2].x_c[0].lc_i.i1b ),
    .S(\y_c[2].x_c[0].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[2].x_c[0].lc_i.lmux  (.A0(\y_c[2].x_c[0].lc_i.i0 ),
    .A1(\y_c[2].x_c[0].lc_i.i1 ),
    .S(\y_c[2].x_c[0].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[2].x_c[0].lc_i.s0muxa0  (.A(\y_c[0].x_c[0].lc_i.B ),
    .B(\y_c[2].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[0].lc_i.s0muxa1  (.A0(\y_c[1].x_c[1].lc_i.B ),
    .A1(\y_c[0].x_c[3].lc_i.T ),
    .S(\y_c[2].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[0].lc_i.s0muxb  (.A0(\y_c[2].x_c[0].lc_i.s0a ),
    .A1(\y_c[2].x_c[0].lc_i.s0b ),
    .S(\y_c[2].x_c[0].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[2].x_c[0].lc_i.sinv  (.A(\y_c[2].x_c[0].lc_i.s0s ),
    .B(\y_c[2].x_c[0].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_2 \y_c[2].x_c[1].lc_i.dff.dff  (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(\y_c[2].x_c[1].lc_i.muxo_n ),
    .SET_B(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[1].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[2].x_c[1].lc_i.dff.ffsel  (.A0(\y_c[2].x_c[1].lc_i.muxo_n ),
    .A1(\y_c[2].x_c[1].lc_i.dff.dffo_n ),
    .S(\y_c[2].x_c[1].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[1].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[1].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net198),
    .GATE_N(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[1].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[1].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(\y_c[0].x_c[1].lc_i.cfg_data[1] ),
    .GATE_N(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[1].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[1].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net192),
    .GATE_N(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[1].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[1].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net187),
    .GATE_N(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[1].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[1].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net198),
    .GATE_N(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[1].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[1].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(\y_c[0].x_c[1].lc_i.cfg_data[1] ),
    .GATE_N(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[1].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[1].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net190),
    .GATE_N(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[1].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[1].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net185),
    .GATE_N(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[1].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[2].x_c[1].lc_i.i0muxa0  (.A(net41),
    .B(\y_c[2].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[1].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[1].lc_i.i0muxa1  (.A0(net35),
    .A1(\y_c[1].x_c[0].lc_i.B ),
    .S(\y_c[2].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[1].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[2].x_c[1].lc_i.i0muxb  (.A0(\y_c[2].x_c[1].lc_i.i0a ),
    .A1(\y_c[2].x_c[1].lc_i.i0b ),
    .S(\y_c[2].x_c[1].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[1].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[2].x_c[1].lc_i.i1muxa0  (.A(\y_c[2].x_c[1].lc_i.cfg[2] ),
    .B(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[2].x_c[1].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[1].lc_i.i1muxa1  (.A0(\y_c[2].x_c[1].lc_i.B ),
    .A1(net35),
    .S(\y_c[2].x_c[1].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[1].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[1].lc_i.i1muxb  (.A0(\y_c[2].x_c[1].lc_i.i1a ),
    .A1(\y_c[2].x_c[1].lc_i.i1b ),
    .S(\y_c[2].x_c[1].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[1].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[2].x_c[1].lc_i.lmux  (.A0(\y_c[2].x_c[1].lc_i.i0 ),
    .A1(\y_c[2].x_c[1].lc_i.i1 ),
    .S(\y_c[2].x_c[1].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[1].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[2].x_c[1].lc_i.s0muxa0  (.A(net42),
    .B(\y_c[2].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[1].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[1].lc_i.s0muxa1  (.A0(net35),
    .A1(net39),
    .S(\y_c[2].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[1].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[1].lc_i.s0muxb  (.A0(\y_c[2].x_c[1].lc_i.s0a ),
    .A1(\y_c[2].x_c[1].lc_i.s0b ),
    .S(\y_c[2].x_c[1].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[1].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[2].x_c[1].lc_i.sinv  (.A(\y_c[2].x_c[1].lc_i.s0s ),
    .B(\y_c[2].x_c[1].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[1].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_2 \y_c[2].x_c[2].lc_i.dff.dff  (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[2].x_c[2].lc_i.muxo_n ),
    .SET_B(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[2].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[2].x_c[2].lc_i.dff.ffsel  (.A0(\y_c[2].x_c[2].lc_i.muxo_n ),
    .A1(\y_c[2].x_c[2].lc_i.dff.dffo_n ),
    .S(\y_c[2].x_c[2].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[2].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[2].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net182),
    .GATE_N(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[2].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[2].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(\y_c[0].x_c[2].lc_i.cfg_data[1] ),
    .GATE_N(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[2].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[2].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net177),
    .GATE_N(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[2].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[2].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net175),
    .GATE_N(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[2].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[2].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net182),
    .GATE_N(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[2].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[2].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net181),
    .GATE_N(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[2].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[2].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net177),
    .GATE_N(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[2].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[2].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net174),
    .GATE_N(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[2].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[2].x_c[2].lc_i.i0muxa0  (.A(\y_c[0].x_c[2].lc_i.B ),
    .B(\y_c[2].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[2].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[2].lc_i.i0muxa1  (.A0(net48),
    .A1(net38),
    .S(\y_c[2].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[2].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[2].x_c[2].lc_i.i0muxb  (.A0(\y_c[2].x_c[2].lc_i.i0a ),
    .A1(\y_c[2].x_c[2].lc_i.i0b ),
    .S(\y_c[2].x_c[2].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[2].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[2].x_c[2].lc_i.i1muxa0  (.A(\y_c[2].x_c[2].lc_i.cfg[2] ),
    .B(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[2].x_c[2].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[2].lc_i.i1muxa1  (.A0(net34),
    .A1(net48),
    .S(\y_c[2].x_c[2].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[2].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[2].lc_i.i1muxb  (.A0(\y_c[2].x_c[2].lc_i.i1a ),
    .A1(\y_c[2].x_c[2].lc_i.i1b ),
    .S(\y_c[2].x_c[2].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[2].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[2].x_c[2].lc_i.lmux  (.A0(\y_c[2].x_c[2].lc_i.i0 ),
    .A1(\y_c[2].x_c[2].lc_i.i1 ),
    .S(\y_c[2].x_c[2].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[2].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[2].x_c[2].lc_i.s0muxa0  (.A(net44),
    .B(\y_c[2].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[2].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[2].lc_i.s0muxa1  (.A0(\y_c[1].x_c[3].lc_i.B ),
    .A1(\y_c[1].x_c[1].lc_i.B ),
    .S(\y_c[2].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[2].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[2].lc_i.s0muxb  (.A0(\y_c[2].x_c[2].lc_i.s0a ),
    .A1(\y_c[2].x_c[2].lc_i.s0b ),
    .S(\y_c[2].x_c[2].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[2].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[2].x_c[2].lc_i.sinv  (.A(\y_c[2].x_c[2].lc_i.s0s ),
    .B(\y_c[2].x_c[2].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[2].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[2].x_c[3].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[2].x_c[3].lc_i.muxo_n ),
    .SET_B(net140),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[3].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[2].x_c[3].lc_i.dff.ffsel  (.A0(\y_c[2].x_c[3].lc_i.muxo_n ),
    .A1(\y_c[2].x_c[3].lc_i.dff.dffo_n ),
    .S(\y_c[2].x_c[3].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[3].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[3].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net171),
    .GATE_N(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[3].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[3].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net168),
    .GATE_N(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[3].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[3].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net164),
    .GATE_N(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[3].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[3].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net160),
    .GATE_N(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[3].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[3].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net171),
    .GATE_N(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[3].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[3].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net168),
    .GATE_N(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[3].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[3].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net164),
    .GATE_N(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[3].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[3].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net161),
    .GATE_N(\y_c[2].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[3].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[2].x_c[3].lc_i.i0muxa0  (.A(net46),
    .B(\y_c[2].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[3].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[3].lc_i.i0muxa1  (.A0(\y_c[1].x_c[4].lc_i.B ),
    .A1(net36),
    .S(\y_c[2].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[3].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[2].x_c[3].lc_i.i0muxb  (.A0(\y_c[2].x_c[3].lc_i.i0a ),
    .A1(\y_c[2].x_c[3].lc_i.i0b ),
    .S(\y_c[2].x_c[3].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[3].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[2].x_c[3].lc_i.i1muxa0  (.A(\y_c[2].x_c[3].lc_i.cfg[2] ),
    .B(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[2].x_c[3].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[3].lc_i.i1muxa1  (.A0(net19),
    .A1(net50),
    .S(\y_c[2].x_c[3].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[3].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[3].lc_i.i1muxb  (.A0(\y_c[2].x_c[3].lc_i.i1a ),
    .A1(\y_c[2].x_c[3].lc_i.i1b ),
    .S(\y_c[2].x_c[3].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[3].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[2].x_c[3].lc_i.lmux  (.A0(\y_c[2].x_c[3].lc_i.i0 ),
    .A1(\y_c[2].x_c[3].lc_i.i1 ),
    .S(\y_c[2].x_c[3].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[3].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[2].x_c[3].lc_i.s0muxa0  (.A(net46),
    .B(\y_c[2].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[3].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[3].lc_i.s0muxa1  (.A0(net50),
    .A1(net36),
    .S(\y_c[2].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[3].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[3].lc_i.s0muxb  (.A0(\y_c[2].x_c[3].lc_i.s0a ),
    .A1(\y_c[2].x_c[3].lc_i.s0b ),
    .S(\y_c[2].x_c[3].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[3].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[2].x_c[3].lc_i.sinv  (.A(\y_c[2].x_c[3].lc_i.s0s ),
    .B(\y_c[2].x_c[3].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[3].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_2 \y_c[2].x_c[4].lc_i.dff.dff  (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(\y_c[2].x_c[4].lc_i.muxo_n ),
    .SET_B(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[4].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[2].x_c[4].lc_i.dff.ffsel  (.A0(\y_c[2].x_c[4].lc_i.muxo_n ),
    .A1(\y_c[2].x_c[4].lc_i.dff.dffo_n ),
    .S(\y_c[2].x_c[4].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[1].x_c[4].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[4].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net158),
    .GATE_N(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[4].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[4].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net155),
    .GATE_N(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[4].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[4].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net151),
    .GATE_N(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[4].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[4].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net148),
    .GATE_N(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[4].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[4].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net158),
    .GATE_N(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[4].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[4].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net155),
    .GATE_N(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[4].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[2].x_c[4].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net151),
    .GATE_N(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[4].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_2 \y_c[2].x_c[4].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net149),
    .GATE_N(\y_c[2].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[2].x_c[4].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[2].x_c[4].lc_i.i0muxa0  (.A(net51),
    .B(\y_c[2].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[4].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[4].lc_i.i0muxa1  (.A0(net50),
    .A1(net47),
    .S(\y_c[2].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[4].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[2].x_c[4].lc_i.i0muxb  (.A0(\y_c[2].x_c[4].lc_i.i0a ),
    .A1(\y_c[2].x_c[4].lc_i.i0b ),
    .S(\y_c[2].x_c[4].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[4].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[2].x_c[4].lc_i.i1muxa0  (.A(\y_c[2].x_c[4].lc_i.cfg[2] ),
    .B(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[2].x_c[4].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[4].lc_i.i1muxa1  (.A0(net14),
    .A1(net49),
    .S(\y_c[2].x_c[4].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[4].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[4].lc_i.i1muxb  (.A0(\y_c[2].x_c[4].lc_i.i1a ),
    .A1(\y_c[2].x_c[4].lc_i.i1b ),
    .S(\y_c[2].x_c[4].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[4].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[2].x_c[4].lc_i.lmux  (.A0(\y_c[2].x_c[4].lc_i.i0 ),
    .A1(\y_c[2].x_c[4].lc_i.i1 ),
    .S(\y_c[2].x_c[4].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[4].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[2].x_c[4].lc_i.s0muxa0  (.A(net51),
    .B(\y_c[2].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[4].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[4].lc_i.s0muxa1  (.A0(net49),
    .A1(net47),
    .S(\y_c[2].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[4].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[2].x_c[4].lc_i.s0muxb  (.A0(\y_c[2].x_c[4].lc_i.s0a ),
    .A1(\y_c[2].x_c[4].lc_i.s0b ),
    .S(\y_c[2].x_c[4].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[4].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[2].x_c[4].lc_i.sinv  (.A(\y_c[2].x_c[4].lc_i.s0s ),
    .B(\y_c[2].x_c[4].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[4].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[3].x_c[0].lc_i.dff.dff  (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(\y_c[3].x_c[0].lc_i.muxo_n ),
    .SET_B(net143),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[0].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_2 \y_c[3].x_c[0].lc_i.dff.ffsel  (.A0(\y_c[3].x_c[0].lc_i.muxo_n ),
    .A1(\y_c[3].x_c[0].lc_i.dff.dffo_n ),
    .S(\y_c[3].x_c[0].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[0].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[0].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net210),
    .GATE_N(\y_c[3].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[0].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[0].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net206),
    .GATE_N(\y_c[3].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[0].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[0].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net202),
    .GATE_N(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[0].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[0].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net201),
    .GATE_N(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[0].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[0].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net210),
    .GATE_N(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[0].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[0].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net207),
    .GATE_N(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[0].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[0].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net203),
    .GATE_N(\y_c[3].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[0].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[0].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net199),
    .GATE_N(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[0].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[3].x_c[0].lc_i.i0muxa0  (.A(net39),
    .B(\y_c[3].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[0].lc_i.i0muxa1  (.A0(net32),
    .A1(\y_c[0].x_c[4].lc_i.T ),
    .S(\y_c[3].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[3].x_c[0].lc_i.i0muxb  (.A0(\y_c[3].x_c[0].lc_i.i0a ),
    .A1(\y_c[3].x_c[0].lc_i.i0b ),
    .S(\y_c[3].x_c[0].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[3].x_c[0].lc_i.i1muxa0  (.A(\y_c[3].x_c[0].lc_i.cfg[2] ),
    .B(\y_c[0].x_c[4].lc_i.T ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[3].x_c[0].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[0].lc_i.i1muxa1  (.A0(\y_c[3].x_c[0].lc_i.B ),
    .A1(net32),
    .S(\y_c[3].x_c[0].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[3].x_c[0].lc_i.i1muxb  (.A0(\y_c[3].x_c[0].lc_i.i1a ),
    .A1(\y_c[3].x_c[0].lc_i.i1b ),
    .S(\y_c[3].x_c[0].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[3].x_c[0].lc_i.lmux  (.A0(\y_c[3].x_c[0].lc_i.i0 ),
    .A1(\y_c[3].x_c[0].lc_i.i1 ),
    .S(\y_c[3].x_c[0].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[3].x_c[0].lc_i.s0muxa0  (.A(net39),
    .B(\y_c[3].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_2 \y_c[3].x_c[0].lc_i.s0muxa1  (.A0(\y_c[2].x_c[1].lc_i.B ),
    .A1(\y_c[0].x_c[4].lc_i.T ),
    .S(\y_c[3].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_4 \y_c[3].x_c[0].lc_i.s0muxb  (.A0(\y_c[3].x_c[0].lc_i.s0a ),
    .A1(\y_c[3].x_c[0].lc_i.s0b ),
    .S(\y_c[3].x_c[0].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[3].x_c[0].lc_i.sinv  (.A(\y_c[3].x_c[0].lc_i.s0s ),
    .B(\y_c[3].x_c[0].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[3].x_c[1].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[3].x_c[1].lc_i.muxo_n ),
    .SET_B(net141),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[1].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[3].x_c[1].lc_i.dff.ffsel  (.A0(\y_c[3].x_c[1].lc_i.muxo_n ),
    .A1(\y_c[3].x_c[1].lc_i.dff.dffo_n ),
    .S(\y_c[3].x_c[1].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[1].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[1].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net196),
    .GATE_N(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[1].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[1].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net193),
    .GATE_N(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[1].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[1].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net190),
    .GATE_N(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[1].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[1].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net187),
    .GATE_N(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[1].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[1].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net196),
    .GATE_N(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[1].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[1].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net193),
    .GATE_N(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[1].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[1].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net192),
    .GATE_N(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[1].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[1].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net185),
    .GATE_N(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[1].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[3].x_c[1].lc_i.i0muxa0  (.A(net37),
    .B(\y_c[3].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[1].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[1].lc_i.i0muxa1  (.A0(\y_c[2].x_c[2].lc_i.B ),
    .A1(net30),
    .S(\y_c[3].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[1].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[3].x_c[1].lc_i.i0muxb  (.A0(\y_c[3].x_c[1].lc_i.i0a ),
    .A1(\y_c[3].x_c[1].lc_i.i0b ),
    .S(\y_c[3].x_c[1].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[1].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[3].x_c[1].lc_i.i1muxa0  (.A(\y_c[3].x_c[1].lc_i.cfg[2] ),
    .B(\y_c[2].x_c[0].lc_i.B ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[3].x_c[1].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[1].lc_i.i1muxa1  (.A0(\y_c[3].x_c[1].lc_i.B ),
    .A1(\y_c[2].x_c[2].lc_i.B ),
    .S(\y_c[3].x_c[1].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[1].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[1].lc_i.i1muxb  (.A0(\y_c[3].x_c[1].lc_i.i1a ),
    .A1(\y_c[3].x_c[1].lc_i.i1b ),
    .S(\y_c[3].x_c[1].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[1].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[3].x_c[1].lc_i.lmux  (.A0(\y_c[3].x_c[1].lc_i.i0 ),
    .A1(\y_c[3].x_c[1].lc_i.i1 ),
    .S(\y_c[3].x_c[1].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[1].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[3].x_c[1].lc_i.s0muxa0  (.A(net38),
    .B(\y_c[3].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[1].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[1].lc_i.s0muxa1  (.A0(net34),
    .A1(net30),
    .S(\y_c[3].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[1].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[3].x_c[1].lc_i.s0muxb  (.A0(\y_c[3].x_c[1].lc_i.s0a ),
    .A1(\y_c[3].x_c[1].lc_i.s0b ),
    .S(\y_c[3].x_c[1].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[1].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[3].x_c[1].lc_i.sinv  (.A(\y_c[3].x_c[1].lc_i.s0s ),
    .B(\y_c[3].x_c[1].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[1].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[3].x_c[2].lc_i.dff.dff  (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(\y_c[3].x_c[2].lc_i.muxo_n ),
    .SET_B(_12_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[2].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[3].x_c[2].lc_i.dff.ffsel  (.A0(\y_c[3].x_c[2].lc_i.muxo_n ),
    .A1(\y_c[3].x_c[2].lc_i.dff.dffo_n ),
    .S(\y_c[3].x_c[2].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[2].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[2].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net182),
    .GATE_N(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[2].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[2].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net181),
    .GATE_N(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[2].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[2].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net176),
    .GATE_N(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[2].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[2].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net174),
    .GATE_N(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[2].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[2].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net182),
    .GATE_N(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[2].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[2].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net181),
    .GATE_N(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[2].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[2].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net176),
    .GATE_N(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[2].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[2].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net173),
    .GATE_N(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[2].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[3].x_c[2].lc_i.i0muxa0  (.A(\y_c[1].x_c[2].lc_i.B ),
    .B(\y_c[3].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[2].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[2].lc_i.i0muxa1  (.A0(net19),
    .A1(net31),
    .S(\y_c[3].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[2].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[2].lc_i.i0muxb  (.A0(\y_c[3].x_c[2].lc_i.i0a ),
    .A1(\y_c[3].x_c[2].lc_i.i0b ),
    .S(\y_c[3].x_c[2].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[2].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[3].x_c[2].lc_i.i1muxa0  (.A(\y_c[3].x_c[2].lc_i.cfg[2] ),
    .B(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[3].x_c[2].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[2].lc_i.i1muxa1  (.A0(\y_c[3].x_c[2].lc_i.B ),
    .A1(\y_c[2].x_c[3].lc_i.B ),
    .S(\y_c[3].x_c[2].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[2].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[2].lc_i.i1muxb  (.A0(\y_c[3].x_c[2].lc_i.i1a ),
    .A1(\y_c[3].x_c[2].lc_i.i1b ),
    .S(\y_c[3].x_c[2].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[2].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[3].x_c[2].lc_i.lmux  (.A0(\y_c[3].x_c[2].lc_i.i0 ),
    .A1(\y_c[3].x_c[2].lc_i.i1 ),
    .S(\y_c[3].x_c[2].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[2].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[3].x_c[2].lc_i.s0muxa0  (.A(\y_c[1].x_c[2].lc_i.B ),
    .B(\y_c[3].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[2].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[2].lc_i.s0muxa1  (.A0(\y_c[2].x_c[3].lc_i.B ),
    .A1(net31),
    .S(\y_c[3].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[2].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[3].x_c[2].lc_i.s0muxb  (.A0(\y_c[3].x_c[2].lc_i.s0a ),
    .A1(\y_c[3].x_c[2].lc_i.s0b ),
    .S(\y_c[3].x_c[2].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[2].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[3].x_c[2].lc_i.sinv  (.A(\y_c[3].x_c[2].lc_i.s0s ),
    .B(\y_c[3].x_c[2].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[2].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[3].x_c[3].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[3].x_c[3].lc_i.muxo_n ),
    .SET_B(net140),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[3].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[3].x_c[3].lc_i.dff.ffsel  (.A0(\y_c[3].x_c[3].lc_i.muxo_n ),
    .A1(\y_c[3].x_c[3].lc_i.dff.dffo_n ),
    .S(\y_c[3].x_c[3].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[3].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[3].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net172),
    .GATE_N(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[3].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[3].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net167),
    .GATE_N(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[3].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[3].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net164),
    .GATE_N(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[3].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[3].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net160),
    .GATE_N(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[3].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[3].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net171),
    .GATE_N(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[3].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[3].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net167),
    .GATE_N(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[3].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[3].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net164),
    .GATE_N(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[3].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[3].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net162),
    .GATE_N(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[3].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[3].x_c[3].lc_i.i0muxa0  (.A(net48),
    .B(\y_c[3].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[3].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[3].lc_i.i0muxa1  (.A0(\y_c[2].x_c[4].lc_i.B ),
    .A1(net33),
    .S(\y_c[3].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[3].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[3].lc_i.i0muxb  (.A0(\y_c[3].x_c[3].lc_i.i0a ),
    .A1(\y_c[3].x_c[3].lc_i.i0b ),
    .S(\y_c[3].x_c[3].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[3].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[3].x_c[3].lc_i.i1muxa0  (.A(\y_c[3].x_c[3].lc_i.cfg[2] ),
    .B(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[3].x_c[3].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[3].lc_i.i1muxa1  (.A0(\y_c[3].x_c[3].lc_i.B ),
    .A1(\y_c[2].x_c[4].lc_i.B ),
    .S(\y_c[3].x_c[3].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[3].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[3].x_c[3].lc_i.i1muxb  (.A0(\y_c[3].x_c[3].lc_i.i1a ),
    .A1(\y_c[3].x_c[3].lc_i.i1b ),
    .S(\y_c[3].x_c[3].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[3].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[3].x_c[3].lc_i.lmux  (.A0(\y_c[3].x_c[3].lc_i.i0 ),
    .A1(\y_c[3].x_c[3].lc_i.i1 ),
    .S(\y_c[3].x_c[3].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[3].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[3].x_c[3].lc_i.s0muxa0  (.A(net47),
    .B(\y_c[3].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[3].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[3].lc_i.s0muxa1  (.A0(\y_c[2].x_c[4].lc_i.B ),
    .A1(net33),
    .S(\y_c[3].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[3].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[3].x_c[3].lc_i.s0muxb  (.A0(\y_c[3].x_c[3].lc_i.s0a ),
    .A1(\y_c[3].x_c[3].lc_i.s0b ),
    .S(\y_c[3].x_c[3].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[3].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[3].x_c[3].lc_i.sinv  (.A(\y_c[3].x_c[3].lc_i.s0s ),
    .B(\y_c[3].x_c[3].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[3].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[3].x_c[4].lc_i.dff.dff  (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[3].x_c[4].lc_i.muxo_n ),
    .SET_B(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[4].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[3].x_c[4].lc_i.dff.ffsel  (.A0(\y_c[3].x_c[4].lc_i.muxo_n ),
    .A1(\y_c[3].x_c[4].lc_i.dff.dffo_n ),
    .S(\y_c[3].x_c[4].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[2].x_c[4].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[4].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net159),
    .GATE_N(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[4].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[4].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net156),
    .GATE_N(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[4].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[4].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net152),
    .GATE_N(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[4].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[4].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net148),
    .GATE_N(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[4].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[4].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net158),
    .GATE_N(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[4].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[4].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net155),
    .GATE_N(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[4].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[4].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net151),
    .GATE_N(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[4].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[3].x_c[4].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net146),
    .GATE_N(\y_c[3].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[3].x_c[4].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[3].x_c[4].lc_i.i0muxa0  (.A(net49),
    .B(\y_c[3].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[4].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[4].lc_i.i0muxa1  (.A0(net14),
    .A1(net18),
    .S(\y_c[3].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[4].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[4].lc_i.i0muxb  (.A0(\y_c[3].x_c[4].lc_i.i0a ),
    .A1(\y_c[3].x_c[4].lc_i.i0b ),
    .S(\y_c[3].x_c[4].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[4].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[3].x_c[4].lc_i.i1muxa0  (.A(\y_c[3].x_c[4].lc_i.cfg[2] ),
    .B(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[3].x_c[4].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[4].lc_i.i1muxa1  (.A0(net11),
    .A1(net14),
    .S(\y_c[3].x_c[4].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[4].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[3].x_c[4].lc_i.i1muxb  (.A0(\y_c[3].x_c[4].lc_i.i1a ),
    .A1(\y_c[3].x_c[4].lc_i.i1b ),
    .S(\y_c[3].x_c[4].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[4].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[3].x_c[4].lc_i.lmux  (.A0(\y_c[3].x_c[4].lc_i.i0 ),
    .A1(\y_c[3].x_c[4].lc_i.i1 ),
    .S(\y_c[3].x_c[4].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[4].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[3].x_c[4].lc_i.s0muxa0  (.A(net49),
    .B(\y_c[3].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[4].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[3].x_c[4].lc_i.s0muxa1  (.A0(net14),
    .A1(net18),
    .S(\y_c[3].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[4].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[3].x_c[4].lc_i.s0muxb  (.A0(\y_c[3].x_c[4].lc_i.s0a ),
    .A1(\y_c[3].x_c[4].lc_i.s0b ),
    .S(\y_c[3].x_c[4].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[4].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[3].x_c[4].lc_i.sinv  (.A(\y_c[3].x_c[4].lc_i.s0s ),
    .B(\y_c[3].x_c[4].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[4].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[4].x_c[0].lc_i.dff.dff  (.CLK(clknet_2_3__leaf_io_in[0]),
    .D(\y_c[4].x_c[0].lc_i.muxo_n ),
    .SET_B(net143),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[0].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[0].lc_i.dff.ffsel  (.A0(\y_c[4].x_c[0].lc_i.muxo_n ),
    .A1(\y_c[4].x_c[0].lc_i.dff.dffo_n ),
    .S(\y_c[4].x_c[0].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[0].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[0].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(\y_c[0].x_c[0].lc_i.cfg_data[0] ),
    .GATE_N(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[0].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[0].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net207),
    .GATE_N(\y_c[4].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[0].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[0].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net202),
    .GATE_N(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[0].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[0].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net201),
    .GATE_N(\y_c[4].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[0].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[0].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net210),
    .GATE_N(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[0].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[0].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net207),
    .GATE_N(\y_c[4].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[0].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[0].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net202),
    .GATE_N(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[0].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_2 \y_c[4].x_c[0].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net201),
    .GATE_N(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[0].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[4].x_c[0].lc_i.i0muxa0  (.A(net30),
    .B(\y_c[4].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[0].lc_i.i0muxa1  (.A0(\y_c[3].x_c[1].lc_i.B ),
    .A1(\y_c[4].x_c[0].lc_i.L ),
    .S(\y_c[4].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[0].lc_i.i0muxb  (.A0(\y_c[4].x_c[0].lc_i.i0a ),
    .A1(\y_c[4].x_c[0].lc_i.i0b ),
    .S(\y_c[4].x_c[0].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[4].x_c[0].lc_i.i1muxa0  (.A(\y_c[4].x_c[0].lc_i.cfg[2] ),
    .B(\y_c[4].x_c[0].lc_i.L ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[4].x_c[0].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[0].lc_i.i1muxa1  (.A0(net28),
    .A1(net12),
    .S(\y_c[4].x_c[0].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[0].lc_i.i1muxb  (.A0(\y_c[4].x_c[0].lc_i.i1a ),
    .A1(\y_c[4].x_c[0].lc_i.i1b ),
    .S(\y_c[4].x_c[0].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[0].lc_i.lmux  (.A0(\y_c[4].x_c[0].lc_i.i0 ),
    .A1(\y_c[4].x_c[0].lc_i.i1 ),
    .S(\y_c[4].x_c[0].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[4].x_c[0].lc_i.s0muxa0  (.A(net30),
    .B(\y_c[4].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[0].lc_i.s0muxa1  (.A0(net13),
    .A1(\y_c[4].x_c[0].lc_i.L ),
    .S(\y_c[4].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[4].x_c[0].lc_i.s0muxb  (.A0(\y_c[4].x_c[0].lc_i.s0a ),
    .A1(\y_c[4].x_c[0].lc_i.s0b ),
    .S(\y_c[4].x_c[0].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[4].x_c[0].lc_i.sinv  (.A(\y_c[4].x_c[0].lc_i.s0s ),
    .B(\y_c[4].x_c[0].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[4].x_c[1].lc_i.dff.dff  (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[4].x_c[1].lc_i.muxo_n ),
    .SET_B(net141),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[1].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[1].lc_i.dff.ffsel  (.A0(\y_c[4].x_c[1].lc_i.muxo_n ),
    .A1(\y_c[4].x_c[1].lc_i.dff.dffo_n ),
    .S(\y_c[4].x_c[1].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[1].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[1].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net196),
    .GATE_N(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[1].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[1].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net193),
    .GATE_N(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[1].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[1].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net191),
    .GATE_N(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[1].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[1].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net188),
    .GATE_N(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[1].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[1].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net196),
    .GATE_N(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[1].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[1].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net193),
    .GATE_N(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[1].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[1].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net191),
    .GATE_N(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[1].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[1].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net188),
    .GATE_N(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[1].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[4].x_c[1].lc_i.i0muxa0  (.A(net31),
    .B(\y_c[4].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[1].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[1].lc_i.i0muxa1  (.A0(\y_c[3].x_c[2].lc_i.B ),
    .A1(net29),
    .S(\y_c[4].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[1].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[4].x_c[1].lc_i.i0muxb  (.A0(\y_c[4].x_c[1].lc_i.i0a ),
    .A1(\y_c[4].x_c[1].lc_i.i0b ),
    .S(\y_c[4].x_c[1].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[1].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[4].x_c[1].lc_i.i1muxa0  (.A(\y_c[4].x_c[1].lc_i.cfg[2] ),
    .B(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[4].x_c[1].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_2 \y_c[4].x_c[1].lc_i.i1muxa1  (.A0(net26),
    .A1(net16),
    .S(\y_c[4].x_c[1].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[1].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[1].lc_i.i1muxb  (.A0(\y_c[4].x_c[1].lc_i.i1a ),
    .A1(\y_c[4].x_c[1].lc_i.i1b ),
    .S(\y_c[4].x_c[1].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[1].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[1].lc_i.lmux  (.A0(\y_c[4].x_c[1].lc_i.i0 ),
    .A1(\y_c[4].x_c[1].lc_i.i1 ),
    .S(\y_c[4].x_c[1].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[1].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[4].x_c[1].lc_i.s0muxa0  (.A(net31),
    .B(\y_c[4].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[1].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[1].lc_i.s0muxa1  (.A0(net17),
    .A1(net29),
    .S(\y_c[4].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[1].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[4].x_c[1].lc_i.s0muxb  (.A0(\y_c[4].x_c[1].lc_i.s0a ),
    .A1(\y_c[4].x_c[1].lc_i.s0b ),
    .S(\y_c[4].x_c[1].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[1].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[4].x_c[1].lc_i.sinv  (.A(\y_c[4].x_c[1].lc_i.s0s ),
    .B(\y_c[4].x_c[1].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[1].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[4].x_c[2].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[4].x_c[2].lc_i.muxo_n ),
    .SET_B(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[2].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[2].lc_i.dff.ffsel  (.A0(\y_c[4].x_c[2].lc_i.muxo_n ),
    .A1(\y_c[4].x_c[2].lc_i.dff.dffo_n ),
    .S(\y_c[4].x_c[2].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[2].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[2].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net183),
    .GATE_N(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[2].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[2].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net179),
    .GATE_N(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[2].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[2].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net176),
    .GATE_N(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[2].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[2].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(\y_c[0].x_c[2].lc_i.cfg_data[3] ),
    .GATE_N(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[2].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[2].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net183),
    .GATE_N(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[2].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[2].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net179),
    .GATE_N(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[2].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[2].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net176),
    .GATE_N(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[2].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[2].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net175),
    .GATE_N(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[2].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[4].x_c[2].lc_i.i0muxa0  (.A(net33),
    .B(\y_c[4].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[2].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[2].lc_i.i0muxa1  (.A0(net21),
    .A1(net13),
    .S(\y_c[4].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[2].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[2].lc_i.i0muxb  (.A0(\y_c[4].x_c[2].lc_i.i0a ),
    .A1(\y_c[4].x_c[2].lc_i.i0b ),
    .S(\y_c[4].x_c[2].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[2].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[4].x_c[2].lc_i.i1muxa0  (.A(\y_c[4].x_c[2].lc_i.cfg[2] ),
    .B(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[4].x_c[2].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[2].lc_i.i1muxa1  (.A0(net24),
    .A1(net20),
    .S(\y_c[4].x_c[2].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[2].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[2].lc_i.i1muxb  (.A0(\y_c[4].x_c[2].lc_i.i1a ),
    .A1(\y_c[4].x_c[2].lc_i.i1b ),
    .S(\y_c[4].x_c[2].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[2].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[2].lc_i.lmux  (.A0(\y_c[4].x_c[2].lc_i.i0 ),
    .A1(\y_c[4].x_c[2].lc_i.i1 ),
    .S(\y_c[4].x_c[2].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[2].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[4].x_c[2].lc_i.s0muxa0  (.A(net33),
    .B(\y_c[4].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[2].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[2].lc_i.s0muxa1  (.A0(net21),
    .A1(net12),
    .S(\y_c[4].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[2].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[4].x_c[2].lc_i.s0muxb  (.A0(\y_c[4].x_c[2].lc_i.s0a ),
    .A1(\y_c[4].x_c[2].lc_i.s0b ),
    .S(\y_c[4].x_c[2].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[2].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[4].x_c[2].lc_i.sinv  (.A(\y_c[4].x_c[2].lc_i.s0s ),
    .B(\y_c[4].x_c[2].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[2].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[4].x_c[3].lc_i.dff.dff  (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[4].x_c[3].lc_i.muxo_n ),
    .SET_B(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[3].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[3].lc_i.dff.ffsel  (.A0(\y_c[4].x_c[3].lc_i.muxo_n ),
    .A1(\y_c[4].x_c[3].lc_i.dff.dffo_n ),
    .S(\y_c[4].x_c[3].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[3].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[3].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net172),
    .GATE_N(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[3].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[3].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net167),
    .GATE_N(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[3].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[3].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net165),
    .GATE_N(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[3].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[3].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net160),
    .GATE_N(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[3].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[3].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net172),
    .GATE_N(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[3].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[3].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net167),
    .GATE_N(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[3].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[3].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net165),
    .GATE_N(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[3].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[3].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net161),
    .GATE_N(\y_c[4].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[3].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[4].x_c[3].lc_i.i0muxa0  (.A(net18),
    .B(\y_c[4].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[3].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[3].lc_i.i0muxa1  (.A0(net11),
    .A1(net17),
    .S(\y_c[4].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[3].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[3].lc_i.i0muxb  (.A0(\y_c[4].x_c[3].lc_i.i0a ),
    .A1(\y_c[4].x_c[3].lc_i.i0b ),
    .S(\y_c[4].x_c[3].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[3].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[4].x_c[3].lc_i.i1muxa0  (.A(\y_c[4].x_c[3].lc_i.cfg[2] ),
    .B(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[4].x_c[3].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[3].lc_i.i1muxa1  (.A0(\y_c[4].x_c[3].lc_i.B ),
    .A1(\y_c[3].x_c[4].lc_i.B ),
    .S(\y_c[4].x_c[3].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[3].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[4].x_c[3].lc_i.i1muxb  (.A0(\y_c[4].x_c[3].lc_i.i1a ),
    .A1(\y_c[4].x_c[3].lc_i.i1b ),
    .S(\y_c[4].x_c[3].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[3].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[3].lc_i.lmux  (.A0(\y_c[4].x_c[3].lc_i.i0 ),
    .A1(\y_c[4].x_c[3].lc_i.i1 ),
    .S(\y_c[4].x_c[3].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[3].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[4].x_c[3].lc_i.s0muxa0  (.A(net18),
    .B(\y_c[4].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[3].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[3].lc_i.s0muxa1  (.A0(net11),
    .A1(net17),
    .S(\y_c[4].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[3].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[4].x_c[3].lc_i.s0muxb  (.A0(\y_c[4].x_c[3].lc_i.s0a ),
    .A1(\y_c[4].x_c[3].lc_i.s0b ),
    .S(\y_c[4].x_c[3].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[3].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[4].x_c[3].lc_i.sinv  (.A(\y_c[4].x_c[3].lc_i.s0s ),
    .B(\y_c[4].x_c[3].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[3].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[4].x_c[4].lc_i.dff.dff  (.CLK(clknet_2_2__leaf_io_in[0]),
    .D(\y_c[4].x_c[4].lc_i.muxo_n ),
    .SET_B(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[4].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[4].lc_i.dff.ffsel  (.A0(\y_c[4].x_c[4].lc_i.muxo_n ),
    .A1(\y_c[4].x_c[4].lc_i.dff.dffo_n ),
    .S(\y_c[4].x_c[4].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[3].x_c[4].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[4].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net159),
    .GATE_N(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[4].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[4].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net156),
    .GATE_N(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[4].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[4].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net153),
    .GATE_N(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[4].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[4].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net148),
    .GATE_N(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[4].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[4].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(net159),
    .GATE_N(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[4].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[4].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net156),
    .GATE_N(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[4].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[4].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net152),
    .GATE_N(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[4].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[4].x_c[4].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net147),
    .GATE_N(\y_c[4].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[4].x_c[4].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[4].x_c[4].lc_i.i0muxa0  (.A(net15),
    .B(\y_c[4].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[4].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[4].lc_i.i0muxa1  (.A0(\y_c[3].x_c[4].lc_i.B ),
    .A1(net20),
    .S(\y_c[4].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[4].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[4].lc_i.i0muxb  (.A0(\y_c[4].x_c[4].lc_i.i0a ),
    .A1(\y_c[4].x_c[4].lc_i.i0b ),
    .S(\y_c[4].x_c[4].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[4].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[4].x_c[4].lc_i.i1muxa0  (.A(\y_c[4].x_c[4].lc_i.cfg[2] ),
    .B(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[4].x_c[4].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[4].lc_i.i1muxa1  (.A0(\y_c[4].x_c[4].lc_i.B ),
    .A1(net10),
    .S(\y_c[4].x_c[4].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[4].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[4].lc_i.i1muxb  (.A0(\y_c[4].x_c[4].lc_i.i1a ),
    .A1(\y_c[4].x_c[4].lc_i.i1b ),
    .S(\y_c[4].x_c[4].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[4].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[4].lc_i.lmux  (.A0(\y_c[4].x_c[4].lc_i.i0 ),
    .A1(\y_c[4].x_c[4].lc_i.i1 ),
    .S(\y_c[4].x_c[4].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[4].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[4].x_c[4].lc_i.s0muxa0  (.A(net15),
    .B(\y_c[4].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[4].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[4].x_c[4].lc_i.s0muxa1  (.A0(net11),
    .A1(net21),
    .S(\y_c[4].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[4].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_4 \y_c[4].x_c[4].lc_i.s0muxb  (.A0(\y_c[4].x_c[4].lc_i.s0a ),
    .A1(\y_c[4].x_c[4].lc_i.s0b ),
    .S(\y_c[4].x_c[4].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[4].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[4].x_c[4].lc_i.sinv  (.A(\y_c[4].x_c[4].lc_i.s0s ),
    .B(\y_c[4].x_c[4].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[4].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[5].x_c[0].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[5].x_c[0].lc_i.muxo_n ),
    .SET_B(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[0].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[5].x_c[0].lc_i.dff.ffsel  (.A0(\y_c[5].x_c[0].lc_i.muxo_n ),
    .A1(\y_c[5].x_c[0].lc_i.dff.dffo_n ),
    .S(\y_c[5].x_c[0].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[0].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[0].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(\y_c[0].x_c[0].lc_i.cfg_data[0] ),
    .GATE_N(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[0].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[0].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(\y_c[0].x_c[0].lc_i.cfg_data[1] ),
    .GATE_N(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[0].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[0].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net202),
    .GATE_N(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[0].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[0].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net201),
    .GATE_N(\y_c[5].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[0].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[0].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(\y_c[0].x_c[0].lc_i.cfg_data[0] ),
    .GATE_N(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[0].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[0].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(\y_c[0].x_c[0].lc_i.cfg_data[1] ),
    .GATE_N(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[0].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[0].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(\y_c[0].x_c[0].lc_i.cfg_data[2] ),
    .GATE_N(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[0].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[0].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net199),
    .GATE_N(\y_c[5].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[0].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[5].x_c[0].lc_i.i0muxa0  (.A(\y_c[3].x_c[0].lc_i.B ),
    .B(\y_c[5].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[0].lc_i.i0muxa1  (.A0(net27),
    .A1(\y_c[5].x_c[0].lc_i.L ),
    .S(\y_c[5].x_c[0].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[5].x_c[0].lc_i.i0muxb  (.A0(\y_c[5].x_c[0].lc_i.i0a ),
    .A1(\y_c[5].x_c[0].lc_i.i0b ),
    .S(\y_c[5].x_c[0].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[5].x_c[0].lc_i.i1muxa0  (.A(\y_c[5].x_c[0].lc_i.cfg[2] ),
    .B(\y_c[5].x_c[0].lc_i.L ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[5].x_c[0].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[0].lc_i.i1muxa1  (.A0(net28),
    .A1(net27),
    .S(\y_c[5].x_c[0].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[0].lc_i.i1muxb  (.A0(\y_c[5].x_c[0].lc_i.i1a ),
    .A1(\y_c[5].x_c[0].lc_i.i1b ),
    .S(\y_c[5].x_c[0].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[5].x_c[0].lc_i.lmux  (.A0(\y_c[5].x_c[0].lc_i.i0 ),
    .A1(\y_c[5].x_c[0].lc_i.i1 ),
    .S(\y_c[5].x_c[0].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[5].x_c[0].lc_i.s0muxa0  (.A(net29),
    .B(\y_c[5].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[0].lc_i.s0muxa1  (.A0(\y_c[4].x_c[1].lc_i.B ),
    .A1(\y_c[5].x_c[0].lc_i.L ),
    .S(\y_c[5].x_c[0].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[5].x_c[0].lc_i.s0muxb  (.A0(\y_c[5].x_c[0].lc_i.s0a ),
    .A1(\y_c[5].x_c[0].lc_i.s0b ),
    .S(\y_c[5].x_c[0].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[5].x_c[0].lc_i.sinv  (.A(\y_c[5].x_c[0].lc_i.s0s ),
    .B(\y_c[5].x_c[0].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[0].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[5].x_c[1].lc_i.dff.dff  (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[5].x_c[1].lc_i.muxo_n ),
    .SET_B(net136),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[1].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_2 \y_c[5].x_c[1].lc_i.dff.ffsel  (.A0(\y_c[5].x_c[1].lc_i.muxo_n ),
    .A1(\y_c[5].x_c[1].lc_i.dff.dffo_n ),
    .S(\y_c[5].x_c[1].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[1].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[1].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(\y_c[0].x_c[1].lc_i.cfg_data[0] ),
    .GATE_N(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[1].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[1].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net195),
    .GATE_N(net124),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[1].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[1].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net191),
    .GATE_N(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[1].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[1].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net188),
    .GATE_N(\y_c[5].x_c[0].lc_i.cfg_strb[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[1].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[1].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(\y_c[0].x_c[1].lc_i.cfg_data[0] ),
    .GATE_N(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[1].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[1].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net195),
    .GATE_N(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[1].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[1].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net191),
    .GATE_N(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[1].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[1].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net186),
    .GATE_N(\y_c[5].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[1].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[5].x_c[1].lc_i.i0muxa0  (.A(net13),
    .B(\y_c[5].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[1].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[1].lc_i.i0muxa1  (.A0(net25),
    .A1(net28),
    .S(\y_c[5].x_c[1].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[1].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[1].lc_i.i0muxb  (.A0(\y_c[5].x_c[1].lc_i.i0a ),
    .A1(\y_c[5].x_c[1].lc_i.i0b ),
    .S(\y_c[5].x_c[1].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[1].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[5].x_c[1].lc_i.i1muxa0  (.A(\y_c[5].x_c[1].lc_i.cfg[2] ),
    .B(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[5].x_c[1].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[1].lc_i.i1muxa1  (.A0(net27),
    .A1(\y_c[4].x_c[2].lc_i.B ),
    .S(\y_c[5].x_c[1].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[1].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[1].lc_i.i1muxb  (.A0(\y_c[5].x_c[1].lc_i.i1a ),
    .A1(\y_c[5].x_c[1].lc_i.i1b ),
    .S(\y_c[5].x_c[1].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[1].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[5].x_c[1].lc_i.lmux  (.A0(\y_c[5].x_c[1].lc_i.i0 ),
    .A1(\y_c[5].x_c[1].lc_i.i1 ),
    .S(\y_c[5].x_c[1].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[1].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[5].x_c[1].lc_i.s0muxa0  (.A(net12),
    .B(\y_c[5].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[1].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_2 \y_c[5].x_c[1].lc_i.s0muxa1  (.A0(net25),
    .A1(\y_c[4].x_c[0].lc_i.B ),
    .S(\y_c[5].x_c[1].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[1].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_4 \y_c[5].x_c[1].lc_i.s0muxb  (.A0(\y_c[5].x_c[1].lc_i.s0a ),
    .A1(\y_c[5].x_c[1].lc_i.s0b ),
    .S(\y_c[5].x_c[1].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[1].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[5].x_c[1].lc_i.sinv  (.A(\y_c[5].x_c[1].lc_i.s0s ),
    .B(\y_c[5].x_c[1].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[1].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[5].x_c[2].lc_i.dff.dff  (.CLK(clknet_2_0__leaf_io_in[0]),
    .D(\y_c[5].x_c[2].lc_i.muxo_n ),
    .SET_B(net136),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[2].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[5].x_c[2].lc_i.dff.ffsel  (.A0(\y_c[5].x_c[2].lc_i.muxo_n ),
    .A1(\y_c[5].x_c[2].lc_i.dff.dffo_n ),
    .S(\y_c[5].x_c[2].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[2].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[2].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(net183),
    .GATE_N(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[2].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[2].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net179),
    .GATE_N(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[2].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[2].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net178),
    .GATE_N(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[2].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[2].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(\y_c[0].x_c[2].lc_i.cfg_data[3] ),
    .GATE_N(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[2].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[2].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(\y_c[0].x_c[2].lc_i.cfg_data[0] ),
    .GATE_N(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[2].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[2].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net179),
    .GATE_N(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[2].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[2].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net178),
    .GATE_N(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[2].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[2].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net175),
    .GATE_N(\y_c[5].x_c[0].lc_i.cfg_strb[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[2].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[5].x_c[2].lc_i.i0muxa0  (.A(net16),
    .B(\y_c[5].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[2].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[2].lc_i.i0muxa1  (.A0(net23),
    .A1(net26),
    .S(\y_c[5].x_c[2].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[2].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[2].lc_i.i0muxb  (.A0(\y_c[5].x_c[2].lc_i.i0a ),
    .A1(\y_c[5].x_c[2].lc_i.i0b ),
    .S(\y_c[5].x_c[2].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[2].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[5].x_c[2].lc_i.i1muxa0  (.A(\y_c[5].x_c[2].lc_i.cfg[2] ),
    .B(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[5].x_c[2].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[2].lc_i.i1muxa1  (.A0(\y_c[4].x_c[2].lc_i.B ),
    .A1(\y_c[4].x_c[3].lc_i.B ),
    .S(\y_c[5].x_c[2].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[2].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_4 \y_c[5].x_c[2].lc_i.i1muxb  (.A0(\y_c[5].x_c[2].lc_i.i1a ),
    .A1(\y_c[5].x_c[2].lc_i.i1b ),
    .S(\y_c[5].x_c[2].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[2].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[5].x_c[2].lc_i.lmux  (.A0(\y_c[5].x_c[2].lc_i.i0 ),
    .A1(\y_c[5].x_c[2].lc_i.i1 ),
    .S(\y_c[5].x_c[2].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[2].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[5].x_c[2].lc_i.s0muxa0  (.A(net16),
    .B(\y_c[5].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[2].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[2].lc_i.s0muxa1  (.A0(net22),
    .A1(net26),
    .S(\y_c[5].x_c[2].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[2].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[5].x_c[2].lc_i.s0muxb  (.A0(\y_c[5].x_c[2].lc_i.s0a ),
    .A1(\y_c[5].x_c[2].lc_i.s0b ),
    .S(\y_c[5].x_c[2].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[2].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[5].x_c[2].lc_i.sinv  (.A(\y_c[5].x_c[2].lc_i.s0s ),
    .B(\y_c[5].x_c[2].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[2].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[5].x_c[3].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[5].x_c[3].lc_i.muxo_n ),
    .SET_B(net136),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[3].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_2 \y_c[5].x_c[3].lc_i.dff.ffsel  (.A0(\y_c[5].x_c[3].lc_i.muxo_n ),
    .A1(\y_c[5].x_c[3].lc_i.dff.dffo_n ),
    .S(\y_c[5].x_c[3].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[3].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[3].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(\y_c[0].x_c[3].lc_i.cfg_data[0] ),
    .GATE_N(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[3].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[3].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(net169),
    .GATE_N(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[3].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[3].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(\y_c[0].x_c[3].lc_i.cfg_data[2] ),
    .GATE_N(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[3].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[3].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net160),
    .GATE_N(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[3].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[3].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(\y_c[0].x_c[3].lc_i.cfg_data[0] ),
    .GATE_N(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[3].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[3].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(net169),
    .GATE_N(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[3].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[3].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net165),
    .GATE_N(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[3].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[3].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net161),
    .GATE_N(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[3].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[5].x_c[3].lc_i.i0muxa0  (.A(\y_c[3].x_c[3].lc_i.B ),
    .B(\y_c[5].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[3].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[3].lc_i.i0muxa1  (.A0(net9),
    .A1(net24),
    .S(\y_c[5].x_c[3].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[3].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[3].lc_i.i0muxb  (.A0(\y_c[5].x_c[3].lc_i.i0a ),
    .A1(\y_c[5].x_c[3].lc_i.i0b ),
    .S(\y_c[5].x_c[3].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[3].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[5].x_c[3].lc_i.i1muxa0  (.A(\y_c[5].x_c[3].lc_i.cfg[2] ),
    .B(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[5].x_c[3].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[3].lc_i.i1muxa1  (.A0(net23),
    .A1(net9),
    .S(\y_c[5].x_c[3].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[3].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[3].lc_i.i1muxb  (.A0(\y_c[5].x_c[3].lc_i.i1a ),
    .A1(\y_c[5].x_c[3].lc_i.i1b ),
    .S(\y_c[5].x_c[3].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[3].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[5].x_c[3].lc_i.lmux  (.A0(\y_c[5].x_c[3].lc_i.i0 ),
    .A1(\y_c[5].x_c[3].lc_i.i1 ),
    .S(\y_c[5].x_c[3].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[3].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[5].x_c[3].lc_i.s0muxa0  (.A(net20),
    .B(\y_c[5].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[3].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[3].lc_i.s0muxa1  (.A0(net9),
    .A1(net24),
    .S(\y_c[5].x_c[3].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[3].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[5].x_c[3].lc_i.s0muxb  (.A0(\y_c[5].x_c[3].lc_i.s0a ),
    .A1(\y_c[5].x_c[3].lc_i.s0b ),
    .S(\y_c[5].x_c[3].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[3].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_2 \y_c[5].x_c[3].lc_i.sinv  (.A(\y_c[5].x_c[3].lc_i.s0s ),
    .B(\y_c[5].x_c[3].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[3].lc_i.s0 ));
 sky130_fd_sc_hd__dfsbp_1 \y_c[5].x_c[4].lc_i.dff.dff  (.CLK(clknet_2_1__leaf_io_in[0]),
    .D(\y_c[5].x_c[4].lc_i.muxo_n ),
    .SET_B(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[4].lc_i.dff.dffo_n ));
 sky130_fd_sc_hd__mux2i_4 \y_c[5].x_c[4].lc_i.dff.ffsel  (.A0(\y_c[5].x_c[4].lc_i.muxo_n ),
    .A1(\y_c[5].x_c[4].lc_i.dff.dffo_n ),
    .S(\y_c[5].x_c[4].lc_i.cfg[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[4].x_c[4].lc_i.B ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[4].lc_i.genblk1[0].genblk1[0].cfg_lat_i  (.D(\y_c[0].x_c[4].lc_i.cfg_data[0] ),
    .GATE_N(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[4].lc_i.cfg[0] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[4].lc_i.genblk1[0].genblk1[1].cfg_lat_i  (.D(\y_c[0].x_c[4].lc_i.cfg_data[1] ),
    .GATE_N(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[4].lc_i.cfg[1] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[4].lc_i.genblk1[0].genblk1[2].cfg_lat_i  (.D(net153),
    .GATE_N(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[4].lc_i.cfg[2] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[4].lc_i.genblk1[0].genblk1[3].cfg_lat_i  (.D(net149),
    .GATE_N(net124),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[4].lc_i.cfg[3] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[4].lc_i.genblk1[1].genblk1[0].cfg_lat_i  (.D(\y_c[0].x_c[4].lc_i.cfg_data[0] ),
    .GATE_N(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[4].lc_i.cfg[4] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[4].lc_i.genblk1[1].genblk1[1].cfg_lat_i  (.D(\y_c[0].x_c[4].lc_i.cfg_data[1] ),
    .GATE_N(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[4].lc_i.cfg[5] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[4].lc_i.genblk1[1].genblk1[2].cfg_lat_i  (.D(net152),
    .GATE_N(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[4].lc_i.cfg[6] ));
 sky130_fd_sc_hd__dlxtn_1 \y_c[5].x_c[4].lc_i.genblk1[1].genblk1[3].cfg_lat_i  (.D(net147),
    .GATE_N(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\y_c[5].x_c[4].lc_i.cfg[7] ));
 sky130_fd_sc_hd__nand2_1 \y_c[5].x_c[4].lc_i.i0muxa0  (.A(net10),
    .B(\y_c[5].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[4].lc_i.i0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[4].lc_i.i0muxa1  (.A0(net8),
    .A1(net22),
    .S(\y_c[5].x_c[4].lc_i.cfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[4].lc_i.i0b ));
 sky130_fd_sc_hd__mux2i_2 \y_c[5].x_c[4].lc_i.i0muxb  (.A0(\y_c[5].x_c[4].lc_i.i0a ),
    .A1(\y_c[5].x_c[4].lc_i.i0b ),
    .S(\y_c[5].x_c[4].lc_i.cfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[4].lc_i.i0 ));
 sky130_fd_sc_hd__and2_1 \y_c[5].x_c[4].lc_i.i1muxa0  (.A(\y_c[5].x_c[4].lc_i.cfg[2] ),
    .B(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\y_c[5].x_c[4].lc_i.i1a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[4].lc_i.i1muxa1  (.A0(net8),
    .A1(net8),
    .S(\y_c[5].x_c[4].lc_i.cfg[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[4].lc_i.i1b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[4].lc_i.i1muxb  (.A0(\y_c[5].x_c[4].lc_i.i1a ),
    .A1(\y_c[5].x_c[4].lc_i.i1b ),
    .S(\y_c[5].x_c[4].lc_i.cfg[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[4].lc_i.i1 ));
 sky130_fd_sc_hd__mux2i_4 \y_c[5].x_c[4].lc_i.lmux  (.A0(\y_c[5].x_c[4].lc_i.i0 ),
    .A1(\y_c[5].x_c[4].lc_i.i1 ),
    .S(\y_c[5].x_c[4].lc_i.s0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[4].lc_i.muxo_n ));
 sky130_fd_sc_hd__nand2_1 \y_c[5].x_c[4].lc_i.s0muxa0  (.A(net10),
    .B(\y_c[5].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[4].lc_i.s0a ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[4].lc_i.s0muxa1  (.A0(\y_c[4].x_c[4].lc_i.B ),
    .A1(net22),
    .S(\y_c[5].x_c[4].lc_i.cfg[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[4].lc_i.s0b ));
 sky130_fd_sc_hd__mux2i_1 \y_c[5].x_c[4].lc_i.s0muxb  (.A0(\y_c[5].x_c[4].lc_i.s0a ),
    .A1(\y_c[5].x_c[4].lc_i.s0b ),
    .S(\y_c[5].x_c[4].lc_i.cfg[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[4].lc_i.s0s ));
 sky130_fd_sc_hd__xnor2_1 \y_c[5].x_c[4].lc_i.sinv  (.A(\y_c[5].x_c[4].lc_i.s0s ),
    .B(\y_c[5].x_c[4].lc_i.cfg[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\y_c[5].x_c[4].lc_i.s0 ));
endmodule
