VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_module_347688030570545747
  CLASS BLOCK ;
  FOREIGN user_module_347688030570545747 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 120.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 2.000 4.040 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.000 11.520 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.000 19.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.000 26.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.000 33.960 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.000 41.440 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.000 48.920 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.000 56.400 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 2.000 63.880 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 2.000 71.360 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.000 78.840 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.000 86.320 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.000 93.800 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.000 101.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 2.000 108.760 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.000 116.240 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.590 5.200 16.190 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.330 5.200 35.930 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.070 5.200 55.670 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.810 5.200 75.410 114.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.460 5.200 26.060 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.200 5.200 45.800 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.940 5.200 65.540 114.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 84.180 114.325 ;
      LAYER met1 ;
        RECT 5.520 5.200 84.180 114.480 ;
      LAYER met2 ;
        RECT 6.990 3.555 75.380 116.125 ;
      LAYER met3 ;
        RECT 2.400 115.240 75.400 116.105 ;
        RECT 2.000 109.160 75.400 115.240 ;
        RECT 2.400 107.760 75.400 109.160 ;
        RECT 2.000 101.680 75.400 107.760 ;
        RECT 2.400 100.280 75.400 101.680 ;
        RECT 2.000 94.200 75.400 100.280 ;
        RECT 2.400 92.800 75.400 94.200 ;
        RECT 2.000 86.720 75.400 92.800 ;
        RECT 2.400 85.320 75.400 86.720 ;
        RECT 2.000 79.240 75.400 85.320 ;
        RECT 2.400 77.840 75.400 79.240 ;
        RECT 2.000 71.760 75.400 77.840 ;
        RECT 2.400 70.360 75.400 71.760 ;
        RECT 2.000 64.280 75.400 70.360 ;
        RECT 2.400 62.880 75.400 64.280 ;
        RECT 2.000 56.800 75.400 62.880 ;
        RECT 2.400 55.400 75.400 56.800 ;
        RECT 2.000 49.320 75.400 55.400 ;
        RECT 2.400 47.920 75.400 49.320 ;
        RECT 2.000 41.840 75.400 47.920 ;
        RECT 2.400 40.440 75.400 41.840 ;
        RECT 2.000 34.360 75.400 40.440 ;
        RECT 2.400 32.960 75.400 34.360 ;
        RECT 2.000 26.880 75.400 32.960 ;
        RECT 2.400 25.480 75.400 26.880 ;
        RECT 2.000 19.400 75.400 25.480 ;
        RECT 2.400 18.000 75.400 19.400 ;
        RECT 2.000 11.920 75.400 18.000 ;
        RECT 2.400 10.520 75.400 11.920 ;
        RECT 2.000 4.440 75.400 10.520 ;
        RECT 2.400 3.575 75.400 4.440 ;
  END
END user_module_347688030570545747
END LIBRARY

