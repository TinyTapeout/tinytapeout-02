/* Automatically generated from https://wokwi.com/projects/347144898258928211 */

`default_nettype none

module user_module_347144898258928211(
  input [7:0] io_in,
  output [7:0] io_out
);
  wire net1 = io_in[0];
  wire net2 = io_in[6];
  wire net3 = io_in[7];
  wire net4;
  wire net5 = 1'b0;
  wire net6 = 1'b1;
  wire net7 = 1'b1;
  wire net8;
  wire net9;
  wire net10 = 1'b1;
  wire net11;
  wire net12;
  wire net13 = 1'b1;
  wire net14;
  wire net15;
  wire net16 = 1'b1;
  wire net17;
  wire net18;
  wire net19 = 1'b1;
  wire net20;
  wire net21;
  wire net22 = 1'b0;
  wire net23;
  wire net24;
  wire net25 = 1'b0;
  wire net26;
  wire net27;
  wire net28 = 1'b0;
  wire net29;
  wire net30;
  wire net31 = 1'b1;
  wire net32;
  wire net33;
  wire net34 = 1'b0;
  wire net35;
  wire net36;
  wire net37 = 1'b1;
  wire net38;
  wire net39;
  wire net40 = 1'b0;
  wire net41;
  wire net42;
  wire net43 = 1'b1;
  wire net44;
  wire net45;
  wire net46 = 1'b0;
  wire net47;
  wire net48;
  wire net49 = 1'b1;
  wire net50;
  wire net51;
  wire net52 = 1'b1;
  wire net53;
  wire net54;
  wire net55 = 1'b1;
  wire net56;
  wire net57;
  wire net58 = 1'b1;
  wire net59;
  wire net60 = 1'b0;
  wire net61 = 1'b0;
  wire net62 = 1'b0;
  wire net63;
  wire net64;
  wire net65 = 1'b1;
  wire net66;
  wire net67;
  wire net68 = 1'b1;
  wire net69;
  wire net70;
  wire net71 = 1'b1;
  wire net72;
  wire net73;
  wire net74 = 1'b1;
  wire net75;
  wire net76;
  wire net77 = 1'b0;
  wire net78;
  wire net79;
  wire net80 = 1'b1;
  wire net81;
  wire net82;
  wire net83 = 1'b0;
  wire net84;
  wire net85;
  wire net86 = 1'b0;
  wire net87;
  wire net88;
  wire net89 = 1'b1;
  wire net90;
  wire net91;
  wire net92 = 1'b0;
  wire net93;
  wire net94;
  wire net95 = 1'b1;
  wire net96;
  wire net97;
  wire net98 = 1'b1;
  wire net99;
  wire net100;
  wire net101 = 1'b0;
  wire net102;
  wire net103;
  wire net104 = 1'b1;
  wire net105;
  wire net106;
  wire net107 = 1'b1;
  wire net108;
  wire net109;
  wire net110 = 1'b1;
  wire net111;
  wire net112;
  wire net113 = 1'b1;
  wire net114;
  wire net115 = 1'b0;
  wire net116;
  wire net117 = 1'b1;
  wire net118;
  wire net119;
  wire net120 = 1'b1;
  wire net121;
  wire net122;
  wire net123 = 1'b1;
  wire net124;
  wire net125;
  wire net126 = 1'b1;
  wire net127;
  wire net128;
  wire net129 = 1'b1;
  wire net130;
  wire net131;
  wire net132 = 1'b1;
  wire net133;
  wire net134;
  wire net135 = 1'b1;
  wire net136;
  wire net137;
  wire net138 = 1'b1;
  wire net139;
  wire net140;
  wire net141 = 1'b1;
  wire net142;
  wire net143;
  wire net144 = 1'b1;
  wire net145;
  wire net146;
  wire net147 = 1'b1;
  wire net148;
  wire net149;
  wire net150 = 1'b1;
  wire net151;
  wire net152;
  wire net153 = 1'b0;
  wire net154;
  wire net155;
  wire net156 = 1'b0;
  wire net157;
  wire net158;
  wire net159 = 1'b1;
  wire net160;
  wire net161;
  wire net162 = 1'b1;
  wire net163;
  wire net164;
  wire net165 = 1'b1;
  wire net166;
  wire net167;
  wire net168 = 1'b0;
  wire net169;
  wire net170;
  wire net171 = 1'b1;
  wire net172;
  wire net173;
  wire net174 = 1'b1;
  wire net175;
  wire net176;
  wire net177 = 1'b0;
  wire net178;
  wire net179;
  wire net180 = 1'b1;
  wire net181;
  wire net182;
  wire net183 = 1'b1;
  wire net184;
  wire net185;
  wire net186 = 1'b1;
  wire net187;
  wire net188;
  wire net189 = 1'b1;
  wire net190;
  wire net191 = 1'b0;
  wire net192;
  wire net193 = 1'b1;
  wire net194;
  wire net195;
  wire net196 = 1'b1;
  wire net197;
  wire net198;
  wire net199 = 1'b1;
  wire net200;
  wire net201;
  wire net202 = 1'b1;
  wire net203;
  wire net204;
  wire net205 = 1'b1;
  wire net206;
  wire net207;
  wire net208 = 1'b1;
  wire net209;
  wire net210;
  wire net211 = 1'b1;
  wire net212;
  wire net213;
  wire net214 = 1'b1;
  wire net215;
  wire net216;
  wire net217 = 1'b0;
  wire net218;
  wire net219;
  wire net220 = 1'b1;
  wire net221;
  wire net222;
  wire net223 = 1'b0;
  wire net224;
  wire net225;
  wire net226 = 1'b0;
  wire net227;
  wire net228;
  wire net229 = 1'b1;
  wire net230;
  wire net231;
  wire net232 = 1'b1;
  wire net233;
  wire net234;
  wire net235 = 1'b1;
  wire net236;
  wire net237;
  wire net238 = 1'b1;
  wire net239;
  wire net240;
  wire net241 = 1'b0;
  wire net242;
  wire net243;
  wire net244 = 1'b1;
  wire net245;
  wire net246;
  wire net247 = 1'b1;
  wire net248;
  wire net249;
  wire net250 = 1'b1;
  wire net251;
  wire net252;
  wire net253 = 1'b1;
  wire net254;
  wire net255 = 1'b0;
  wire net256;
  wire net257 = 1'b1;
  wire net258;
  wire net259;
  wire net260 = 1'b1;
  wire net261;
  wire net262;
  wire net263 = 1'b1;
  wire net264;
  wire net265;
  wire net266 = 1'b1;
  wire net267;
  wire net268;
  wire net269 = 1'b1;
  wire net270;
  wire net271;
  wire net272 = 1'b1;
  wire net273;
  wire net274;
  wire net275 = 1'b1;
  wire net276;
  wire net277;
  wire net278 = 1'b1;
  wire net279;
  wire net280;
  wire net281 = 1'b0;
  wire net282;
  wire net283;
  wire net284 = 1'b0;
  wire net285;
  wire net286;
  wire net287 = 1'b1;
  wire net288;
  wire net289;
  wire net290 = 1'b0;
  wire net291;
  wire net292;
  wire net293 = 1'b1;
  wire net294;
  wire net295;
  wire net296 = 1'b0;
  wire net297;
  wire net298;
  wire net299 = 1'b0;
  wire net300;
  wire net301;
  wire net302 = 1'b0;
  wire net303;
  wire net304;
  wire net305 = 1'b0;
  wire net306;
  wire net307;
  wire net308 = 1'b1;
  wire net309;
  wire net310;
  wire net311 = 1'b1;
  wire net312;
  wire net313;
  wire net314 = 1'b1;
  wire net315;
  wire net316;
  wire net317 = 1'b1;
  wire net318 = 1'b0;
  wire net319;
  wire net320 = 1'b1;
  wire net321;
  wire net322;
  wire net323 = 1'b1;
  wire net324;
  wire net325;
  wire net326 = 1'b1;
  wire net327;
  wire net328;
  wire net329 = 1'b1;
  wire net330 = 1'b1;

  assign io_out[0] = net3;
  assign io_out[1] = net2;
  assign io_out[7] = net4;

  dff_cell flop1 (
    .d (net8),
    .clk (net1),
    .q (net9)
  );
  mux_cell mux1 (
    .a (net10),
    .b (net11),
    .sel (net2),
    .out (net8)
  );
  dff_cell flop3 (
    .d (net12),
    .clk (net1),
    .q (net11)
  );
  mux_cell mux3 (
    .a (net13),
    .b (net14),
    .sel (net2),
    .out (net12)
  );
  dff_cell flop4 (
    .d (net15),
    .clk (net1),
    .q (net14)
  );
  mux_cell mux4 (
    .a (net16),
    .b (net17),
    .sel (net2),
    .out (net15)
  );
  dff_cell flop5 (
    .d (net18),
    .clk (net1),
    .q (net17)
  );
  mux_cell mux5 (
    .a (net19),
    .b (net20),
    .sel (net2),
    .out (net18)
  );
  dff_cell flop6 (
    .d (net21),
    .clk (net1),
    .q (net20)
  );
  mux_cell mux6 (
    .a (net22),
    .b (net23),
    .sel (net2),
    .out (net21)
  );
  dff_cell flop7 (
    .d (net24),
    .clk (net1),
    .q (net23)
  );
  mux_cell mux7 (
    .a (net25),
    .b (net26),
    .sel (net2),
    .out (net24)
  );
  dff_cell flop8 (
    .d (net27),
    .clk (net1),
    .q (net26)
  );
  mux_cell mux8 (
    .a (net28),
    .b (net29),
    .sel (net2),
    .out (net27)
  );
  dff_cell flop9 (
    .d (net30),
    .clk (net1),
    .q (net29)
  );
  mux_cell mux9 (
    .a (net31),
    .b (net32),
    .sel (net2),
    .out (net30)
  );
  dff_cell flop10 (
    .d (net33),
    .clk (net1),
    .q (net32)
  );
  mux_cell mux10 (
    .a (net34),
    .b (net35),
    .sel (net2),
    .out (net33)
  );
  dff_cell flop11 (
    .d (net36),
    .clk (net1),
    .q (net35)
  );
  mux_cell mux11 (
    .a (net37),
    .b (net38),
    .sel (net2),
    .out (net36)
  );
  dff_cell flop12 (
    .d (net39),
    .clk (net1),
    .q (net38)
  );
  mux_cell mux12 (
    .a (net40),
    .b (net41),
    .sel (net2),
    .out (net39)
  );
  dff_cell flop13 (
    .d (net42),
    .clk (net1),
    .q (net41)
  );
  mux_cell mux13 (
    .a (net43),
    .b (net44),
    .sel (net2),
    .out (net42)
  );
  dff_cell flop14 (
    .d (net45),
    .clk (net1),
    .q (net44)
  );
  mux_cell mux14 (
    .a (net46),
    .b (net47),
    .sel (net2),
    .out (net45)
  );
  dff_cell flop15 (
    .d (net48),
    .clk (net1),
    .q (net47)
  );
  mux_cell mux15 (
    .a (net49),
    .b (net50),
    .sel (net2),
    .out (net48)
  );
  dff_cell flop16 (
    .d (net51),
    .clk (net1),
    .q (net50)
  );
  mux_cell mux16 (
    .a (net52),
    .b (net53),
    .sel (net2),
    .out (net51)
  );
  dff_cell flop17 (
    .d (net54),
    .clk (net1),
    .q (net53)
  );
  mux_cell mux17 (
    .a (net55),
    .b (net56),
    .sel (net2),
    .out (net54)
  );
  dff_cell flop18 (
    .d (net57),
    .clk (net1),
    .q (net56)
  );
  mux_cell mux18 (
    .a (net58),
    .b (net59),
    .sel (net2),
    .out (net57)
  );
  dff_cell flop2 (
    .d (net63),
    .clk (net1),
    .q (net64)
  );
  mux_cell mux19 (
    .a (net65),
    .b (net66),
    .sel (net2),
    .out (net63)
  );
  dff_cell flop19 (
    .d (net67),
    .clk (net1),
    .q (net66)
  );
  mux_cell mux20 (
    .a (net68),
    .b (net69),
    .sel (net2),
    .out (net67)
  );
  dff_cell flop20 (
    .d (net70),
    .clk (net1),
    .q (net69)
  );
  mux_cell mux21 (
    .a (net71),
    .b (net72),
    .sel (net2),
    .out (net70)
  );
  dff_cell flop21 (
    .d (net73),
    .clk (net1),
    .q (net72)
  );
  mux_cell mux22 (
    .a (net74),
    .b (net75),
    .sel (net2),
    .out (net73)
  );
  dff_cell flop22 (
    .d (net76),
    .clk (net1),
    .q (net75)
  );
  mux_cell mux23 (
    .a (net77),
    .b (net78),
    .sel (net2),
    .out (net76)
  );
  dff_cell flop23 (
    .d (net79),
    .clk (net1),
    .q (net78)
  );
  mux_cell mux24 (
    .a (net80),
    .b (net81),
    .sel (net2),
    .out (net79)
  );
  dff_cell flop24 (
    .d (net82),
    .clk (net1),
    .q (net81)
  );
  mux_cell mux25 (
    .a (net83),
    .b (net84),
    .sel (net2),
    .out (net82)
  );
  dff_cell flop25 (
    .d (net85),
    .clk (net1),
    .q (net84)
  );
  mux_cell mux26 (
    .a (net86),
    .b (net87),
    .sel (net2),
    .out (net85)
  );
  dff_cell flop26 (
    .d (net88),
    .clk (net1),
    .q (net87)
  );
  mux_cell mux27 (
    .a (net89),
    .b (net90),
    .sel (net2),
    .out (net88)
  );
  dff_cell flop27 (
    .d (net91),
    .clk (net1),
    .q (net90)
  );
  mux_cell mux28 (
    .a (net92),
    .b (net93),
    .sel (net2),
    .out (net91)
  );
  dff_cell flop28 (
    .d (net94),
    .clk (net1),
    .q (net93)
  );
  mux_cell mux29 (
    .a (net95),
    .b (net96),
    .sel (net2),
    .out (net94)
  );
  dff_cell flop29 (
    .d (net97),
    .clk (net1),
    .q (net96)
  );
  mux_cell mux30 (
    .a (net98),
    .b (net99),
    .sel (net2),
    .out (net97)
  );
  dff_cell flop30 (
    .d (net100),
    .clk (net1),
    .q (net99)
  );
  mux_cell mux31 (
    .a (net101),
    .b (net102),
    .sel (net2),
    .out (net100)
  );
  dff_cell flop31 (
    .d (net103),
    .clk (net1),
    .q (net102)
  );
  mux_cell mux32 (
    .a (net104),
    .b (net105),
    .sel (net2),
    .out (net103)
  );
  dff_cell flop32 (
    .d (net106),
    .clk (net1),
    .q (net105)
  );
  mux_cell mux33 (
    .a (net107),
    .b (net108),
    .sel (net2),
    .out (net106)
  );
  dff_cell flop33 (
    .d (net109),
    .clk (net1),
    .q (net108)
  );
  mux_cell mux34 (
    .a (net110),
    .b (net111),
    .sel (net2),
    .out (net109)
  );
  dff_cell flop34 (
    .d (net112),
    .clk (net1),
    .q (net111)
  );
  mux_cell mux35 (
    .a (net113),
    .b (net114),
    .sel (net2),
    .out (net112)
  );
  dff_cell flop35 (
    .d (net116),
    .clk (net1),
    .q (net59)
  );
  mux_cell mux36 (
    .a (net117),
    .b (net118),
    .sel (net2),
    .out (net116)
  );
  dff_cell flop36 (
    .d (net119),
    .clk (net1),
    .q (net118)
  );
  mux_cell mux37 (
    .a (net120),
    .b (net121),
    .sel (net2),
    .out (net119)
  );
  dff_cell flop37 (
    .d (net122),
    .clk (net1),
    .q (net121)
  );
  mux_cell mux38 (
    .a (net123),
    .b (net124),
    .sel (net2),
    .out (net122)
  );
  dff_cell flop38 (
    .d (net125),
    .clk (net1),
    .q (net124)
  );
  mux_cell mux39 (
    .a (net126),
    .b (net64),
    .sel (net2),
    .out (net125)
  );
  dff_cell flop39 (
    .d (net127),
    .clk (net1),
    .q (net128)
  );
  mux_cell mux40 (
    .a (net129),
    .b (net130),
    .sel (net2),
    .out (net127)
  );
  dff_cell flop40 (
    .d (net131),
    .clk (net1),
    .q (net130)
  );
  mux_cell mux41 (
    .a (net132),
    .b (net133),
    .sel (net2),
    .out (net131)
  );
  dff_cell flop41 (
    .d (net134),
    .clk (net1),
    .q (net133)
  );
  mux_cell mux42 (
    .a (net135),
    .b (net136),
    .sel (net2),
    .out (net134)
  );
  dff_cell flop42 (
    .d (net137),
    .clk (net1),
    .q (net136)
  );
  mux_cell mux43 (
    .a (net138),
    .b (net9),
    .sel (net2),
    .out (net137)
  );
  dff_cell flop43 (
    .d (net139),
    .clk (net1),
    .q (net140)
  );
  mux_cell mux44 (
    .a (net141),
    .b (net142),
    .sel (net2),
    .out (net139)
  );
  dff_cell flop44 (
    .d (net143),
    .clk (net1),
    .q (net142)
  );
  mux_cell mux45 (
    .a (net144),
    .b (net145),
    .sel (net2),
    .out (net143)
  );
  dff_cell flop45 (
    .d (net146),
    .clk (net1),
    .q (net145)
  );
  mux_cell mux46 (
    .a (net147),
    .b (net148),
    .sel (net2),
    .out (net146)
  );
  dff_cell flop46 (
    .d (net149),
    .clk (net1),
    .q (net148)
  );
  mux_cell mux47 (
    .a (net150),
    .b (net151),
    .sel (net2),
    .out (net149)
  );
  dff_cell flop47 (
    .d (net152),
    .clk (net1),
    .q (net151)
  );
  mux_cell mux48 (
    .a (net153),
    .b (net154),
    .sel (net2),
    .out (net152)
  );
  dff_cell flop48 (
    .d (net155),
    .clk (net1),
    .q (net154)
  );
  mux_cell mux49 (
    .a (net156),
    .b (net157),
    .sel (net2),
    .out (net155)
  );
  dff_cell flop49 (
    .d (net158),
    .clk (net1),
    .q (net157)
  );
  mux_cell mux50 (
    .a (net159),
    .b (net160),
    .sel (net2),
    .out (net158)
  );
  dff_cell flop50 (
    .d (net161),
    .clk (net1),
    .q (net160)
  );
  mux_cell mux51 (
    .a (net162),
    .b (net163),
    .sel (net2),
    .out (net161)
  );
  dff_cell flop51 (
    .d (net164),
    .clk (net1),
    .q (net163)
  );
  mux_cell mux52 (
    .a (net165),
    .b (net166),
    .sel (net2),
    .out (net164)
  );
  dff_cell flop52 (
    .d (net167),
    .clk (net1),
    .q (net166)
  );
  mux_cell mux53 (
    .a (net168),
    .b (net169),
    .sel (net2),
    .out (net167)
  );
  dff_cell flop53 (
    .d (net170),
    .clk (net1),
    .q (net169)
  );
  mux_cell mux54 (
    .a (net171),
    .b (net172),
    .sel (net2),
    .out (net170)
  );
  dff_cell flop54 (
    .d (net173),
    .clk (net1),
    .q (net172)
  );
  mux_cell mux55 (
    .a (net174),
    .b (net175),
    .sel (net2),
    .out (net173)
  );
  dff_cell flop55 (
    .d (net176),
    .clk (net1),
    .q (net175)
  );
  mux_cell mux56 (
    .a (net177),
    .b (net178),
    .sel (net2),
    .out (net176)
  );
  dff_cell flop56 (
    .d (net179),
    .clk (net1),
    .q (net178)
  );
  mux_cell mux57 (
    .a (net180),
    .b (net181),
    .sel (net2),
    .out (net179)
  );
  dff_cell flop57 (
    .d (net182),
    .clk (net1),
    .q (net181)
  );
  mux_cell mux58 (
    .a (net183),
    .b (net184),
    .sel (net2),
    .out (net182)
  );
  dff_cell flop58 (
    .d (net185),
    .clk (net1),
    .q (net184)
  );
  mux_cell mux59 (
    .a (net186),
    .b (net187),
    .sel (net2),
    .out (net185)
  );
  dff_cell flop59 (
    .d (net188),
    .clk (net1),
    .q (net187)
  );
  mux_cell mux60 (
    .a (net189),
    .b (net190),
    .sel (net2),
    .out (net188)
  );
  dff_cell flop60 (
    .d (net192),
    .clk (net1),
    .q (net114)
  );
  mux_cell mux61 (
    .a (net193),
    .b (net194),
    .sel (net2),
    .out (net192)
  );
  dff_cell flop61 (
    .d (net195),
    .clk (net1),
    .q (net194)
  );
  mux_cell mux62 (
    .a (net196),
    .b (net197),
    .sel (net2),
    .out (net195)
  );
  dff_cell flop62 (
    .d (net198),
    .clk (net1),
    .q (net197)
  );
  mux_cell mux63 (
    .a (net199),
    .b (net200),
    .sel (net2),
    .out (net198)
  );
  dff_cell flop63 (
    .d (net201),
    .clk (net1),
    .q (net200)
  );
  mux_cell mux64 (
    .a (net202),
    .b (net140),
    .sel (net2),
    .out (net201)
  );
  dff_cell flop64 (
    .d (net203),
    .clk (net1),
    .q (net204)
  );
  mux_cell mux65 (
    .a (net205),
    .b (net206),
    .sel (net2),
    .out (net203)
  );
  dff_cell flop65 (
    .d (net207),
    .clk (net1),
    .q (net206)
  );
  mux_cell mux66 (
    .a (net208),
    .b (net209),
    .sel (net2),
    .out (net207)
  );
  dff_cell flop66 (
    .d (net210),
    .clk (net1),
    .q (net209)
  );
  mux_cell mux67 (
    .a (net211),
    .b (net212),
    .sel (net2),
    .out (net210)
  );
  dff_cell flop67 (
    .d (net213),
    .clk (net1),
    .q (net212)
  );
  mux_cell mux68 (
    .a (net214),
    .b (net215),
    .sel (net2),
    .out (net213)
  );
  dff_cell flop68 (
    .d (net216),
    .clk (net1),
    .q (net215)
  );
  mux_cell mux69 (
    .a (net217),
    .b (net218),
    .sel (net2),
    .out (net216)
  );
  dff_cell flop69 (
    .d (net219),
    .clk (net1),
    .q (net218)
  );
  mux_cell mux70 (
    .a (net220),
    .b (net221),
    .sel (net2),
    .out (net219)
  );
  dff_cell flop70 (
    .d (net222),
    .clk (net1),
    .q (net221)
  );
  mux_cell mux71 (
    .a (net223),
    .b (net224),
    .sel (net2),
    .out (net222)
  );
  dff_cell flop71 (
    .d (net225),
    .clk (net1),
    .q (net224)
  );
  mux_cell mux72 (
    .a (net226),
    .b (net227),
    .sel (net2),
    .out (net225)
  );
  dff_cell flop72 (
    .d (net228),
    .clk (net1),
    .q (net227)
  );
  mux_cell mux73 (
    .a (net229),
    .b (net230),
    .sel (net2),
    .out (net228)
  );
  dff_cell flop73 (
    .d (net231),
    .clk (net1),
    .q (net230)
  );
  mux_cell mux74 (
    .a (net232),
    .b (net233),
    .sel (net2),
    .out (net231)
  );
  dff_cell flop74 (
    .d (net234),
    .clk (net1),
    .q (net233)
  );
  mux_cell mux75 (
    .a (net235),
    .b (net236),
    .sel (net2),
    .out (net234)
  );
  dff_cell flop75 (
    .d (net237),
    .clk (net1),
    .q (net236)
  );
  mux_cell mux76 (
    .a (net238),
    .b (net239),
    .sel (net2),
    .out (net237)
  );
  dff_cell flop76 (
    .d (net240),
    .clk (net1),
    .q (net239)
  );
  mux_cell mux77 (
    .a (net241),
    .b (net242),
    .sel (net2),
    .out (net240)
  );
  dff_cell flop77 (
    .d (net243),
    .clk (net1),
    .q (net242)
  );
  mux_cell mux78 (
    .a (net244),
    .b (net245),
    .sel (net2),
    .out (net243)
  );
  dff_cell flop78 (
    .d (net246),
    .clk (net1),
    .q (net245)
  );
  mux_cell mux79 (
    .a (net247),
    .b (net248),
    .sel (net2),
    .out (net246)
  );
  dff_cell flop79 (
    .d (net249),
    .clk (net1),
    .q (net248)
  );
  mux_cell mux80 (
    .a (net250),
    .b (net251),
    .sel (net2),
    .out (net249)
  );
  dff_cell flop80 (
    .d (net252),
    .clk (net1),
    .q (net251)
  );
  mux_cell mux81 (
    .a (net253),
    .b (net254),
    .sel (net2),
    .out (net252)
  );
  dff_cell flop81 (
    .d (net256),
    .clk (net1),
    .q (net190)
  );
  mux_cell mux82 (
    .a (net257),
    .b (net258),
    .sel (net2),
    .out (net256)
  );
  dff_cell flop82 (
    .d (net259),
    .clk (net1),
    .q (net258)
  );
  mux_cell mux83 (
    .a (net260),
    .b (net261),
    .sel (net2),
    .out (net259)
  );
  dff_cell flop83 (
    .d (net262),
    .clk (net1),
    .q (net261)
  );
  mux_cell mux84 (
    .a (net263),
    .b (net264),
    .sel (net2),
    .out (net262)
  );
  dff_cell flop84 (
    .d (net265),
    .clk (net1),
    .q (net264)
  );
  mux_cell mux85 (
    .a (net266),
    .b (net204),
    .sel (net2),
    .out (net265)
  );
  dff_cell flop85 (
    .d (net267),
    .clk (net1),
    .q (net268)
  );
  mux_cell mux86 (
    .a (net269),
    .b (net270),
    .sel (net2),
    .out (net267)
  );
  dff_cell flop86 (
    .d (net271),
    .clk (net1),
    .q (net270)
  );
  mux_cell mux87 (
    .a (net272),
    .b (net273),
    .sel (net2),
    .out (net271)
  );
  dff_cell flop87 (
    .d (net274),
    .clk (net1),
    .q (net273)
  );
  mux_cell mux88 (
    .a (net275),
    .b (net276),
    .sel (net2),
    .out (net274)
  );
  dff_cell flop88 (
    .d (net277),
    .clk (net1),
    .q (net276)
  );
  mux_cell mux89 (
    .a (net278),
    .b (net279),
    .sel (net2),
    .out (net277)
  );
  dff_cell flop89 (
    .d (net280),
    .clk (net1),
    .q (net279)
  );
  mux_cell mux90 (
    .a (net281),
    .b (net282),
    .sel (net2),
    .out (net280)
  );
  dff_cell flop90 (
    .d (net283),
    .clk (net1),
    .q (net282)
  );
  mux_cell mux91 (
    .a (net284),
    .b (net285),
    .sel (net2),
    .out (net283)
  );
  dff_cell flop91 (
    .d (net286),
    .clk (net1),
    .q (net285)
  );
  mux_cell mux92 (
    .a (net287),
    .b (net288),
    .sel (net2),
    .out (net286)
  );
  dff_cell flop92 (
    .d (net289),
    .clk (net1),
    .q (net288)
  );
  mux_cell mux93 (
    .a (net290),
    .b (net291),
    .sel (net2),
    .out (net289)
  );
  dff_cell flop93 (
    .d (net292),
    .clk (net1),
    .q (net291)
  );
  mux_cell mux94 (
    .a (net293),
    .b (net294),
    .sel (net2),
    .out (net292)
  );
  dff_cell flop94 (
    .d (net295),
    .clk (net1),
    .q (net294)
  );
  mux_cell mux95 (
    .a (net296),
    .b (net297),
    .sel (net2),
    .out (net295)
  );
  dff_cell flop95 (
    .d (net298),
    .clk (net1),
    .q (net297)
  );
  mux_cell mux96 (
    .a (net299),
    .b (net300),
    .sel (net2),
    .out (net298)
  );
  dff_cell flop96 (
    .d (net301),
    .clk (net1),
    .q (net300)
  );
  mux_cell mux97 (
    .a (net302),
    .b (net303),
    .sel (net2),
    .out (net301)
  );
  dff_cell flop97 (
    .d (net304),
    .clk (net1),
    .q (net303)
  );
  mux_cell mux98 (
    .a (net305),
    .b (net306),
    .sel (net2),
    .out (net304)
  );
  dff_cell flop98 (
    .d (net307),
    .clk (net1),
    .q (net306)
  );
  mux_cell mux99 (
    .a (net308),
    .b (net309),
    .sel (net2),
    .out (net307)
  );
  dff_cell flop99 (
    .d (net310),
    .clk (net1),
    .q (net309)
  );
  mux_cell mux100 (
    .a (net311),
    .b (net312),
    .sel (net2),
    .out (net310)
  );
  dff_cell flop100 (
    .d (net313),
    .clk (net1),
    .q (net312)
  );
  mux_cell mux101 (
    .a (net314),
    .b (net315),
    .sel (net2),
    .out (net313)
  );
  dff_cell flop101 (
    .d (net316),
    .clk (net1),
    .q (net315)
  );
  mux_cell mux102 (
    .a (net317),
    .b (net4),
    .sel (net2),
    .out (net316)
  );
  dff_cell flop102 (
    .d (net319),
    .clk (net1),
    .q (net254)
  );
  mux_cell mux103 (
    .a (net320),
    .b (net321),
    .sel (net2),
    .out (net319)
  );
  dff_cell flop103 (
    .d (net322),
    .clk (net1),
    .q (net321)
  );
  mux_cell mux104 (
    .a (net323),
    .b (net324),
    .sel (net2),
    .out (net322)
  );
  dff_cell flop104 (
    .d (net325),
    .clk (net1),
    .q (net324)
  );
  mux_cell mux105 (
    .a (net326),
    .b (net327),
    .sel (net2),
    .out (net325)
  );
  dff_cell flop105 (
    .d (net328),
    .clk (net1),
    .q (net327)
  );
  mux_cell mux106 (
    .a (net329),
    .b (net268),
    .sel (net2),
    .out (net328)
  );
  mux_cell mux2 (
    .a (net330),
    .b (net128),
    .sel (net3),
    .out (net4)
  );
endmodule
