magic
tech sky130B
magscale 1 2
timestamp 1669906244
<< obsli1 >>
rect 1104 1071 4876 22865
<< obsm1 >>
rect 1104 1040 4954 22896
<< obsm2 >>
rect 1124 711 4948 23225
<< metal3 >>
rect 5200 23128 6000 23248
rect 0 22312 800 22432
rect 5200 21632 6000 21752
rect 5200 20136 6000 20256
rect 0 19320 800 19440
rect 5200 18640 6000 18760
rect 5200 17144 6000 17264
rect 0 16328 800 16448
rect 5200 15648 6000 15768
rect 5200 14152 6000 14272
rect 0 13336 800 13456
rect 5200 12656 6000 12776
rect 5200 11160 6000 11280
rect 0 10344 800 10464
rect 5200 9664 6000 9784
rect 5200 8168 6000 8288
rect 0 7352 800 7472
rect 5200 6672 6000 6792
rect 5200 5176 6000 5296
rect 0 4360 800 4480
rect 5200 3680 6000 3800
rect 5200 2184 6000 2304
rect 0 1368 800 1488
rect 5200 688 6000 808
<< obsm3 >>
rect 798 23048 5120 23221
rect 798 22512 5200 23048
rect 880 22232 5200 22512
rect 798 21832 5200 22232
rect 798 21552 5120 21832
rect 798 20336 5200 21552
rect 798 20056 5120 20336
rect 798 19520 5200 20056
rect 880 19240 5200 19520
rect 798 18840 5200 19240
rect 798 18560 5120 18840
rect 798 17344 5200 18560
rect 798 17064 5120 17344
rect 798 16528 5200 17064
rect 880 16248 5200 16528
rect 798 15848 5200 16248
rect 798 15568 5120 15848
rect 798 14352 5200 15568
rect 798 14072 5120 14352
rect 798 13536 5200 14072
rect 880 13256 5200 13536
rect 798 12856 5200 13256
rect 798 12576 5120 12856
rect 798 11360 5200 12576
rect 798 11080 5120 11360
rect 798 10544 5200 11080
rect 880 10264 5200 10544
rect 798 9864 5200 10264
rect 798 9584 5120 9864
rect 798 8368 5200 9584
rect 798 8088 5120 8368
rect 798 7552 5200 8088
rect 880 7272 5200 7552
rect 798 6872 5200 7272
rect 798 6592 5120 6872
rect 798 5376 5200 6592
rect 798 5096 5120 5376
rect 798 4560 5200 5096
rect 880 4280 5200 4560
rect 798 3880 5200 4280
rect 798 3600 5120 3880
rect 798 2384 5200 3600
rect 798 2104 5120 2384
rect 798 1568 5200 2104
rect 880 1288 5200 1568
rect 798 888 5200 1288
rect 798 715 5120 888
<< metal4 >>
rect 1418 1040 1738 22896
rect 1892 1040 2212 22896
rect 2366 1040 2686 22896
rect 2840 1040 3160 22896
rect 3314 1040 3634 22896
rect 3788 1040 4108 22896
rect 4262 1040 4582 22896
<< labels >>
rlabel metal3 s 0 1368 800 1488 6 clk_in
port 1 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 clk_out
port 2 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 data_in
port 3 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 data_out
port 4 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 latch_enable_in
port 5 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 latch_enable_out
port 6 nsew signal output
rlabel metal3 s 5200 688 6000 808 6 module_data_in[0]
port 7 nsew signal output
rlabel metal3 s 5200 2184 6000 2304 6 module_data_in[1]
port 8 nsew signal output
rlabel metal3 s 5200 3680 6000 3800 6 module_data_in[2]
port 9 nsew signal output
rlabel metal3 s 5200 5176 6000 5296 6 module_data_in[3]
port 10 nsew signal output
rlabel metal3 s 5200 6672 6000 6792 6 module_data_in[4]
port 11 nsew signal output
rlabel metal3 s 5200 8168 6000 8288 6 module_data_in[5]
port 12 nsew signal output
rlabel metal3 s 5200 9664 6000 9784 6 module_data_in[6]
port 13 nsew signal output
rlabel metal3 s 5200 11160 6000 11280 6 module_data_in[7]
port 14 nsew signal output
rlabel metal3 s 5200 12656 6000 12776 6 module_data_out[0]
port 15 nsew signal input
rlabel metal3 s 5200 14152 6000 14272 6 module_data_out[1]
port 16 nsew signal input
rlabel metal3 s 5200 15648 6000 15768 6 module_data_out[2]
port 17 nsew signal input
rlabel metal3 s 5200 17144 6000 17264 6 module_data_out[3]
port 18 nsew signal input
rlabel metal3 s 5200 18640 6000 18760 6 module_data_out[4]
port 19 nsew signal input
rlabel metal3 s 5200 20136 6000 20256 6 module_data_out[5]
port 20 nsew signal input
rlabel metal3 s 5200 21632 6000 21752 6 module_data_out[6]
port 21 nsew signal input
rlabel metal3 s 5200 23128 6000 23248 6 module_data_out[7]
port 22 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 scan_select_in
port 23 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 scan_select_out
port 24 nsew signal output
rlabel metal4 s 1418 1040 1738 22896 6 vccd1
port 25 nsew power bidirectional
rlabel metal4 s 2366 1040 2686 22896 6 vccd1
port 25 nsew power bidirectional
rlabel metal4 s 3314 1040 3634 22896 6 vccd1
port 25 nsew power bidirectional
rlabel metal4 s 4262 1040 4582 22896 6 vccd1
port 25 nsew power bidirectional
rlabel metal4 s 1892 1040 2212 22896 6 vssd1
port 26 nsew ground bidirectional
rlabel metal4 s 2840 1040 3160 22896 6 vssd1
port 26 nsew ground bidirectional
rlabel metal4 s 3788 1040 4108 22896 6 vssd1
port 26 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 6000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 361192
string GDS_FILE /home/matt/work/asic-workshop/shuttle8/tinytapeout-02/openlane/scanchain/runs/22_12_01_15_49/results/signoff/scanchain.magic.gds
string GDS_START 86034
<< end >>

