VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chrisruk_matrix
  CLASS BLOCK ;
  FOREIGN chrisruk_matrix ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 120.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 2.000 4.040 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.000 11.520 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.000 19.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.000 26.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.000 33.960 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.000 41.440 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.000 48.920 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.000 56.400 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 2.000 63.880 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 2.000 71.360 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.000 78.840 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.000 86.320 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.000 93.800 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.000 101.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 2.000 108.760 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.000 116.240 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.590 5.200 16.190 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.330 5.200 35.930 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.070 5.200 55.670 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.810 5.200 75.410 114.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.460 5.200 26.060 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.200 5.200 45.800 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.940 5.200 65.540 114.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 84.180 114.325 ;
      LAYER met1 ;
        RECT 0.070 3.440 85.950 114.480 ;
      LAYER met2 ;
        RECT 0.100 3.410 85.930 116.125 ;
      LAYER met3 ;
        RECT 2.400 115.240 85.955 116.105 ;
        RECT 0.270 109.160 85.955 115.240 ;
        RECT 2.400 107.760 85.955 109.160 ;
        RECT 0.270 101.680 85.955 107.760 ;
        RECT 2.400 100.280 85.955 101.680 ;
        RECT 0.270 94.200 85.955 100.280 ;
        RECT 2.400 92.800 85.955 94.200 ;
        RECT 0.270 86.720 85.955 92.800 ;
        RECT 2.400 85.320 85.955 86.720 ;
        RECT 0.270 79.240 85.955 85.320 ;
        RECT 2.400 77.840 85.955 79.240 ;
        RECT 0.270 71.760 85.955 77.840 ;
        RECT 2.400 70.360 85.955 71.760 ;
        RECT 0.270 64.280 85.955 70.360 ;
        RECT 2.400 62.880 85.955 64.280 ;
        RECT 0.270 56.800 85.955 62.880 ;
        RECT 2.400 55.400 85.955 56.800 ;
        RECT 0.270 49.320 85.955 55.400 ;
        RECT 2.400 47.920 85.955 49.320 ;
        RECT 0.270 41.840 85.955 47.920 ;
        RECT 2.400 40.440 85.955 41.840 ;
        RECT 0.270 34.360 85.955 40.440 ;
        RECT 2.400 32.960 85.955 34.360 ;
        RECT 0.270 26.880 85.955 32.960 ;
        RECT 2.400 25.480 85.955 26.880 ;
        RECT 0.270 19.400 85.955 25.480 ;
        RECT 2.400 18.000 85.955 19.400 ;
        RECT 0.270 11.920 85.955 18.000 ;
        RECT 2.400 10.520 85.955 11.920 ;
        RECT 0.270 4.440 85.955 10.520 ;
        RECT 2.400 3.575 85.955 4.440 ;
      LAYER met4 ;
        RECT 0.295 4.800 14.190 104.545 ;
        RECT 16.590 4.800 24.060 104.545 ;
        RECT 26.460 4.800 33.930 104.545 ;
        RECT 36.330 4.800 43.800 104.545 ;
        RECT 46.200 4.800 53.670 104.545 ;
        RECT 56.070 4.800 63.540 104.545 ;
        RECT 65.940 4.800 73.410 104.545 ;
        RECT 75.810 4.800 84.345 104.545 ;
        RECT 0.295 3.575 84.345 4.800 ;
  END
END chrisruk_matrix
END LIBRARY

