VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fraserbc_simon
  CLASS BLOCK ;
  FOREIGN fraserbc_simon ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 120.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 2.000 4.040 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.000 11.520 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.000 19.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.000 26.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.000 33.960 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.000 41.440 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.000 48.920 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.000 56.400 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 2.000 63.880 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 2.000 71.360 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.000 78.840 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.000 86.320 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.000 93.800 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.000 101.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 2.000 108.760 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.000 116.240 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.550 5.200 16.150 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.215 5.200 35.815 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.880 5.200 55.480 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.545 5.200 75.145 114.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.380 5.200 25.980 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.045 5.200 45.645 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.710 5.200 65.310 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.375 5.200 84.975 114.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 84.180 114.325 ;
      LAYER met1 ;
        RECT 0.070 2.080 90.000 119.920 ;
      LAYER met2 ;
        RECT 0.090 2.050 90.000 119.670 ;
      LAYER met3 ;
        RECT 2.400 115.240 89.890 116.105 ;
        RECT 0.065 109.160 89.890 115.240 ;
        RECT 2.400 107.760 89.890 109.160 ;
        RECT 0.065 101.680 89.890 107.760 ;
        RECT 2.400 100.280 89.890 101.680 ;
        RECT 0.065 94.200 89.890 100.280 ;
        RECT 2.400 92.800 89.890 94.200 ;
        RECT 0.065 86.720 89.890 92.800 ;
        RECT 2.400 85.320 89.890 86.720 ;
        RECT 0.065 79.240 89.890 85.320 ;
        RECT 2.400 77.840 89.890 79.240 ;
        RECT 0.065 71.760 89.890 77.840 ;
        RECT 2.400 70.360 89.890 71.760 ;
        RECT 0.065 64.280 89.890 70.360 ;
        RECT 2.400 62.880 89.890 64.280 ;
        RECT 0.065 56.800 89.890 62.880 ;
        RECT 2.400 55.400 89.890 56.800 ;
        RECT 0.065 49.320 89.890 55.400 ;
        RECT 2.400 47.920 89.890 49.320 ;
        RECT 0.065 41.840 89.890 47.920 ;
        RECT 2.400 40.440 89.890 41.840 ;
        RECT 0.065 34.360 89.890 40.440 ;
        RECT 2.400 32.960 89.890 34.360 ;
        RECT 0.065 26.880 89.890 32.960 ;
        RECT 2.400 25.480 89.890 26.880 ;
        RECT 0.065 19.400 89.890 25.480 ;
        RECT 2.400 18.000 89.890 19.400 ;
        RECT 0.065 11.920 89.890 18.000 ;
        RECT 2.400 10.520 89.890 11.920 ;
        RECT 0.065 4.440 89.890 10.520 ;
        RECT 2.400 3.040 89.890 4.440 ;
        RECT 0.065 2.215 89.890 3.040 ;
      LAYER met4 ;
        RECT 0.295 114.880 89.865 116.105 ;
        RECT 0.295 4.800 14.150 114.880 ;
        RECT 16.550 4.800 23.980 114.880 ;
        RECT 26.380 4.800 33.815 114.880 ;
        RECT 36.215 4.800 43.645 114.880 ;
        RECT 46.045 4.800 53.480 114.880 ;
        RECT 55.880 4.800 63.310 114.880 ;
        RECT 65.710 4.800 73.145 114.880 ;
        RECT 75.545 4.800 82.975 114.880 ;
        RECT 85.375 4.800 89.865 114.880 ;
        RECT 0.295 2.895 89.865 4.800 ;
  END
END fraserbc_simon
END LIBRARY

