module c_tt2_mrcs_test (vccd1,
    vssd1,
    io_in,
    io_out);
 input vccd1;
 input vssd1;
 input [7:0] io_in;
 output [7:0] io_out;

 wire net2;
 wire \SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ;
 wire \SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ;
 wire \SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.out_0 ;
 wire \SavedGate_1.LogicGate_0.in_0 ;
 wire \SavedGate_2.SavedGate_0.LogicGate_0.in_0 ;
 wire \SavedGate_2.SavedGate_0.LogicGate_0.out_0 ;
 wire \SavedGate_4.LogicGate_0.in_0 ;
 wire \SavedGate_4.LogicGate_0.out_0 ;
 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire \clknet_0_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ;
 wire \clknet_0_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ;
 wire \clknet_0_SavedGate_1.LogicGate_0.in_0 ;
 wire \clknet_0_SavedGate_2.SavedGate_0.LogicGate_0.in_0 ;
 wire \clknet_0_SavedGate_4.LogicGate_0.in_0 ;
 wire \clknet_0_SavedGate_4.LogicGate_0.out_0 ;
 wire clknet_0__01_;
 wire clknet_0__02_;
 wire clknet_0__04_;
 wire \clknet_1_0__leaf_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ;
 wire \clknet_1_0__leaf_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ;
 wire \clknet_1_0__leaf_SavedGate_1.LogicGate_0.in_0 ;
 wire \clknet_1_0__leaf_SavedGate_2.SavedGate_0.LogicGate_0.in_0 ;
 wire \clknet_1_0__leaf_SavedGate_4.LogicGate_0.in_0 ;
 wire \clknet_1_0__leaf_SavedGate_4.LogicGate_0.out_0 ;
 wire clknet_1_0__leaf__01_;
 wire clknet_1_0__leaf__02_;
 wire clknet_1_0__leaf__04_;
 wire \clknet_1_1__leaf_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ;
 wire \clknet_1_1__leaf_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ;
 wire \clknet_1_1__leaf_SavedGate_1.LogicGate_0.in_0 ;
 wire \clknet_1_1__leaf_SavedGate_2.SavedGate_0.LogicGate_0.in_0 ;
 wire \clknet_1_1__leaf_SavedGate_4.LogicGate_0.in_0 ;
 wire \clknet_1_1__leaf_SavedGate_4.LogicGate_0.out_0 ;
 wire clknet_1_1__leaf__01_;
 wire clknet_1_1__leaf__02_;
 wire clknet_1_1__leaf__04_;
 wire net1;
 wire [0:0] clknet_0_io_in;
 wire [0:0] clknet_1_0__leaf_io_in;
 wire [0:0] clknet_1_1__leaf_io_in;

 sky130_fd_sc_hd__decap_3 FILLER_0_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_10_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_10_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_10_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_10_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_10_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_11_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_11_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_11_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_11_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_12_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_12_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_12_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_12_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_12_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_13_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_13_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_13_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_13_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_14_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_14_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_14_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_14_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_14_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_15_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_15_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_15_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_15_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_16_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_16_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_16_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_16_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_16_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_17_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_17_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_17_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_17_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_18_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_18_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_18_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_18_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_18_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_19_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_19_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_19_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_19_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_1_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_1_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_20_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_20_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_20_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_20_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_20_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_21_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_21_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_21_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_21_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_22_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_22_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_22_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_22_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_22_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_22_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_23_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_23_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_23_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_23_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_24_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_24_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_24_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_24_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_24_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_25_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_25_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_25_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_25_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_26_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_26_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_26_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_26_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_26_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_27_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_27_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_27_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_27_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_28_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_28_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_28_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_28_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_28_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_28_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_29_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_29_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_29_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_29_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_2_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_2_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_2_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_2_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_2_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_30_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_30_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_30_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_38 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_50 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_62 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_30_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_30_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_30_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_31_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_31_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_31_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_31_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_32_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_32_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_32_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_32_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_32 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_44 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_56 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_68 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_32_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_32_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_33_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_33_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_33_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_33_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_34_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_34_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_34_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_34_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_34_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_34_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_35_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_35_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_35_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_35_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_61 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_73 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_35_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_36_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_36_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_36_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_36_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_36_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_36_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_36_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_36_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_36_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_37_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_37_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_60 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_37_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_72 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_84 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_37_96 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_38_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_38_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_38_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_38_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_38_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_38_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_39_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_39_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_39_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_39_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_39_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_3_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_3_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_3_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_40_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_40_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_40_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_40_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_54 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_66 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_40_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_40_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_41_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_41_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_41_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_41_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_42_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_42_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_42_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_42_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_42 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_54 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_66 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_42_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_42_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_43_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_43_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_43_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_36 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_43_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_43_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_44_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_44_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_44_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_44_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_44_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_44_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_44_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_44_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_44_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_44_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_33 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_45 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_44_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_44_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_45_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_45_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_35 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_45_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_45_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_45_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_46_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_46_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_46_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_46_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_46_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_46_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_47_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_47_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_35 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_47_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_47_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_47_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_48_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_48_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_48_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_48_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_48_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_48_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_49_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_49_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_49_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_49_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_4_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_4_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_4_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_4_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_4_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_50_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_50_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_50_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_50_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_50_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_51_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_51_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_51_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_51_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_52_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_52_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_52_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_52_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_52_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_53_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_53_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_53_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_53_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_54_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_54_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_54_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_54_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_54_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_55_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_55_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_55_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_55_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_56_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_56_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_56_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_56_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_56_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_57_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_57_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_57_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_6 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 FILLER_57_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_57_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_11 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_23 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_5_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_5_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_35 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_5_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_5_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_5_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_6_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_6_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_6_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_6_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_6_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_7_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_7_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_7_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_7_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_109 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_121 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_141 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_153 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_165 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_177 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_197 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_209 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_221 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_233 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_253 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_265 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_277 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_8 FILLER_8_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_29 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__fill_2 FILLER_8_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_41 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_53 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_65 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_8_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_8_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_85 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_8_97 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_113 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_125 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_137 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_149 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_15 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_169 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_181 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_193 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_205 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_225 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_237 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_249 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_261 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_27 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_281 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_6 FILLER_9_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_3 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_39 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_4 FILLER_9_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_9_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_57 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_69 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_81 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_ef_sc_hd__decap_12 FILLER_9_93 (.VGND(vssd1),
    .VPWR(vccd1),
    .VPB(vccd1),
    .VNB(vssd1));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__mux2_2 _05_ (.A0(net1),
    .A1(\clknet_1_0__leaf_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ),
    .S(clknet_1_0__leaf_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_00_));
 sky130_fd_sc_hd__buf_1 _06_ (.A(_00_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ));
 sky130_fd_sc_hd__buf_1 _07_ (.A(clknet_1_1__leaf_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_01_));
 sky130_fd_sc_hd__nand2_2 _08_ (.A(clknet_1_0__leaf__01_),
    .B(\clknet_1_1__leaf_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_02_));
 sky130_fd_sc_hd__o21a_2 _09_ (.A1(clknet_1_0__leaf__01_),
    .A2(\clknet_1_1__leaf_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ),
    .B1(clknet_1_1__leaf__02_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__nand2_2 _10_ (.A(\clknet_1_0__leaf_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ),
    .B(clknet_1_0__leaf__02_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.out_0 ));
 sky130_fd_sc_hd__mux2_2 _11_ (.A0(net1),
    .A1(\clknet_1_0__leaf_SavedGate_1.LogicGate_0.in_0 ),
    .S(clknet_1_0__leaf_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_03_));
 sky130_fd_sc_hd__buf_1 _12_ (.A(_03_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SavedGate_1.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__nand2_2 _13_ (.A(clknet_1_0__leaf__01_),
    .B(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_04_));
 sky130_fd_sc_hd__o21a_2 _14_ (.A1(clknet_1_1__leaf__01_),
    .A2(\clknet_1_0__leaf_SavedGate_2.SavedGate_0.LogicGate_0.in_0 ),
    .B1(clknet_1_0__leaf__04_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SavedGate_2.SavedGate_0.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__nand2_2 _15_ (.A(\clknet_1_0__leaf_SavedGate_2.SavedGate_0.LogicGate_0.in_0 ),
    .B(clknet_1_1__leaf__04_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\SavedGate_2.SavedGate_0.LogicGate_0.out_0 ));
 sky130_fd_sc_hd__nand2_2 _16_ (.A(clknet_1_1__leaf__01_),
    .B(\clknet_1_0__leaf_SavedGate_4.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\SavedGate_4.LogicGate_0.out_0 ));
 sky130_fd_sc_hd__nand2_2 _17_ (.A(net1),
    .B(\clknet_1_0__leaf_SavedGate_4.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\SavedGate_4.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__buf_2 _19_ (.A(\clknet_1_1__leaf_SavedGate_1.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 _20_ (.A(\SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_2 _21_ (.A(\clknet_1_0__leaf_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_2 _22_ (.A(\SavedGate_2.SavedGate_0.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_2 _23_ (.A(\clknet_1_1__leaf_SavedGate_2.SavedGate_0.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_2 _24_ (.A(\clknet_1_1__leaf_SavedGate_4.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_2 _25_ (.A(\clknet_1_1__leaf_SavedGate_4.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(io_out[6]));
 sky130_fd_sc_hd__conb_1 c_tt2_mrcs_test_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net2));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0  (.A(\SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_0_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0  (.A(\SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_0_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_SavedGate_1.LogicGate_0.in_0  (.A(\SavedGate_1.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_0_SavedGate_1.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_SavedGate_2.SavedGate_0.LogicGate_0.in_0  (.A(\SavedGate_2.SavedGate_0.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_0_SavedGate_2.SavedGate_0.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_SavedGate_4.LogicGate_0.in_0  (.A(\SavedGate_4.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_0_SavedGate_4.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_SavedGate_4.LogicGate_0.out_0  (.A(\SavedGate_4.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_0_SavedGate_4.LogicGate_0.out_0 ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__01_ (.A(_01_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0__01_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__02_ (.A(_02_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0__02_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04_ (.A(_04_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0__04_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_io_in[0]  (.A(io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_0_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0  (.A(\clknet_0_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_0__leaf_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0  (.A(\clknet_0_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_0__leaf_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_SavedGate_1.LogicGate_0.in_0  (.A(\clknet_0_SavedGate_1.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_0__leaf_SavedGate_1.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_SavedGate_2.SavedGate_0.LogicGate_0.in_0  (.A(\clknet_0_SavedGate_2.SavedGate_0.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_0__leaf_SavedGate_2.SavedGate_0.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_SavedGate_4.LogicGate_0.in_0  (.A(\clknet_0_SavedGate_4.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_0__leaf_SavedGate_4.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_SavedGate_4.LogicGate_0.out_0  (.A(\clknet_0_SavedGate_4.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_0__leaf_SavedGate_4.LogicGate_0.out_0 ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__01_ (.A(clknet_0__01_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_0__leaf__01_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__02_ (.A(clknet_0__02_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_0__leaf__02_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04_ (.A(clknet_0__04_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_0__leaf__04_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_0__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0  (.A(\clknet_0_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_1__leaf_SavedGate_0.SavedGate_0.SavedGate_0.LogicGate_0.out_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0  (.A(\clknet_0_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_1__leaf_SavedGate_0.SavedGate_1.SavedGate_0.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_SavedGate_1.LogicGate_0.in_0  (.A(\clknet_0_SavedGate_1.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_1__leaf_SavedGate_1.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_SavedGate_2.SavedGate_0.LogicGate_0.in_0  (.A(\clknet_0_SavedGate_2.SavedGate_0.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_1__leaf_SavedGate_2.SavedGate_0.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_SavedGate_4.LogicGate_0.in_0  (.A(\clknet_0_SavedGate_4.LogicGate_0.in_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_1__leaf_SavedGate_4.LogicGate_0.in_0 ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_SavedGate_4.LogicGate_0.out_0  (.A(\clknet_0_SavedGate_4.LogicGate_0.out_0 ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\clknet_1_1__leaf_SavedGate_4.LogicGate_0.out_0 ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__01_ (.A(clknet_0__01_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_1__leaf__01_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__02_ (.A(clknet_0__02_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_1__leaf__02_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04_ (.A(clknet_0__04_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_1__leaf__04_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_io_in[0]  (.A(clknet_0_io_in[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(clknet_1_1__leaf_io_in[0]));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_in[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1));
 assign io_out[7] = net2;
endmodule
