VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO chase_the_beat
  CLASS BLOCK ;
  FOREIGN chase_the_beat ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 120.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 2.000 4.040 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.000 11.520 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.000 19.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.000 26.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.000 33.960 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.000 41.440 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.000 48.920 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.000 56.400 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 2.000 63.880 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 2.000 71.360 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.000 78.840 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.000 86.320 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.000 93.800 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.000 101.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 2.000 108.760 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.000 116.240 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.590 5.200 16.190 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.330 5.200 35.930 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.070 5.200 55.670 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.810 5.200 75.410 114.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.460 5.200 26.060 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.200 5.200 45.800 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.940 5.200 65.540 114.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 84.180 114.325 ;
      LAYER met1 ;
        RECT 5.520 5.200 84.180 114.480 ;
      LAYER met2 ;
        RECT 6.530 3.555 78.570 116.125 ;
      LAYER met3 ;
        RECT 2.400 115.240 78.595 116.105 ;
        RECT 2.000 109.160 78.595 115.240 ;
        RECT 2.400 107.760 78.595 109.160 ;
        RECT 2.000 101.680 78.595 107.760 ;
        RECT 2.400 100.280 78.595 101.680 ;
        RECT 2.000 94.200 78.595 100.280 ;
        RECT 2.400 92.800 78.595 94.200 ;
        RECT 2.000 86.720 78.595 92.800 ;
        RECT 2.400 85.320 78.595 86.720 ;
        RECT 2.000 79.240 78.595 85.320 ;
        RECT 2.400 77.840 78.595 79.240 ;
        RECT 2.000 71.760 78.595 77.840 ;
        RECT 2.400 70.360 78.595 71.760 ;
        RECT 2.000 64.280 78.595 70.360 ;
        RECT 2.400 62.880 78.595 64.280 ;
        RECT 2.000 56.800 78.595 62.880 ;
        RECT 2.400 55.400 78.595 56.800 ;
        RECT 2.000 49.320 78.595 55.400 ;
        RECT 2.400 47.920 78.595 49.320 ;
        RECT 2.000 41.840 78.595 47.920 ;
        RECT 2.400 40.440 78.595 41.840 ;
        RECT 2.000 34.360 78.595 40.440 ;
        RECT 2.400 32.960 78.595 34.360 ;
        RECT 2.000 26.880 78.595 32.960 ;
        RECT 2.400 25.480 78.595 26.880 ;
        RECT 2.000 19.400 78.595 25.480 ;
        RECT 2.400 18.000 78.595 19.400 ;
        RECT 2.000 11.920 78.595 18.000 ;
        RECT 2.400 10.520 78.595 11.920 ;
        RECT 2.000 4.440 78.595 10.520 ;
        RECT 2.400 3.575 78.595 4.440 ;
      LAYER met4 ;
        RECT 16.855 17.855 24.060 88.225 ;
        RECT 26.460 17.855 33.930 88.225 ;
        RECT 36.330 17.855 43.800 88.225 ;
        RECT 46.200 17.855 53.670 88.225 ;
        RECT 56.070 17.855 63.540 88.225 ;
        RECT 65.940 17.855 68.705 88.225 ;
  END
END chase_the_beat
END LIBRARY

