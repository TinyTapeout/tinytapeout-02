/* Automatically generated from https://wokwi.com/projects/349953952950780498 */

`default_nettype none

module user_module_349953952950780498(
  input [7:0] io_in,
  output [7:0] io_out
);
  wire net1 = io_in[0];
  wire net2 = io_in[1];
  wire net3 = io_in[2];
  wire net4 = io_in[3];
  wire net5 = io_in[4];
  wire net6 = io_in[5];
  wire net7 = io_in[6];
  wire net8 = io_in[7];
  wire net9;
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16;
  wire net17 = 1'b1;
  wire net18 = 1'b1;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24 = 1'b0;
  wire net25;
  wire net26 = 1'b0;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35 = 1'b0;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41 = 1'b0;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48 = 1'b0;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53 = 1'b0;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60 = 1'b0;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66 = 1'b0;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71 = 1'b0;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78 = 1'b0;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83 = 1'b0;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90 = 1'b0;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131 = 1'b0;
  wire net132;
  wire net133 = 1'b0;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205 = 1'b0;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247 = 1'b0;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284;
  wire net285;
  wire net286;
  wire net287;
  wire net288;
  wire net289;
  wire net290;
  wire net291;
  wire net292;
  wire net293;
  wire net294;
  wire net295;
  wire net296;
  wire net297;
  wire net298;
  wire net299;
  wire net300;
  wire net301;
  wire net302;
  wire net303 = 1'b0;
  wire net304;
  wire net305;
  wire net306;
  wire net307;
  wire net308;
  wire net309;
  wire net310;
  wire net311;
  wire net312;
  wire net313;
  wire net314;
  wire net315;
  wire net316;
  wire net317;
  wire net318;
  wire net319;
  wire net320;
  wire net321;
  wire net322;
  wire net323;
  wire net324;
  wire net325;
  wire net326;
  wire net327;
  wire net328;
  wire net329;
  wire net330;
  wire net331;
  wire net332;
  wire net333;
  wire net334;
  wire net335;
  wire net336;
  wire net337;
  wire net338;
  wire net339;
  wire net340;
  wire net341;
  wire net342;
  wire net343;
  wire net344;
  wire net345;
  wire net346;
  wire net347;
  wire net348;
  wire net349;
  wire net350;
  wire net351;
  wire net352;
  wire net353;
  wire net354;
  wire net355;
  wire net356;
  wire net357;
  wire net358;
  wire net359;
  wire net360;
  wire net361;
  wire net362;
  wire net363;
  wire net364;
  wire net365;
  wire net366;
  wire net367;
  wire net368;
  wire net369;

  assign io_out[0] = net9;
  assign io_out[1] = net10;
  assign io_out[2] = net11;
  assign io_out[3] = net12;
  assign io_out[4] = net13;
  assign io_out[5] = net14;
  assign io_out[6] = net15;
  assign io_out[7] = net16;

  dff_cell flipflop2 (
    .d (net19),
    .clk (net1),
    .q (net20)
  );
  dff_cell flipflop3 (
    .d (net21),
    .clk (net1),
    .q (net22)
  );
  buffer_cell gate12 (
    .in (net7)
  );
  mux_cell mux2 (
    .a (net23),
    .b (net24),
    .sel (net22),
    .out (net25)
  );
  mux_cell mux3 (
    .a (net20),
    .b (net26),
    .sel (net22),
    .out (net27)
  );
  and_cell gate13 (
    .a (net22),
    .b (net28)
  );
  and_cell gate14 (
    .a (net29),
    .b (net20),
    .out (net30)
  );
  not_cell gate17 (
    .in (net22),
    .out (net29)
  );
  dff_cell flipflop4 (
    .d (net31),
    .clk (net1),
    .q (net32)
  );
  buffer_cell gate19 (
    .in (net33),
    .out (net34)
  );
  mux_cell mux4 (
    .a (net35),
    .b (net34),
    .sel (net36),
    .out (net31)
  );
  dff_cell flipflop5 (
    .d (net37),
    .clk (net1),
    .q (net38)
  );
  buffer_cell gate22 (
    .in (net39),
    .out (net40)
  );
  mux_cell mux5 (
    .a (net41),
    .b (net40),
    .sel (net36),
    .out (net37)
  );
  buffer_cell gate24 (
    .in (net32),
    .out (net42)
  );
  buffer_cell gate25 (
    .in (net38),
    .out (net43)
  );
  dff_cell flipflop6 (
    .d (net44),
    .clk (net1),
    .q (net45)
  );
  buffer_cell gate26 (
    .in (net46),
    .out (net47)
  );
  mux_cell mux6 (
    .a (net48),
    .b (net47),
    .sel (net36),
    .out (net44)
  );
  dff_cell flipflop7 (
    .d (net49),
    .clk (net1),
    .q (net50)
  );
  buffer_cell gate28 (
    .in (net51),
    .out (net52)
  );
  mux_cell mux7 (
    .a (net53),
    .b (net52),
    .sel (net36),
    .out (net49)
  );
  buffer_cell gate30 (
    .in (net45),
    .out (net54)
  );
  buffer_cell gate31 (
    .in (net50),
    .out (net55)
  );
  dff_cell flipflop9 (
    .d (net56),
    .clk (net1),
    .q (net57)
  );
  buffer_cell gate32 (
    .in (net58),
    .out (net59)
  );
  mux_cell mux8 (
    .a (net60),
    .b (net59),
    .sel (net36),
    .out (net56)
  );
  buffer_cell gate34 (
    .in (net57),
    .out (net61)
  );
  dff_cell flipflop8 (
    .d (net62),
    .clk (net1),
    .q (net63)
  );
  buffer_cell gate35 (
    .in (net64),
    .out (net65)
  );
  mux_cell mux9 (
    .a (net66),
    .b (net65),
    .sel (net30),
    .out (net62)
  );
  dff_cell flipflop10 (
    .d (net67),
    .clk (net1),
    .q (net68)
  );
  buffer_cell gate37 (
    .in (net69),
    .out (net70)
  );
  mux_cell mux10 (
    .a (net71),
    .b (net70),
    .sel (net30),
    .out (net67)
  );
  buffer_cell gate39 (
    .in (net63),
    .out (net72)
  );
  buffer_cell gate40 (
    .in (net68),
    .out (net73)
  );
  dff_cell flipflop11 (
    .d (net74),
    .clk (net1),
    .q (net75)
  );
  buffer_cell gate41 (
    .in (net76),
    .out (net77)
  );
  mux_cell mux11 (
    .a (net78),
    .b (net77),
    .sel (net30),
    .out (net74)
  );
  dff_cell flipflop12 (
    .d (net79),
    .clk (net1),
    .q (net80)
  );
  buffer_cell gate43 (
    .in (net81),
    .out (net82)
  );
  mux_cell mux12 (
    .a (net83),
    .b (net82),
    .sel (net30),
    .out (net79)
  );
  buffer_cell gate45 (
    .in (net75),
    .out (net84)
  );
  buffer_cell gate46 (
    .in (net80),
    .out (net85)
  );
  dff_cell flipflop13 (
    .d (net86),
    .clk (net1),
    .q (net87)
  );
  buffer_cell gate47 (
    .in (net88),
    .out (net89)
  );
  mux_cell mux13 (
    .a (net90),
    .b (net89),
    .sel (net30),
    .out (net86)
  );
  buffer_cell gate49 (
    .in (net87),
    .out (net91)
  );
  not_cell gate51 (
    .in (net92),
    .out (net36)
  );
  or_cell gate52 (
    .a (net22),
    .b (net20),
    .out (net92)
  );
  dff_cell flipflop14 (
    .d (net93),
    .clk (net1),
    .q (net94)
  );
  buffer_cell gate15 (
    .in (net95),
    .out (net96)
  );
  mux_cell mux14 (
    .a (net94),
    .b (net96),
    .sel (net30),
    .out (net93)
  );
  buffer_cell gate16 (
    .in (net94),
    .out (net97)
  );
  dff_cell flipflop15 (
    .d (net98),
    .clk (net1),
    .q (net99)
  );
  buffer_cell gate18 (
    .in (net100),
    .out (net101)
  );
  mux_cell mux15 (
    .a (net99),
    .b (net101),
    .sel (net30),
    .out (net98)
  );
  buffer_cell gate20 (
    .in (net99),
    .out (net102)
  );
  dff_cell flipflop16 (
    .d (net103),
    .clk (net1),
    .q (net104)
  );
  buffer_cell gate23 (
    .in (net105),
    .out (net106)
  );
  mux_cell mux16 (
    .a (net104),
    .b (net106),
    .sel (net30),
    .out (net103)
  );
  buffer_cell gate27 (
    .in (net104),
    .out (net107)
  );
  dff_cell flipflop17 (
    .d (net108),
    .clk (net1),
    .q (net109)
  );
  buffer_cell gate29 (
    .in (net110),
    .out (net111)
  );
  mux_cell mux17 (
    .a (net109),
    .b (net111),
    .sel (net30),
    .out (net108)
  );
  buffer_cell gate36 (
    .in (net109),
    .out (net112)
  );
  dff_cell flipflop18 (
    .d (net113),
    .clk (net1),
    .q (net114)
  );
  buffer_cell gate38 (
    .in (net115),
    .out (net116)
  );
  mux_cell mux18 (
    .a (net114),
    .b (net116),
    .sel (net30),
    .out (net113)
  );
  buffer_cell gate42 (
    .in (net114),
    .out (net117)
  );
  dff_cell flipflop19 (
    .d (net118),
    .clk (net1),
    .q (net119)
  );
  buffer_cell gate44 (
    .in (net120),
    .out (net121)
  );
  mux_cell mux19 (
    .a (net119),
    .b (net121),
    .sel (net30),
    .out (net118)
  );
  buffer_cell gate48 (
    .in (net119),
    .out (net122)
  );
  and_cell gate62 (
    .a (net123),
    .b (net36),
    .out (net33)
  );
  and_cell gate63 (
    .a (net124),
    .b (net36),
    .out (net39)
  );
  and_cell gate64 (
    .a (net125),
    .b (net36),
    .out (net46)
  );
  and_cell gate66 (
    .a (net126),
    .b (net36),
    .out (net58)
  );
  and_cell gate67 (
    .a (net127),
    .b (net36),
    .out (net51)
  );
  and_cell gate65 (
    .a (net123),
    .b (net30),
    .out (net64)
  );
  and_cell gate68 (
    .a (net124),
    .b (net30),
    .out (net69)
  );
  and_cell gate69 (
    .a (net125),
    .b (net30),
    .out (net76)
  );
  and_cell gate70 (
    .a (net126),
    .b (net30),
    .out (net88)
  );
  and_cell gate71 (
    .a (net127),
    .b (net30),
    .out (net81)
  );
  buffer_cell gate72 (
    .in (net2),
    .out (net123)
  );
  buffer_cell gate73 (
    .in (net3),
    .out (net124)
  );
  buffer_cell gate74 (
    .in (net4),
    .out (net125)
  );
  buffer_cell gate75 (
    .in (net5),
    .out (net127)
  );
  buffer_cell gate76 (
    .in (net6),
    .out (net126)
  );
  buffer_cell gate78 (
    .in (net8),
    .out (net128)
  );
  and_cell gate79 (
    .a (net2),
    .b (net129),
    .out (net130)
  );
  mux_cell mux20 (
    .a (net131),
    .b (net107),
    .sel (net128),
    .out (net132)
  );
  mux_cell mux21 (
    .a (net133),
    .b (net112),
    .sel (net128),
    .out (net134)
  );
  mux_cell mux22 (
    .a (net97),
    .b (net117),
    .sel (net128),
    .out (net135)
  );
  mux_cell mux23 (
    .a (net102),
    .b (net122),
    .sel (net128),
    .out (net136)
  );
  buffer_cell gate33 (
    .in (net132),
    .out (net137)
  );
  buffer_cell gate50 (
    .in (net134),
    .out (net138)
  );
  buffer_cell gate53 (
    .in (net136),
    .out (net139)
  );
  buffer_cell gate54 (
    .in (net135),
    .out (net140)
  );
  not_cell gate55 (
    .in (net139),
    .out (net141)
  );
  not_cell gate56 (
    .in (net140),
    .out (net142)
  );
  not_cell gate57 (
    .in (net138),
    .out (net143)
  );
  not_cell gate58 (
    .in (net137),
    .out (net144)
  );
  and_cell gate61 (
    .a (net139),
    .b (net145),
    .out (net146)
  );
  and_cell gate77 (
    .a (net144),
    .b (net138),
    .out (net145)
  );
  or_cell gate80 (
    .a (net147),
    .b (net148),
    .out (net9)
  );
  and_cell gate81 (
    .a (net137),
    .b (net141),
    .out (net149)
  );
  and_cell gate82 (
    .a (net142),
    .b (net150),
    .out (net151)
  );
  and_cell gate138 (
    .a (net143),
    .b (net137),
    .out (net150)
  );
  and_cell gate139 (
    .a (net140),
    .b (net144),
    .out (net152)
  );
  and_cell gate140 (
    .a (net138),
    .b (net140),
    .out (net153)
  );
  or_cell gate141 (
    .a (net154),
    .b (net153),
    .out (net155)
  );
  or_cell gate142 (
    .a (net152),
    .b (net146),
    .out (net156)
  );
  or_cell gate143 (
    .a (net151),
    .b (net149),
    .out (net148)
  );
  or_cell gate144 (
    .a (net155),
    .b (net156),
    .out (net147)
  );
  and_cell gate145 (
    .a (net137),
    .b (net157),
    .out (net158)
  );
  and_cell gate146 (
    .a (net142),
    .b (net139),
    .out (net157)
  );
  and_cell gate147 (
    .a (net143),
    .b (net141),
    .out (net154)
  );
  and_cell gate148 (
    .a (net144),
    .b (net159),
    .out (net160)
  );
  and_cell gate149 (
    .a (net142),
    .b (net141),
    .out (net159)
  );
  and_cell gate150 (
    .a (net144),
    .b (net140),
    .out (net161)
  );
  and_cell gate151 (
    .a (net161),
    .b (net139),
    .out (net162)
  );
  and_cell gate152 (
    .a (net144),
    .b (net143),
    .out (net163)
  );
  or_cell gate153 (
    .a (net158),
    .b (net163),
    .out (net164)
  );
  or_cell gate154 (
    .a (net162),
    .b (net160),
    .out (net165)
  );
  or_cell gate155 (
    .a (net164),
    .b (net165),
    .out (net166)
  );
  or_cell gate156 (
    .a (net166),
    .b (net154),
    .out (net10)
  );
  and_cell gate157 (
    .a (net137),
    .b (net143),
    .out (net167)
  );
  and_cell gate158 (
    .a (net144),
    .b (net138),
    .out (net168)
  );
  and_cell gate159 (
    .a (net144),
    .b (net142),
    .out (net169)
  );
  and_cell gate160 (
    .a (net144),
    .b (net139),
    .out (net170)
  );
  and_cell gate161 (
    .a (net139),
    .b (net142),
    .out (net171)
  );
  or_cell gate162 (
    .a (net167),
    .b (net168),
    .out (net172)
  );
  or_cell gate163 (
    .a (net169),
    .b (net170),
    .out (net173)
  );
  or_cell gate164 (
    .a (net172),
    .b (net173),
    .out (net174)
  );
  or_cell gate165 (
    .a (net174),
    .b (net171),
    .out (net11)
  );
  and_cell gate166 (
    .a (net138),
    .b (net142),
    .out (net175)
  );
  and_cell gate167 (
    .a (net144),
    .b (net140),
    .out (net176)
  );
  and_cell gate168 (
    .a (net137),
    .b (net138),
    .out (net177)
  );
  and_cell gate169 (
    .a (net175),
    .b (net139),
    .out (net178)
  );
  and_cell gate170 (
    .a (net176),
    .b (net141),
    .out (net179)
  );
  and_cell gate171 (
    .a (net177),
    .b (net141),
    .out (net180)
  );
  and_cell gate172 (
    .a (net143),
    .b (net142),
    .out (net181)
  );
  and_cell gate173 (
    .a (net143),
    .b (net140),
    .out (net182)
  );
  and_cell gate174 (
    .a (net181),
    .b (net141),
    .out (net183)
  );
  and_cell gate175 (
    .a (net182),
    .b (net139),
    .out (net184)
  );
  or_cell gate176 (
    .a (net180),
    .b (net179),
    .out (net185)
  );
  or_cell gate177 (
    .a (net178),
    .b (net184),
    .out (net186)
  );
  or_cell gate178 (
    .a (net185),
    .b (net186),
    .out (net187)
  );
  or_cell gate179 (
    .a (net187),
    .b (net183),
    .out (net12)
  );
  and_cell gate180 (
    .a (net137),
    .b (net140),
    .out (net188)
  );
  and_cell gate181 (
    .a (net137),
    .b (net138),
    .out (net189)
  );
  and_cell gate182 (
    .a (net140),
    .b (net141),
    .out (net190)
  );
  or_cell gate183 (
    .a (net189),
    .b (net188),
    .out (net191)
  );
  or_cell gate184 (
    .a (net154),
    .b (net190),
    .out (net192)
  );
  or_cell gate185 (
    .a (net191),
    .b (net192),
    .out (net13)
  );
  and_cell gate186 (
    .a (net137),
    .b (net143),
    .out (net193)
  );
  and_cell gate187 (
    .a (net169),
    .b (net138),
    .out (net194)
  );
  and_cell gate188 (
    .a (net138),
    .b (net141),
    .out (net195)
  );
  or_cell gate189 (
    .a (net193),
    .b (net188),
    .out (net196)
  );
  or_cell gate190 (
    .a (net194),
    .b (net195),
    .out (net197)
  );
  or_cell gate191 (
    .a (net196),
    .b (net197),
    .out (net198)
  );
  or_cell gate192 (
    .a (net198),
    .b (net159),
    .out (net14)
  );
  and_cell gate193 (
    .a (net193),
    .b (net199),
    .out (net16)
  );
  and_cell gate194 (
    .a (net137),
    .b (net139),
    .out (net200)
  );
  or_cell gate195 (
    .a (net193),
    .b (net194),
    .out (net201)
  );
  or_cell gate196 (
    .a (net200),
    .b (net202),
    .out (net203)
  );
  and_cell gate197 (
    .a (net143),
    .b (net140),
    .out (net202)
  );
  or_cell gate198 (
    .a (net201),
    .b (net203),
    .out (net204)
  );
  or_cell gate199 (
    .a (net190),
    .b (net204),
    .out (net15)
  );
  and_cell gate200 (
    .a (net140),
    .b (net139),
    .out (net199)
  );
  buffer_cell gate60 (
    .in (net206),
    .out (net207)
  );
  buffer_cell gate83 (
    .in (net208),
    .out (net209)
  );
  buffer_cell gate84 (
    .in (net210),
    .out (net211)
  );
  xor_cell gate85 (
    .a (net211),
    .b (net207),
    .out (net212)
  );
  xor_cell gate86 (
    .a (net209),
    .b (net212),
    .out (net213)
  );
  and_cell gate87 (
    .a (net209),
    .b (net207),
    .out (net214)
  );
  and_cell gate88 (
    .a (net209),
    .b (net211),
    .out (net215)
  );
  and_cell gate89 (
    .a (net211),
    .b (net207),
    .out (net216)
  );
  or_cell gate90 (
    .a (net215),
    .b (net214),
    .out (net217)
  );
  or_cell gate91 (
    .a (net216),
    .b (net217),
    .out (net218)
  );
  buffer_cell gate92 (
    .in (net219),
    .out (net220)
  );
  buffer_cell gate93 (
    .in (net221),
    .out (net222)
  );
  buffer_cell gate94 (
    .in (net223),
    .out (net224)
  );
  xor_cell gate95 (
    .a (net224),
    .b (net220),
    .out (net225)
  );
  xor_cell gate96 (
    .a (net222),
    .b (net225),
    .out (net226)
  );
  and_cell gate97 (
    .a (net222),
    .b (net220),
    .out (net227)
  );
  and_cell gate98 (
    .a (net222),
    .b (net224),
    .out (net228)
  );
  and_cell gate99 (
    .a (net224),
    .b (net220),
    .out (net229)
  );
  or_cell gate100 (
    .a (net228),
    .b (net227),
    .out (net230)
  );
  or_cell gate101 (
    .a (net229),
    .b (net230),
    .out (net231)
  );
  buffer_cell gate102 (
    .in (net232),
    .out (net233)
  );
  buffer_cell gate103 (
    .in (net234),
    .out (net235)
  );
  buffer_cell gate104 (
    .in (net231),
    .out (net236)
  );
  xor_cell gate105 (
    .a (net236),
    .b (net233),
    .out (net237)
  );
  xor_cell gate106 (
    .a (net235),
    .b (net237),
    .out (net238)
  );
  and_cell gate107 (
    .a (net235),
    .b (net233),
    .out (net239)
  );
  and_cell gate108 (
    .a (net235),
    .b (net236),
    .out (net240)
  );
  and_cell gate109 (
    .a (net236),
    .b (net233),
    .out (net241)
  );
  or_cell gate110 (
    .a (net240),
    .b (net239),
    .out (net242)
  );
  or_cell gate111 (
    .a (net241),
    .b (net242),
    .out (net210)
  );
  buffer_cell gate112 (
    .in (net243),
    .out (net244)
  );
  buffer_cell gate113 (
    .in (net245),
    .out (net246)
  );
  buffer_cell gate114 (
    .in (net247),
    .out (net248)
  );
  xor_cell gate115 (
    .a (net248),
    .b (net244),
    .out (net249)
  );
  xor_cell gate116 (
    .a (net246),
    .b (net249),
    .out (net250)
  );
  and_cell gate117 (
    .a (net246),
    .b (net244),
    .out (net251)
  );
  and_cell gate118 (
    .a (net246),
    .b (net248),
    .out (net252)
  );
  and_cell gate119 (
    .a (net248),
    .b (net244),
    .out (net253)
  );
  or_cell gate120 (
    .a (net252),
    .b (net251),
    .out (net254)
  );
  or_cell gate121 (
    .a (net253),
    .b (net254),
    .out (net255)
  );
  buffer_cell gate122 (
    .in (net256),
    .out (net257)
  );
  buffer_cell gate123 (
    .in (net258),
    .out (net259)
  );
  buffer_cell gate124 (
    .in (net255),
    .out (net260)
  );
  xor_cell gate125 (
    .a (net260),
    .b (net257),
    .out (net261)
  );
  xor_cell gate126 (
    .a (net259),
    .b (net261),
    .out (net262)
  );
  and_cell gate127 (
    .a (net259),
    .b (net257),
    .out (net263)
  );
  and_cell gate128 (
    .a (net259),
    .b (net260),
    .out (net264)
  );
  and_cell gate129 (
    .a (net260),
    .b (net257),
    .out (net265)
  );
  or_cell gate130 (
    .a (net264),
    .b (net263),
    .out (net266)
  );
  or_cell gate131 (
    .a (net265),
    .b (net266),
    .out (net223)
  );
  xor_cell gate132 (
    .a (net267),
    .b (net268),
    .out (net269)
  );
  xor_cell gate133 (
    .a (net270),
    .b (net269),
    .out (net271)
  );
  and_cell gate134 (
    .a (net272),
    .b (net267),
    .out (net273)
  );
  or_cell gate135 (
    .a (net274),
    .b (net273),
    .out (net275)
  );
  buffer_cell gate136 (
    .in (net276),
    .out (net270)
  );
  buffer_cell gate137 (
    .in (net277),
    .out (net268)
  );
  buffer_cell gate201 (
    .in (net278),
    .out (net267)
  );
  not_cell gate202 (
    .in (net268),
    .out (net272)
  );
  and_cell gate203 (
    .a (net279),
    .b (net270),
    .out (net274)
  );
  not_cell gate204 (
    .in (net269),
    .out (net279)
  );
  xor_cell gate205 (
    .a (net280),
    .b (net281),
    .out (net282)
  );
  xor_cell gate206 (
    .a (net283),
    .b (net282),
    .out (net284)
  );
  and_cell gate207 (
    .a (net285),
    .b (net280),
    .out (net286)
  );
  or_cell gate208 (
    .a (net287),
    .b (net286),
    .out (net288)
  );
  buffer_cell gate209 (
    .in (net289),
    .out (net283)
  );
  buffer_cell gate210 (
    .in (net290),
    .out (net281)
  );
  buffer_cell gate211 (
    .in (net275),
    .out (net280)
  );
  not_cell gate212 (
    .in (net281),
    .out (net285)
  );
  and_cell gate213 (
    .a (net291),
    .b (net283),
    .out (net287)
  );
  not_cell gate214 (
    .in (net282),
    .out (net291)
  );
  xor_cell gate215 (
    .a (net292),
    .b (net293),
    .out (net294)
  );
  xor_cell gate216 (
    .a (net295),
    .b (net294),
    .out (net296)
  );
  and_cell gate217 (
    .a (net297),
    .b (net292),
    .out (net298)
  );
  or_cell gate218 (
    .a (net299),
    .b (net298),
    .out (net300)
  );
  buffer_cell gate219 (
    .in (net301),
    .out (net295)
  );
  buffer_cell gate220 (
    .in (net302),
    .out (net293)
  );
  buffer_cell gate221 (
    .in (net303),
    .out (net292)
  );
  not_cell gate222 (
    .in (net293),
    .out (net297)
  );
  and_cell gate223 (
    .a (net304),
    .b (net295),
    .out (net299)
  );
  not_cell gate224 (
    .in (net294),
    .out (net304)
  );
  xor_cell gate225 (
    .a (net305),
    .b (net306),
    .out (net307)
  );
  xor_cell gate226 (
    .a (net308),
    .b (net307),
    .out (net309)
  );
  and_cell gate227 (
    .a (net310),
    .b (net305),
    .out (net311)
  );
  or_cell gate228 (
    .a (net312),
    .b (net311),
    .out (net278)
  );
  buffer_cell gate229 (
    .in (net313),
    .out (net308)
  );
  buffer_cell gate230 (
    .in (net314),
    .out (net306)
  );
  buffer_cell gate231 (
    .in (net300),
    .out (net305)
  );
  not_cell gate232 (
    .in (net306),
    .out (net310)
  );
  and_cell gate233 (
    .a (net315),
    .b (net308),
    .out (net312)
  );
  not_cell gate234 (
    .in (net307),
    .out (net315)
  );
  xor_cell gate235 (
    .a (net316),
    .b (net317),
    .out (net318)
  );
  xor_cell gate236 (
    .a (net319),
    .b (net318),
    .out (net320)
  );
  and_cell gate237 (
    .a (net321),
    .b (net316),
    .out (net322)
  );
  or_cell gate238 (
    .a (net323),
    .b (net322),
    .out (net324)
  );
  buffer_cell gate239 (
    .in (net325),
    .out (net319)
  );
  buffer_cell gate240 (
    .in (net326),
    .out (net317)
  );
  buffer_cell gate241 (
    .in (net288),
    .out (net316)
  );
  not_cell gate242 (
    .in (net317),
    .out (net321)
  );
  and_cell gate243 (
    .a (net327),
    .b (net319),
    .out (net323)
  );
  not_cell gate244 (
    .in (net318),
    .out (net327)
  );
  and_cell gate245 (
    .a (net328),
    .b (net329),
    .out (net208)
  );
  and_cell gate246 (
    .a (net330),
    .b (net331),
    .out (net206)
  );
  buffer_cell gate247 (
    .in (net61),
    .out (net329)
  );
  buffer_cell gate248 (
    .in (net130),
    .out (net328)
  );
  buffer_cell gate249 (
    .in (net130),
    .out (net331)
  );
  buffer_cell gate250 (
    .in (net91),
    .out (net330)
  );
  and_cell gate251 (
    .a (net332),
    .b (net333),
    .out (net234)
  );
  and_cell gate252 (
    .a (net334),
    .b (net335),
    .out (net232)
  );
  buffer_cell gate253 (
    .in (net55),
    .out (net333)
  );
  buffer_cell gate254 (
    .in (net328),
    .out (net332)
  );
  buffer_cell gate255 (
    .in (net328),
    .out (net335)
  );
  buffer_cell gate256 (
    .in (net85),
    .out (net334)
  );
  and_cell gate257 (
    .a (net336),
    .b (net337),
    .out (net221)
  );
  and_cell gate258 (
    .a (net338),
    .b (net339),
    .out (net219)
  );
  buffer_cell gate259 (
    .in (net54),
    .out (net337)
  );
  buffer_cell gate260 (
    .in (net332),
    .out (net336)
  );
  buffer_cell gate261 (
    .in (net332),
    .out (net339)
  );
  buffer_cell gate262 (
    .in (net84),
    .out (net338)
  );
  and_cell gate263 (
    .a (net340),
    .b (net341),
    .out (net258)
  );
  and_cell gate264 (
    .a (net342),
    .b (net343),
    .out (net256)
  );
  buffer_cell gate265 (
    .in (net43),
    .out (net341)
  );
  buffer_cell gate266 (
    .in (net343),
    .out (net340)
  );
  buffer_cell gate267 (
    .in (net336),
    .out (net343)
  );
  buffer_cell gate268 (
    .in (net73),
    .out (net342)
  );
  and_cell gate269 (
    .a (net344),
    .b (net345),
    .out (net245)
  );
  and_cell gate270 (
    .a (net346),
    .b (net347),
    .out (net243)
  );
  buffer_cell gate271 (
    .in (net42),
    .out (net345)
  );
  buffer_cell gate272 (
    .in (net347),
    .out (net344)
  );
  buffer_cell gate273 (
    .in (net340),
    .out (net347)
  );
  buffer_cell gate274 (
    .in (net72),
    .out (net346)
  );
  and_cell gate275 (
    .a (net348),
    .b (net349),
    .out (net325)
  );
  and_cell gate276 (
    .a (net350),
    .b (net351),
    .out (net326)
  );
  buffer_cell gate277 (
    .in (net61),
    .out (net349)
  );
  buffer_cell gate278 (
    .in (net91),
    .out (net350)
  );
  and_cell gate279 (
    .a (net352),
    .b (net353),
    .out (net289)
  );
  and_cell gate280 (
    .a (net354),
    .b (net355),
    .out (net290)
  );
  buffer_cell gate281 (
    .in (net55),
    .out (net353)
  );
  buffer_cell gate282 (
    .in (net85),
    .out (net354)
  );
  and_cell gate283 (
    .a (net356),
    .b (net357),
    .out (net276)
  );
  and_cell gate284 (
    .a (net358),
    .b (net359),
    .out (net277)
  );
  buffer_cell gate285 (
    .in (net54),
    .out (net357)
  );
  buffer_cell gate286 (
    .in (net84),
    .out (net358)
  );
  and_cell gate287 (
    .a (net360),
    .b (net361),
    .out (net313)
  );
  and_cell gate288 (
    .a (net362),
    .b (net363),
    .out (net314)
  );
  buffer_cell gate289 (
    .in (net43),
    .out (net361)
  );
  buffer_cell gate290 (
    .in (net73),
    .out (net362)
  );
  and_cell gate291 (
    .a (net364),
    .b (net365),
    .out (net301)
  );
  and_cell gate292 (
    .a (net366),
    .b (net367),
    .out (net302)
  );
  buffer_cell gate293 (
    .in (net42),
    .out (net365)
  );
  buffer_cell gate294 (
    .in (net72),
    .out (net366)
  );
  not_cell gate295 (
    .in (net130),
    .out (net348)
  );
  not_cell gate296 (
    .in (net130),
    .out (net351)
  );
  not_cell gate297 (
    .in (net328),
    .out (net352)
  );
  not_cell gate298 (
    .in (net328),
    .out (net355)
  );
  not_cell gate299 (
    .in (net332),
    .out (net356)
  );
  not_cell gate300 (
    .in (net332),
    .out (net359)
  );
  not_cell gate301 (
    .in (net343),
    .out (net360)
  );
  not_cell gate302 (
    .in (net336),
    .out (net363)
  );
  not_cell gate303 (
    .in (net347),
    .out (net364)
  );
  not_cell gate304 (
    .in (net340),
    .out (net367)
  );
  or_cell gate305 (
    .a (net213),
    .b (net320),
    .out (net100)
  );
  or_cell gate306 (
    .a (net284),
    .b (net238),
    .out (net105)
  );
  or_cell gate307 (
    .a (net271),
    .b (net226),
    .out (net110)
  );
  or_cell gate308 (
    .a (net309),
    .b (net262),
    .out (net115)
  );
  or_cell gate309 (
    .a (net296),
    .b (net250),
    .out (net120)
  );
  or_cell gate310 (
    .a (net324),
    .b (net218),
    .out (net95)
  );
  buffer_cell gate311 (
    .in (net7),
    .out (net368)
  );
  mux_cell mux24 (
    .a (net20),
    .b (net25),
    .sel (net368),
    .out (net19)
  );
  mux_cell mux25 (
    .a (net22),
    .b (net27),
    .sel (net368),
    .out (net21)
  );
  or_cell gate312 (
    .a (net30),
    .b (net36),
    .out (net129)
  );
  xor_cell gate5 (
    .a (net22),
    .b (net20),
    .out (net369)
  );
  not_cell gate7 (
    .in (net369),
    .out (net23)
  );
  not_cell gate8 (
    .in (net20),
    .out (net28)
  );
endmodule
