VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_module_341535056611770964
  CLASS BLOCK ;
  FOREIGN user_module_341535056611770964 ;
  ORIGIN 0.000 0.000 ;
  SIZE 160.000 BY 200.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 2.000 8.120 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 2.000 20.360 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 2.000 32.600 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 2.000 44.840 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.000 57.080 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 2.000 69.320 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 2.000 81.560 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.000 93.800 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 2.000 106.040 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 2.000 118.280 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 2.000 130.520 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 2.000 142.760 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 2.000 155.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 2.000 167.240 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 2.000 179.480 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 2.000 191.720 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.340 5.200 24.940 193.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.580 5.200 62.180 193.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.820 5.200 99.420 193.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 135.060 5.200 136.660 193.360 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 41.960 5.200 43.560 193.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.200 5.200 80.800 193.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.440 5.200 118.040 193.360 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 154.100 193.205 ;
      LAYER met1 ;
        RECT 5.520 5.200 154.100 193.360 ;
      LAYER met2 ;
        RECT 6.990 5.255 136.630 193.305 ;
      LAYER met3 ;
        RECT 2.000 192.120 136.650 193.285 ;
        RECT 2.400 190.720 136.650 192.120 ;
        RECT 2.000 179.880 136.650 190.720 ;
        RECT 2.400 178.480 136.650 179.880 ;
        RECT 2.000 167.640 136.650 178.480 ;
        RECT 2.400 166.240 136.650 167.640 ;
        RECT 2.000 155.400 136.650 166.240 ;
        RECT 2.400 154.000 136.650 155.400 ;
        RECT 2.000 143.160 136.650 154.000 ;
        RECT 2.400 141.760 136.650 143.160 ;
        RECT 2.000 130.920 136.650 141.760 ;
        RECT 2.400 129.520 136.650 130.920 ;
        RECT 2.000 118.680 136.650 129.520 ;
        RECT 2.400 117.280 136.650 118.680 ;
        RECT 2.000 106.440 136.650 117.280 ;
        RECT 2.400 105.040 136.650 106.440 ;
        RECT 2.000 94.200 136.650 105.040 ;
        RECT 2.400 92.800 136.650 94.200 ;
        RECT 2.000 81.960 136.650 92.800 ;
        RECT 2.400 80.560 136.650 81.960 ;
        RECT 2.000 69.720 136.650 80.560 ;
        RECT 2.400 68.320 136.650 69.720 ;
        RECT 2.000 57.480 136.650 68.320 ;
        RECT 2.400 56.080 136.650 57.480 ;
        RECT 2.000 45.240 136.650 56.080 ;
        RECT 2.400 43.840 136.650 45.240 ;
        RECT 2.000 33.000 136.650 43.840 ;
        RECT 2.400 31.600 136.650 33.000 ;
        RECT 2.000 20.760 136.650 31.600 ;
        RECT 2.400 19.360 136.650 20.760 ;
        RECT 2.000 8.520 136.650 19.360 ;
        RECT 2.400 7.120 136.650 8.520 ;
        RECT 2.000 5.275 136.650 7.120 ;
  END
END user_module_341535056611770964
END LIBRARY

