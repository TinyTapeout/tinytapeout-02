/* Automatically generated from https://wokwi.com/projects/347894637149553236 */

`default_nettype none

module user_module_347894637149553236(
  input [7:0] io_in,
  output [7:0] io_out
);
  wire net1 = io_in[0];
  wire net2 = io_in[1];
  wire net3 = io_in[2];
  wire net4 = io_in[3];
  wire net5 = io_in[4];
  wire net6 = io_in[5];
  wire net7 = io_in[6];
  wire net8 = io_in[7];
  wire net9;
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16;
  wire net17;
  wire net18;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36 = 1'b0;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117 = 1'b0;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247 = 1'b0;
  wire net248 = 1'b1;
  wire net249 = 1'b0;
  wire net250 = 1'b0;
  wire net251 = 1'b0;
  wire net252;
  wire net253;
  wire net254 = 1'b0;
  wire net255 = 1'b0;
  wire net256;
  wire net257 = 1'b0;
  wire net258 = 1'b0;

  assign io_out[0] = net9;
  assign io_out[1] = net10;
  assign io_out[2] = net11;
  assign io_out[3] = net12;
  assign io_out[4] = net13;
  assign io_out[5] = net14;
  assign io_out[6] = net15;
  assign io_out[7] = net16;

  xor_cell xor1 (
    .a (net17),
    .b (net18),
    .out (net19)
  );
  and_cell and1 (
    .a (net17),
    .b (net18),
    .out (net20)
  );
  xor_cell xor2 (
    .a (net21),
    .b (net22),
    .out (net23)
  );
  xor_cell xor3 (
    .a (net20),
    .b (net23),
    .out (net24)
  );
  and_cell and2 (
    .a (net21),
    .b (net22),
    .out (net25)
  );
  and_cell and3 (
    .a (net20),
    .b (net23),
    .out (net26)
  );
  or_cell or1 (
    .a (net26),
    .b (net25),
    .out (net27)
  );
  xor_cell xor4 (
    .a (net28),
    .b (net29),
    .out (net30)
  );
  xor_cell xor5 (
    .a (net27),
    .b (net30),
    .out (net31)
  );
  and_cell and5 (
    .a (net28),
    .b (net29),
    .out (net32)
  );
  and_cell and6 (
    .a (net27),
    .b (net30),
    .out (net33)
  );
  or_cell or2 (
    .a (net33),
    .b (net32),
    .out (net34)
  );
  xor_cell xor6 (
    .a (net35),
    .b (net36),
    .out (net37)
  );
  xor_cell xor7 (
    .a (net34),
    .b (net37),
    .out (net38)
  );
  and_cell and4 (
    .a (net35),
    .b (net36),
    .out (net39)
  );
  and_cell and7 (
    .a (net34),
    .b (net37),
    .out (net40)
  );
  or_cell or3 (
    .a (net40),
    .b (net39),
    .out (net41)
  );
  and_cell and8 (
    .a (net42),
    .b (net43),
    .out (net44)
  );
  and_cell and9 (
    .a (net45),
    .b (net43),
    .out (net18)
  );
  and_cell and10 (
    .a (net46),
    .b (net43),
    .out (net22)
  );
  and_cell and11 (
    .a (net47),
    .b (net43),
    .out (net29)
  );
  dff_cell flop4 (
    .d (net48),
    .clk (net49),
    .q (net47)
  );
  dff_cell flop1 (
    .d (net50),
    .clk (net49),
    .q (net46)
  );
  dff_cell flop2 (
    .d (net51),
    .clk (net49),
    .q (net45)
  );
  dff_cell flop3 (
    .d (net52),
    .clk (net49),
    .q (net42)
  );
  dff_cell flop9 (
    .d (net5),
    .clk (net1),
    .q (net53)
  );
  dff_cell flop10 (
    .d (net4),
    .clk (net1),
    .q (net54)
  );
  dff_cell flop11 (
    .d (net3),
    .clk (net1),
    .q (net55)
  );
  dff_cell flop12 (
    .d (net2),
    .clk (net1),
    .q (net43)
  );
  and_cell and12 (
    .a (net42),
    .b (net55),
    .out (net17)
  );
  and_cell and13 (
    .a (net45),
    .b (net55),
    .out (net21)
  );
  and_cell and14 (
    .a (net46),
    .b (net55),
    .out (net28)
  );
  and_cell and15 (
    .a (net47),
    .b (net55),
    .out (net35)
  );
  xor_cell xor8 (
    .a (net56),
    .b (net24),
    .out (net57)
  );
  and_cell and16 (
    .a (net56),
    .b (net24),
    .out (net58)
  );
  xor_cell xor9 (
    .a (net59),
    .b (net31),
    .out (net60)
  );
  xor_cell xor10 (
    .a (net58),
    .b (net60),
    .out (net61)
  );
  and_cell and17 (
    .a (net59),
    .b (net31),
    .out (net62)
  );
  and_cell and18 (
    .a (net58),
    .b (net60),
    .out (net63)
  );
  or_cell or4 (
    .a (net63),
    .b (net62),
    .out (net64)
  );
  xor_cell xor11 (
    .a (net65),
    .b (net38),
    .out (net66)
  );
  xor_cell xor12 (
    .a (net64),
    .b (net66),
    .out (net67)
  );
  and_cell and19 (
    .a (net65),
    .b (net38),
    .out (net68)
  );
  and_cell and20 (
    .a (net64),
    .b (net66),
    .out (net69)
  );
  or_cell or5 (
    .a (net69),
    .b (net68),
    .out (net70)
  );
  xor_cell xor13 (
    .a (net71),
    .b (net41),
    .out (net72)
  );
  xor_cell xor14 (
    .a (net70),
    .b (net72),
    .out (net73)
  );
  and_cell and21 (
    .a (net71),
    .b (net41),
    .out (net74)
  );
  and_cell and22 (
    .a (net70),
    .b (net72),
    .out (net75)
  );
  or_cell or6 (
    .a (net75),
    .b (net74),
    .out (net76)
  );
  xor_cell xor15 (
    .a (net77),
    .b (net61),
    .out (net78)
  );
  and_cell and23 (
    .a (net77),
    .b (net61),
    .out (net79)
  );
  xor_cell xor16 (
    .a (net80),
    .b (net67),
    .out (net81)
  );
  xor_cell xor17 (
    .a (net79),
    .b (net81),
    .out (net82)
  );
  and_cell and24 (
    .a (net80),
    .b (net67),
    .out (net83)
  );
  and_cell and25 (
    .a (net79),
    .b (net81),
    .out (net84)
  );
  or_cell or7 (
    .a (net84),
    .b (net83),
    .out (net85)
  );
  xor_cell xor18 (
    .a (net86),
    .b (net73),
    .out (net87)
  );
  xor_cell xor19 (
    .a (net85),
    .b (net87),
    .out (net88)
  );
  and_cell and26 (
    .a (net86),
    .b (net73),
    .out (net89)
  );
  and_cell and27 (
    .a (net85),
    .b (net87),
    .out (net90)
  );
  or_cell or8 (
    .a (net90),
    .b (net89),
    .out (net91)
  );
  xor_cell xor20 (
    .a (net92),
    .b (net76),
    .out (net93)
  );
  xor_cell xor21 (
    .a (net91),
    .b (net93),
    .out (net94)
  );
  and_cell and28 (
    .a (net92),
    .b (net76),
    .out (net95)
  );
  and_cell and29 (
    .a (net91),
    .b (net93),
    .out (net96)
  );
  or_cell or9 (
    .a (net96),
    .b (net95),
    .out (net97)
  );
  and_cell and30 (
    .a (net42),
    .b (net54),
    .out (net56)
  );
  and_cell and31 (
    .a (net45),
    .b (net54),
    .out (net59)
  );
  and_cell and32 (
    .a (net46),
    .b (net54),
    .out (net65)
  );
  and_cell and33 (
    .a (net47),
    .b (net54),
    .out (net71)
  );
  and_cell and34 (
    .a (net42),
    .b (net53),
    .out (net77)
  );
  and_cell and35 (
    .a (net45),
    .b (net53),
    .out (net80)
  );
  and_cell and36 (
    .a (net46),
    .b (net53),
    .out (net86)
  );
  and_cell and37 (
    .a (net47),
    .b (net53),
    .out (net92)
  );
  xor_cell xor22 (
    .a (net98),
    .b (net99),
    .out (net100)
  );
  and_cell and38 (
    .a (net98),
    .b (net99),
    .out (net101)
  );
  xor_cell xor23 (
    .a (net102),
    .b (net103),
    .out (net104)
  );
  xor_cell xor24 (
    .a (net101),
    .b (net104),
    .out (net105)
  );
  and_cell and39 (
    .a (net102),
    .b (net103),
    .out (net106)
  );
  and_cell and40 (
    .a (net101),
    .b (net104),
    .out (net107)
  );
  or_cell or10 (
    .a (net107),
    .b (net106),
    .out (net108)
  );
  xor_cell xor25 (
    .a (net109),
    .b (net110),
    .out (net111)
  );
  xor_cell xor26 (
    .a (net108),
    .b (net111),
    .out (net112)
  );
  and_cell and41 (
    .a (net109),
    .b (net110),
    .out (net113)
  );
  and_cell and42 (
    .a (net108),
    .b (net111),
    .out (net114)
  );
  or_cell or11 (
    .a (net114),
    .b (net113),
    .out (net115)
  );
  xor_cell xor27 (
    .a (net116),
    .b (net117),
    .out (net118)
  );
  xor_cell xor28 (
    .a (net115),
    .b (net118),
    .out (net119)
  );
  and_cell and43 (
    .a (net116),
    .b (net117),
    .out (net120)
  );
  and_cell and44 (
    .a (net115),
    .b (net118),
    .out (net121)
  );
  or_cell or12 (
    .a (net121),
    .b (net120),
    .out (net122)
  );
  and_cell and45 (
    .a (net123),
    .b (net124),
    .out (net125)
  );
  and_cell and46 (
    .a (net126),
    .b (net124),
    .out (net99)
  );
  and_cell and47 (
    .a (net127),
    .b (net124),
    .out (net103)
  );
  and_cell and48 (
    .a (net128),
    .b (net124),
    .out (net110)
  );
  dff_cell flop5 (
    .d (net129),
    .clk (net49),
    .q (net128)
  );
  dff_cell flop6 (
    .d (net130),
    .clk (net49),
    .q (net127)
  );
  dff_cell flop7 (
    .d (net131),
    .clk (net49),
    .q (net126)
  );
  dff_cell flop8 (
    .d (net132),
    .clk (net49),
    .q (net123)
  );
  dff_cell flop13 (
    .d (net53),
    .clk (net1),
    .q (net133)
  );
  dff_cell flop14 (
    .d (net54),
    .clk (net1),
    .q (net134)
  );
  dff_cell flop15 (
    .d (net55),
    .clk (net1),
    .q (net135)
  );
  dff_cell flop16 (
    .d (net43),
    .clk (net1),
    .q (net124)
  );
  and_cell and49 (
    .a (net123),
    .b (net135),
    .out (net98)
  );
  and_cell and50 (
    .a (net126),
    .b (net135),
    .out (net102)
  );
  and_cell and51 (
    .a (net127),
    .b (net135),
    .out (net109)
  );
  and_cell and52 (
    .a (net128),
    .b (net135),
    .out (net116)
  );
  xor_cell xor29 (
    .a (net136),
    .b (net105),
    .out (net137)
  );
  and_cell and53 (
    .a (net136),
    .b (net105),
    .out (net138)
  );
  xor_cell xor30 (
    .a (net139),
    .b (net112),
    .out (net140)
  );
  xor_cell xor31 (
    .a (net138),
    .b (net140),
    .out (net141)
  );
  and_cell and54 (
    .a (net139),
    .b (net112),
    .out (net142)
  );
  and_cell and55 (
    .a (net138),
    .b (net140),
    .out (net143)
  );
  or_cell or13 (
    .a (net143),
    .b (net142),
    .out (net144)
  );
  xor_cell xor32 (
    .a (net145),
    .b (net119),
    .out (net146)
  );
  xor_cell xor33 (
    .a (net144),
    .b (net146),
    .out (net147)
  );
  and_cell and56 (
    .a (net145),
    .b (net119),
    .out (net148)
  );
  and_cell and57 (
    .a (net144),
    .b (net146),
    .out (net149)
  );
  or_cell or14 (
    .a (net149),
    .b (net148),
    .out (net150)
  );
  xor_cell xor34 (
    .a (net151),
    .b (net122),
    .out (net152)
  );
  xor_cell xor35 (
    .a (net150),
    .b (net152),
    .out (net153)
  );
  and_cell and58 (
    .a (net151),
    .b (net122),
    .out (net154)
  );
  and_cell and59 (
    .a (net150),
    .b (net152),
    .out (net155)
  );
  or_cell or15 (
    .a (net155),
    .b (net154),
    .out (net156)
  );
  xor_cell xor36 (
    .a (net157),
    .b (net141),
    .out (net158)
  );
  and_cell and60 (
    .a (net157),
    .b (net141),
    .out (net159)
  );
  xor_cell xor37 (
    .a (net160),
    .b (net147),
    .out (net161)
  );
  xor_cell xor38 (
    .a (net159),
    .b (net161),
    .out (net162)
  );
  and_cell and61 (
    .a (net160),
    .b (net147),
    .out (net163)
  );
  and_cell and62 (
    .a (net159),
    .b (net161),
    .out (net164)
  );
  or_cell or16 (
    .a (net164),
    .b (net163),
    .out (net165)
  );
  xor_cell xor39 (
    .a (net166),
    .b (net153),
    .out (net167)
  );
  xor_cell xor40 (
    .a (net165),
    .b (net167),
    .out (net168)
  );
  and_cell and63 (
    .a (net166),
    .b (net153),
    .out (net169)
  );
  and_cell and64 (
    .a (net165),
    .b (net167),
    .out (net170)
  );
  or_cell or17 (
    .a (net170),
    .b (net169),
    .out (net171)
  );
  xor_cell xor41 (
    .a (net172),
    .b (net156),
    .out (net173)
  );
  xor_cell xor42 (
    .a (net171),
    .b (net173),
    .out (net174)
  );
  and_cell and65 (
    .a (net172),
    .b (net156),
    .out (net175)
  );
  and_cell and66 (
    .a (net171),
    .b (net173),
    .out (net176)
  );
  or_cell or18 (
    .a (net176),
    .b (net175),
    .out (net177)
  );
  and_cell and67 (
    .a (net123),
    .b (net134),
    .out (net136)
  );
  and_cell and68 (
    .a (net126),
    .b (net134),
    .out (net139)
  );
  and_cell and69 (
    .a (net127),
    .b (net134),
    .out (net145)
  );
  and_cell and70 (
    .a (net128),
    .b (net134),
    .out (net151)
  );
  and_cell and71 (
    .a (net123),
    .b (net133),
    .out (net157)
  );
  and_cell and72 (
    .a (net126),
    .b (net133),
    .out (net160)
  );
  and_cell and73 (
    .a (net127),
    .b (net133),
    .out (net166)
  );
  and_cell and74 (
    .a (net128),
    .b (net133),
    .out (net172)
  );
  dff_cell flop17 (
    .d (net44),
    .clk (net1),
    .q (net178)
  );
  dff_cell flop18 (
    .d (net19),
    .clk (net1),
    .q (net179)
  );
  dff_cell flop19 (
    .d (net57),
    .clk (net1),
    .q (net180)
  );
  dff_cell flop20 (
    .d (net78),
    .clk (net1),
    .q (net181)
  );
  dff_cell flop21 (
    .d (net82),
    .clk (net1),
    .q (net182)
  );
  dff_cell flop22 (
    .d (net88),
    .clk (net1),
    .q (net183)
  );
  dff_cell flop23 (
    .d (net94),
    .clk (net1),
    .q (net184)
  );
  dff_cell flop24 (
    .d (net97),
    .clk (net1),
    .q (net185)
  );
  dff_cell flop25 (
    .d (net125),
    .clk (net1),
    .q (net186)
  );
  dff_cell flop26 (
    .d (net100),
    .clk (net1),
    .q (net187)
  );
  dff_cell flop27 (
    .d (net137),
    .clk (net1),
    .q (net188)
  );
  dff_cell flop28 (
    .d (net158),
    .clk (net1),
    .q (net189)
  );
  dff_cell flop29 (
    .d (net162),
    .clk (net1),
    .q (net190)
  );
  dff_cell flop30 (
    .d (net168),
    .clk (net1),
    .q (net191)
  );
  dff_cell flop31 (
    .d (net174),
    .clk (net1),
    .q (net192)
  );
  dff_cell flop32 (
    .d (net177),
    .clk (net1),
    .q (net193)
  );
  xor_cell xor43 (
    .a (net186),
    .b (net178),
    .out (net194)
  );
  and_cell and75 (
    .a (net186),
    .b (net178),
    .out (net195)
  );
  xor_cell xor44 (
    .a (net187),
    .b (net179),
    .out (net196)
  );
  xor_cell xor45 (
    .a (net195),
    .b (net196),
    .out (net197)
  );
  and_cell and76 (
    .a (net187),
    .b (net179),
    .out (net198)
  );
  and_cell and77 (
    .a (net195),
    .b (net196),
    .out (net199)
  );
  or_cell or19 (
    .a (net199),
    .b (net198),
    .out (net200)
  );
  xor_cell xor46 (
    .a (net188),
    .b (net180),
    .out (net201)
  );
  xor_cell xor47 (
    .a (net200),
    .b (net201),
    .out (net202)
  );
  and_cell and78 (
    .a (net188),
    .b (net180),
    .out (net203)
  );
  and_cell and79 (
    .a (net200),
    .b (net201),
    .out (net204)
  );
  or_cell or20 (
    .a (net204),
    .b (net203),
    .out (net205)
  );
  xor_cell xor48 (
    .a (net189),
    .b (net181),
    .out (net206)
  );
  xor_cell xor49 (
    .a (net205),
    .b (net206),
    .out (net207)
  );
  and_cell and80 (
    .a (net189),
    .b (net181),
    .out (net208)
  );
  and_cell and81 (
    .a (net205),
    .b (net206),
    .out (net209)
  );
  or_cell or21 (
    .a (net209),
    .b (net208),
    .out (net210)
  );
  xor_cell xor50 (
    .a (net190),
    .b (net182),
    .out (net211)
  );
  xor_cell xor51 (
    .a (net210),
    .b (net211),
    .out (net212)
  );
  and_cell and82 (
    .a (net190),
    .b (net182),
    .out (net213)
  );
  and_cell and83 (
    .a (net210),
    .b (net211),
    .out (net214)
  );
  or_cell or22 (
    .a (net214),
    .b (net213),
    .out (net215)
  );
  xor_cell xor52 (
    .a (net191),
    .b (net183),
    .out (net216)
  );
  xor_cell xor53 (
    .a (net215),
    .b (net216),
    .out (net217)
  );
  and_cell and84 (
    .a (net191),
    .b (net183),
    .out (net218)
  );
  and_cell and85 (
    .a (net215),
    .b (net216),
    .out (net219)
  );
  or_cell or23 (
    .a (net219),
    .b (net218),
    .out (net220)
  );
  xor_cell xor54 (
    .a (net192),
    .b (net184),
    .out (net221)
  );
  xor_cell xor55 (
    .a (net220),
    .b (net221),
    .out (net222)
  );
  and_cell and86 (
    .a (net192),
    .b (net184),
    .out (net223)
  );
  and_cell and87 (
    .a (net220),
    .b (net221),
    .out (net224)
  );
  or_cell or24 (
    .a (net224),
    .b (net223),
    .out (net225)
  );
  xor_cell xor56 (
    .a (net193),
    .b (net185),
    .out (net226)
  );
  xor_cell xor57 (
    .a (net225),
    .b (net226),
    .out (net227)
  );
  and_cell and88 (
    .a (net193),
    .b (net185),
    .out (net228)
  );
  and_cell and89 (
    .a (net225),
    .b (net226),
    .out (net229)
  );
  or_cell or25 (
    .a (net229),
    .b (net228),
    .out (net230)
  );
  mux_cell mux21 (
    .a (net231),
    .b (net232),
    .sel (net7),
    .out (net9)
  );
  mux_cell mux22 (
    .a (net233),
    .b (net234),
    .sel (net7),
    .out (net10)
  );
  mux_cell mux23 (
    .a (net235),
    .b (net236),
    .sel (net7),
    .out (net11)
  );
  mux_cell mux24 (
    .a (net237),
    .b (net238),
    .sel (net7),
    .out (net12)
  );
  mux_cell mux25 (
    .a (net239),
    .b (net240),
    .sel (net7),
    .out (net13)
  );
  mux_cell mux26 (
    .a (net241),
    .b (net242),
    .sel (net7),
    .out (net14)
  );
  mux_cell mux27 (
    .a (net243),
    .b (net244),
    .sel (net7),
    .out (net15)
  );
  mux_cell mux28 (
    .a (net245),
    .b (net246),
    .sel (net7),
    .out (net16)
  );
  mux_cell mux5 (
    .a (net42),
    .b (net178),
    .sel (net6),
    .out (net232)
  );
  mux_cell mux6 (
    .a (net45),
    .b (net179),
    .sel (net6),
    .out (net234)
  );
  mux_cell mux7 (
    .a (net46),
    .b (net180),
    .sel (net6),
    .out (net236)
  );
  mux_cell mux8 (
    .a (net47),
    .b (net181),
    .sel (net6),
    .out (net238)
  );
  mux_cell mux9 (
    .a (net123),
    .b (net182),
    .sel (net6),
    .out (net240)
  );
  mux_cell mux10 (
    .a (net126),
    .b (net183),
    .sel (net6),
    .out (net242)
  );
  mux_cell mux11 (
    .a (net127),
    .b (net184),
    .sel (net6),
    .out (net244)
  );
  mux_cell mux12 (
    .a (net128),
    .b (net185),
    .sel (net6),
    .out (net246)
  );
  mux_cell mux13 (
    .a (net197),
    .b (net186),
    .sel (net6),
    .out (net231)
  );
  mux_cell mux14 (
    .a (net202),
    .b (net187),
    .sel (net6),
    .out (net233)
  );
  mux_cell mux15 (
    .a (net207),
    .b (net188),
    .sel (net6),
    .out (net235)
  );
  mux_cell mux16 (
    .a (net212),
    .b (net189),
    .sel (net6),
    .out (net237)
  );
  mux_cell mux17 (
    .a (net217),
    .b (net190),
    .sel (net6),
    .out (net239)
  );
  mux_cell mux18 (
    .a (net222),
    .b (net191),
    .sel (net6),
    .out (net241)
  );
  mux_cell mux19 (
    .a (net227),
    .b (net192),
    .sel (net6),
    .out (net243)
  );
  mux_cell mux20 (
    .a (net230),
    .b (net193),
    .sel (net6),
    .out (net245)
  );
  dff_cell flop33 (
    .d (net8),
    .clk (net1),
    .notq (net252)
  );
  and_cell and90 (
    .a (net8),
    .b (net252),
    .out (net49)
  );
  dff_cell flop34 (
    .d (net5),
    .clk (net253),
    .q (net48)
  );
  dff_cell flop35 (
    .d (net4),
    .clk (net253),
    .q (net50)
  );
  dff_cell flop36 (
    .d (net3),
    .clk (net253),
    .q (net51)
  );
  dff_cell flop37 (
    .d (net2),
    .clk (net253),
    .q (net52)
  );
  not_cell not1 (
    .in (net49),
    .out (net253)
  );
  dff_cell flop38 (
    .d (net47),
    .clk (net256),
    .q (net129)
  );
  dff_cell flop39 (
    .d (net46),
    .clk (net256),
    .q (net130)
  );
  dff_cell flop40 (
    .d (net45),
    .clk (net256),
    .q (net131)
  );
  dff_cell flop41 (
    .d (net42),
    .clk (net256),
    .q (net132)
  );
  not_cell not2 (
    .in (net253),
    .out (net256)
  );
endmodule
