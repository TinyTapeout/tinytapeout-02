/* Automatically generated from https://wokwi.com/projects/349901899339661908 */

`default_nettype none

module user_module_349901899339661908(
  input [7:0] io_in,
  output [7:0] io_out
);
  wire net1 = io_in[0];
  wire net2 = io_in[2];
  wire net3 = io_in[3];
  wire net4 = io_in[4];
  wire net5 = io_in[5];
  wire net6 = io_in[6];
  wire net7 = io_in[7];
  wire net8;
  wire net9;
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16 = 1'b1;
  wire net17 = 1'b1;
  wire net18 = 1'b1;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98 = 1'b1;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276 = 1'b0;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284;
  wire net285;
  wire net286;
  wire net287;
  wire net288;
  wire net289;
  wire net290;
  wire net291;
  wire net292;
  wire net293;

  assign io_out[0] = net8;
  assign io_out[1] = net9;
  assign io_out[2] = net10;
  assign io_out[3] = net11;
  assign io_out[4] = net12;
  assign io_out[5] = net13;
  assign io_out[6] = net14;
  assign io_out[7] = net15;

  and_cell gate1 (

  );
  or_cell gate2 (

  );
  xor_cell gate3 (

  );
  nand_cell gate4 (

  );
  not_cell gate5 (

  );
  buffer_cell gate6 (

  );
  mux_cell mux1 (

  );
  dff_cell flipflop1 (

  );
  dff_cell flipflop2 (
    .d (net19),
    .clk (net1),
    .q (net20),
    .notq (net21)
  );
  and_cell gate7 (
    .a (net21),
    .b (net18),
    .out (net22)
  );
  and_cell gate8 (
    .a (net23),
    .b (net20),
    .out (net24)
  );
  or_cell gate9 (
    .a (net22),
    .b (net24),
    .out (net25)
  );
  not_cell gate10 (
    .in (net18),
    .out (net23)
  );
  dff_cell flipflop3 (
    .d (net26),
    .clk (net1),
    .q (net27),
    .notq (net28)
  );
  and_cell gate11 (
    .a (net28),
    .b (net29),
    .out (net30)
  );
  and_cell gate12 (
    .a (net31),
    .b (net27),
    .out (net32)
  );
  or_cell gate13 (
    .a (net30),
    .b (net32),
    .out (net33)
  );
  not_cell gate14 (
    .in (net29),
    .out (net31)
  );
  and_cell gate15 (
    .a (net34),
    .b (net20),
    .out (net35)
  );
  and_cell gate16 (
    .a (net7),
    .b (net21),
    .out (net36)
  );
  or_cell gate17 (
    .a (net35),
    .b (net36),
    .out (net29)
  );
  not_cell gate18 (
    .in (net7),
    .out (net34)
  );
  dff_cell flipflop4 (
    .d (net37),
    .clk (net1),
    .q (net38),
    .notq (net39)
  );
  and_cell gate19 (
    .a (net39),
    .b (net40),
    .out (net41)
  );
  and_cell gate20 (
    .a (net42),
    .b (net38),
    .out (net43)
  );
  or_cell gate21 (
    .a (net41),
    .b (net43),
    .out (net44)
  );
  not_cell gate22 (
    .in (net40),
    .out (net42)
  );
  and_cell gate23 (
    .a (net35),
    .b (net27),
    .out (net45)
  );
  and_cell gate24 (
    .a (net28),
    .b (net36),
    .out (net46)
  );
  or_cell gate25 (
    .a (net45),
    .b (net46),
    .out (net40)
  );
  dff_cell flipflop5 (
    .d (net47),
    .clk (net1),
    .q (net48),
    .notq (net49)
  );
  and_cell gate26 (
    .a (net49),
    .b (net50),
    .out (net51)
  );
  and_cell gate27 (
    .a (net52),
    .b (net48),
    .out (net53)
  );
  or_cell gate28 (
    .a (net51),
    .b (net53),
    .out (net54)
  );
  not_cell gate29 (
    .in (net50),
    .out (net52)
  );
  and_cell gate30 (
    .a (net45),
    .b (net38),
    .out (net55)
  );
  and_cell gate31 (
    .a (net39),
    .b (net46),
    .out (net56)
  );
  or_cell gate32 (
    .a (net55),
    .b (net56),
    .out (net50)
  );
  dff_cell flipflop6 (
    .d (net57),
    .clk (net1),
    .q (net58),
    .notq (net59)
  );
  and_cell gate33 (
    .a (net59),
    .b (net60),
    .out (net61)
  );
  and_cell gate34 (
    .a (net62),
    .b (net58),
    .out (net63)
  );
  or_cell gate35 (
    .a (net61),
    .b (net63),
    .out (net64)
  );
  not_cell gate36 (
    .in (net60),
    .out (net62)
  );
  and_cell gate37 (
    .a (net55),
    .b (net48),
    .out (net65)
  );
  and_cell gate38 (
    .a (net49),
    .b (net56),
    .out (net66)
  );
  or_cell gate39 (
    .a (net65),
    .b (net66),
    .out (net60)
  );
  dff_cell flipflop7 (
    .d (net67),
    .clk (net1),
    .q (net68),
    .notq (net69)
  );
  and_cell gate40 (
    .a (net69),
    .b (net70),
    .out (net71)
  );
  and_cell gate41 (
    .a (net72),
    .b (net68),
    .out (net73)
  );
  or_cell gate42 (
    .a (net71),
    .b (net73),
    .out (net74)
  );
  not_cell gate43 (
    .in (net70),
    .out (net72)
  );
  and_cell gate44 (
    .a (net65),
    .b (net58),
    .out (net75)
  );
  and_cell gate45 (
    .a (net59),
    .b (net66),
    .out (net76)
  );
  or_cell gate46 (
    .a (net75),
    .b (net76),
    .out (net70)
  );
  dff_cell flipflop8 (
    .d (net77),
    .clk (net1),
    .q (net78),
    .notq (net79)
  );
  and_cell gate47 (
    .a (net79),
    .b (net80),
    .out (net81)
  );
  and_cell gate48 (
    .a (net82),
    .b (net78),
    .out (net83)
  );
  or_cell gate49 (
    .a (net81),
    .b (net83),
    .out (net84)
  );
  not_cell gate50 (
    .in (net80),
    .out (net82)
  );
  and_cell gate51 (
    .a (net75),
    .b (net68),
    .out (net85)
  );
  and_cell gate52 (
    .a (net69),
    .b (net76),
    .out (net86)
  );
  or_cell gate53 (
    .a (net85),
    .b (net86),
    .out (net80)
  );
  dff_cell flipflop9 (
    .d (net87),
    .clk (net1),
    .q (net88),
    .notq (net89)
  );
  and_cell gate54 (
    .a (net89),
    .b (net90),
    .out (net91)
  );
  and_cell gate55 (
    .a (net92),
    .b (net88),
    .out (net93)
  );
  or_cell gate56 (
    .a (net91),
    .b (net93),
    .out (net94)
  );
  not_cell gate57 (
    .in (net90),
    .out (net92)
  );
  and_cell gate58 (
    .a (net85),
    .b (net78),
    .out (net95)
  );
  and_cell gate59 (
    .a (net79),
    .b (net86),
    .out (net96)
  );
  or_cell gate60 (
    .a (net95),
    .b (net96),
    .out (net90)
  );
  not_cell gate114 (
    .in (net7),
    .out (net97)
  );
  dff_cell flipflop10 (
    .d (net99),
    .clk (net1),
    .q (net100),
    .notq (net101)
  );
  and_cell gate61 (
    .a (net101),
    .b (net98),
    .out (net102)
  );
  and_cell gate62 (
    .a (net103),
    .b (net100),
    .out (net104)
  );
  or_cell gate63 (
    .a (net102),
    .b (net104),
    .out (net105)
  );
  not_cell gate64 (
    .in (net98),
    .out (net103)
  );
  dff_cell flipflop11 (
    .d (net106),
    .clk (net1),
    .q (net107),
    .notq (net108)
  );
  and_cell gate65 (
    .a (net108),
    .b (net109),
    .out (net110)
  );
  and_cell gate66 (
    .a (net111),
    .b (net107),
    .out (net112)
  );
  or_cell gate67 (
    .a (net110),
    .b (net112),
    .out (net113)
  );
  not_cell gate68 (
    .in (net109),
    .out (net111)
  );
  and_cell gate69 (
    .a (net97),
    .b (net100),
    .out (net114)
  );
  and_cell gate70 (
    .a (net7),
    .b (net101),
    .out (net115)
  );
  or_cell gate71 (
    .a (net114),
    .b (net115),
    .out (net109)
  );
  dff_cell flipflop12 (
    .d (net116),
    .clk (net1),
    .q (net117),
    .notq (net118)
  );
  and_cell gate72 (
    .a (net118),
    .b (net119),
    .out (net120)
  );
  and_cell gate73 (
    .a (net121),
    .b (net117),
    .out (net122)
  );
  or_cell gate74 (
    .a (net120),
    .b (net122),
    .out (net123)
  );
  not_cell gate75 (
    .in (net119),
    .out (net121)
  );
  and_cell gate76 (
    .a (net114),
    .b (net107),
    .out (net124)
  );
  and_cell gate77 (
    .a (net108),
    .b (net115),
    .out (net125)
  );
  or_cell gate78 (
    .a (net124),
    .b (net125),
    .out (net119)
  );
  dff_cell flipflop13 (
    .d (net126),
    .clk (net1),
    .q (net127),
    .notq (net128)
  );
  and_cell gate79 (
    .a (net128),
    .b (net129),
    .out (net130)
  );
  and_cell gate80 (
    .a (net131),
    .b (net127),
    .out (net132)
  );
  or_cell gate81 (
    .a (net130),
    .b (net132),
    .out (net133)
  );
  not_cell gate82 (
    .in (net129),
    .out (net131)
  );
  and_cell gate83 (
    .a (net124),
    .b (net117),
    .out (net134)
  );
  and_cell gate84 (
    .a (net118),
    .b (net125),
    .out (net135)
  );
  or_cell gate85 (
    .a (net134),
    .b (net135),
    .out (net129)
  );
  dff_cell flipflop14 (
    .d (net136),
    .clk (net1),
    .q (net137),
    .notq (net138)
  );
  and_cell gate86 (
    .a (net138),
    .b (net139),
    .out (net140)
  );
  and_cell gate87 (
    .a (net141),
    .b (net137),
    .out (net142)
  );
  or_cell gate88 (
    .a (net140),
    .b (net142),
    .out (net143)
  );
  not_cell gate89 (
    .in (net139),
    .out (net141)
  );
  and_cell gate90 (
    .a (net134),
    .b (net127),
    .out (net144)
  );
  and_cell gate91 (
    .a (net128),
    .b (net135),
    .out (net145)
  );
  or_cell gate92 (
    .a (net144),
    .b (net145),
    .out (net139)
  );
  dff_cell flipflop15 (
    .d (net146),
    .clk (net1),
    .q (net147),
    .notq (net148)
  );
  and_cell gate93 (
    .a (net148),
    .b (net149),
    .out (net150)
  );
  and_cell gate94 (
    .a (net151),
    .b (net147),
    .out (net152)
  );
  or_cell gate95 (
    .a (net150),
    .b (net152),
    .out (net153)
  );
  not_cell gate96 (
    .in (net149),
    .out (net151)
  );
  and_cell gate97 (
    .a (net144),
    .b (net137),
    .out (net154)
  );
  and_cell gate98 (
    .a (net138),
    .b (net145),
    .out (net155)
  );
  or_cell gate99 (
    .a (net154),
    .b (net155),
    .out (net149)
  );
  dff_cell flipflop16 (
    .d (net156),
    .clk (net1),
    .q (net157),
    .notq (net158)
  );
  and_cell gate100 (
    .a (net158),
    .b (net159),
    .out (net160)
  );
  and_cell gate101 (
    .a (net161),
    .b (net157),
    .out (net162)
  );
  or_cell gate102 (
    .a (net160),
    .b (net162),
    .out (net163)
  );
  not_cell gate103 (
    .in (net159),
    .out (net161)
  );
  and_cell gate104 (
    .a (net154),
    .b (net147),
    .out (net164)
  );
  and_cell gate105 (
    .a (net148),
    .b (net155),
    .out (net165)
  );
  or_cell gate106 (
    .a (net164),
    .b (net165),
    .out (net159)
  );
  dff_cell flipflop17 (
    .d (net166),
    .clk (net1),
    .q (net167),
    .notq (net168)
  );
  and_cell gate107 (
    .a (net168),
    .b (net169),
    .out (net170)
  );
  and_cell gate108 (
    .a (net171),
    .b (net167),
    .out (net172)
  );
  or_cell gate109 (
    .a (net170),
    .b (net172),
    .out (net173)
  );
  not_cell gate110 (
    .in (net169),
    .out (net171)
  );
  and_cell gate111 (
    .a (net164),
    .b (net157),
    .out (net174)
  );
  and_cell gate112 (
    .a (net158),
    .b (net165),
    .out (net175)
  );
  or_cell gate113 (
    .a (net174),
    .b (net175),
    .out (net169)
  );
  not_cell gate117 (
    .in (net6),
    .out (net176)
  );
  not_cell gate118 (

  );
  not_cell gate130 (

  );
  not_cell gate131 (

  );
  buffer_cell gate132 (
    .in (net177),
    .out (net178)
  );
  buffer_cell gate133 (
    .in (net179),
    .out (net180)
  );
  buffer_cell gate134 (
    .in (net181),
    .out (net182)
  );
  buffer_cell gate135 (
    .in (net183),
    .out (net184)
  );
  not_cell gate136 (
    .in (net182),
    .out (net185)
  );
  not_cell gate137 (
    .in (net184),
    .out (net186)
  );
  not_cell gate138 (
    .in (net180),
    .out (net187)
  );
  not_cell gate139 (
    .in (net178),
    .out (net188)
  );
  and_cell gate140 (
    .a (net182),
    .b (net189),
    .out (net190)
  );
  and_cell gate141 (
    .a (net188),
    .b (net180),
    .out (net189)
  );
  or_cell gate142 (
    .a (net191),
    .b (net192),
    .out (net8)
  );
  and_cell gate143 (
    .a (net178),
    .b (net185),
    .out (net193)
  );
  and_cell gate144 (
    .a (net186),
    .b (net194),
    .out (net195)
  );
  and_cell gate145 (
    .a (net187),
    .b (net178),
    .out (net194)
  );
  and_cell gate146 (
    .a (net184),
    .b (net188),
    .out (net196)
  );
  and_cell gate147 (
    .a (net180),
    .b (net184),
    .out (net197)
  );
  or_cell gate148 (
    .a (net198),
    .b (net197),
    .out (net199)
  );
  or_cell gate149 (
    .a (net196),
    .b (net190),
    .out (net200)
  );
  or_cell gate150 (
    .a (net195),
    .b (net193),
    .out (net192)
  );
  or_cell gate151 (
    .a (net199),
    .b (net200),
    .out (net191)
  );
  and_cell gate152 (
    .a (net178),
    .b (net201),
    .out (net202)
  );
  and_cell gate153 (
    .a (net186),
    .b (net182),
    .out (net201)
  );
  and_cell gate154 (
    .a (net187),
    .b (net185),
    .out (net198)
  );
  and_cell gate155 (
    .a (net188),
    .b (net203),
    .out (net204)
  );
  and_cell gate156 (
    .a (net186),
    .b (net185),
    .out (net203)
  );
  and_cell gate157 (
    .a (net188),
    .b (net184),
    .out (net205)
  );
  and_cell gate158 (
    .a (net205),
    .b (net182),
    .out (net206)
  );
  and_cell gate159 (
    .a (net188),
    .b (net187),
    .out (net207)
  );
  or_cell gate160 (
    .a (net202),
    .b (net207),
    .out (net208)
  );
  or_cell gate161 (
    .a (net206),
    .b (net204),
    .out (net209)
  );
  or_cell gate162 (
    .a (net208),
    .b (net209),
    .out (net210)
  );
  or_cell gate163 (
    .a (net210),
    .b (net198),
    .out (net9)
  );
  and_cell gate164 (
    .a (net178),
    .b (net187),
    .out (net211)
  );
  and_cell gate165 (
    .a (net188),
    .b (net180),
    .out (net212)
  );
  and_cell gate166 (
    .a (net188),
    .b (net186),
    .out (net213)
  );
  and_cell gate167 (
    .a (net188),
    .b (net182),
    .out (net214)
  );
  and_cell gate168 (
    .a (net182),
    .b (net186),
    .out (net215)
  );
  or_cell gate169 (
    .a (net211),
    .b (net212),
    .out (net216)
  );
  or_cell gate170 (
    .a (net213),
    .b (net214),
    .out (net217)
  );
  or_cell gate171 (
    .a (net216),
    .b (net217),
    .out (net218)
  );
  or_cell gate172 (
    .a (net218),
    .b (net215),
    .out (net10)
  );
  and_cell gate173 (
    .a (net180),
    .b (net186),
    .out (net219)
  );
  and_cell gate174 (
    .a (net188),
    .b (net184),
    .out (net220)
  );
  and_cell gate175 (
    .a (net178),
    .b (net180),
    .out (net221)
  );
  and_cell gate176 (
    .a (net219),
    .b (net182),
    .out (net222)
  );
  and_cell gate177 (
    .a (net220),
    .b (net185),
    .out (net223)
  );
  and_cell gate178 (
    .a (net221),
    .b (net185),
    .out (net224)
  );
  and_cell gate179 (
    .a (net187),
    .b (net186),
    .out (net225)
  );
  and_cell gate180 (
    .a (net187),
    .b (net184),
    .out (net226)
  );
  and_cell gate181 (
    .a (net225),
    .b (net185),
    .out (net227)
  );
  and_cell gate182 (
    .a (net226),
    .b (net182),
    .out (net228)
  );
  or_cell gate183 (
    .a (net224),
    .b (net223),
    .out (net229)
  );
  or_cell gate184 (
    .a (net222),
    .b (net228),
    .out (net230)
  );
  or_cell gate185 (
    .a (net229),
    .b (net230),
    .out (net231)
  );
  or_cell gate186 (
    .a (net231),
    .b (net227),
    .out (net11)
  );
  and_cell gate187 (
    .a (net178),
    .b (net184),
    .out (net232)
  );
  and_cell gate188 (
    .a (net178),
    .b (net180),
    .out (net233)
  );
  and_cell gate189 (
    .a (net184),
    .b (net185),
    .out (net234)
  );
  or_cell gate190 (
    .a (net233),
    .b (net232),
    .out (net235)
  );
  or_cell gate191 (
    .a (net198),
    .b (net234),
    .out (net236)
  );
  or_cell gate192 (
    .a (net235),
    .b (net236),
    .out (net12)
  );
  and_cell gate193 (
    .a (net178),
    .b (net187),
    .out (net237)
  );
  and_cell gate194 (
    .a (net213),
    .b (net180),
    .out (net238)
  );
  and_cell gate195 (
    .a (net180),
    .b (net185),
    .out (net239)
  );
  or_cell gate196 (
    .a (net237),
    .b (net232),
    .out (net240)
  );
  or_cell gate197 (
    .a (net238),
    .b (net239),
    .out (net241)
  );
  or_cell gate198 (
    .a (net240),
    .b (net241),
    .out (net242)
  );
  or_cell gate199 (
    .a (net242),
    .b (net203),
    .out (net13)
  );
  and_cell gate200 (
    .a (net237),
    .b (net243),
    .out (net15)
  );
  and_cell gate201 (
    .a (net178),
    .b (net182),
    .out (net244)
  );
  or_cell gate202 (
    .a (net237),
    .b (net238),
    .out (net245)
  );
  or_cell gate203 (
    .a (net244),
    .b (net246),
    .out (net247)
  );
  and_cell gate204 (
    .a (net187),
    .b (net184),
    .out (net246)
  );
  or_cell gate205 (
    .a (net245),
    .b (net247),
    .out (net248)
  );
  or_cell gate206 (
    .a (net234),
    .b (net248),
    .out (net14)
  );
  and_cell gate207 (
    .a (net184),
    .b (net182),
    .out (net243)
  );
  mux_cell mux5 (
    .a (net20),
    .b (net100),
    .sel (net249),
    .out (net250)
  );
  mux_cell mux6 (
    .a (net48),
    .b (net127),
    .sel (net249),
    .out (net251)
  );
  mux_cell mux7 (
    .a (net38),
    .b (net117),
    .sel (net249),
    .out (net252)
  );
  mux_cell mux8 (
    .a (net27),
    .b (net107),
    .sel (net249),
    .out (net253)
  );
  mux_cell mux9 (
    .a (net58),
    .b (net137),
    .sel (net249),
    .out (net254)
  );
  mux_cell mux10 (
    .a (net88),
    .b (net167),
    .sel (net249),
    .out (net255)
  );
  mux_cell mux11 (
    .a (net78),
    .b (net157),
    .sel (net249),
    .out (net256)
  );
  mux_cell mux12 (
    .a (net68),
    .b (net147),
    .sel (net249),
    .out (net257)
  );
  not_cell not1 (
    .in (net5),
    .out (net249)
  );
  mux_cell mux2 (
    .a (net252),
    .b (net256),
    .sel (net4),
    .out (net179)
  );
  mux_cell mux3 (
    .a (net253),
    .b (net257),
    .sel (net4),
    .out (net183)
  );
  mux_cell mux4 (
    .a (net250),
    .b (net254),
    .sel (net4),
    .out (net181)
  );
  mux_cell mux13 (
    .a (net251),
    .b (net255),
    .sel (net4),
    .out (net177)
  );
  not_cell not2 (
    .in (net3),
    .out (net258)
  );
  and_cell and1 (
    .a (net258),
    .b (net25),
    .out (net259)
  );
  and_cell and2 (
    .a (net258),
    .b (net33),
    .out (net260)
  );
  and_cell and3 (
    .a (net258),
    .b (net44),
    .out (net261)
  );
  and_cell and4 (
    .a (net258),
    .b (net54),
    .out (net262)
  );
  and_cell and5 (
    .a (net258),
    .b (net64),
    .out (net263)
  );
  and_cell and6 (
    .a (net258),
    .b (net74),
    .out (net264)
  );
  and_cell and7 (
    .a (net258),
    .b (net84),
    .out (net265)
  );
  and_cell and8 (
    .a (net258),
    .b (net94),
    .out (net266)
  );
  not_cell not3 (
    .in (net3),
    .out (net267)
  );
  and_cell and9 (
    .a (net267),
    .b (net105),
    .out (net268)
  );
  and_cell and10 (
    .a (net267),
    .b (net113),
    .out (net269)
  );
  and_cell and11 (
    .a (net267),
    .b (net123),
    .out (net270)
  );
  and_cell and12 (
    .a (net267),
    .b (net133),
    .out (net271)
  );
  and_cell and13 (
    .a (net267),
    .b (net143),
    .out (net272)
  );
  and_cell and14 (
    .a (net267),
    .b (net153),
    .out (net273)
  );
  and_cell and15 (
    .a (net267),
    .b (net163),
    .out (net274)
  );
  and_cell and16 (
    .a (net267),
    .b (net173),
    .out (net275)
  );
  mux_cell mux14 (
    .a (net20),
    .b (net259),
    .sel (net277),
    .out (net19)
  );
  and_cell and17 (
    .a (net2),
    .b (net6),
    .out (net277)
  );
  mux_cell mux15 (
    .a (net27),
    .b (net260),
    .sel (net278),
    .out (net26)
  );
  buffer_cell gate115 (
    .in (net277),
    .out (net278)
  );
  mux_cell mux16 (
    .a (net38),
    .b (net261),
    .sel (net279),
    .out (net37)
  );
  buffer_cell gate119 (
    .in (net278),
    .out (net279)
  );
  mux_cell mux17 (
    .a (net48),
    .b (net262),
    .sel (net280),
    .out (net47)
  );
  buffer_cell gate120 (
    .in (net279),
    .out (net280)
  );
  mux_cell mux18 (
    .a (net58),
    .b (net263),
    .sel (net281),
    .out (net57)
  );
  buffer_cell gate121 (
    .in (net280),
    .out (net281)
  );
  mux_cell mux19 (
    .a (net68),
    .b (net264),
    .sel (net282),
    .out (net67)
  );
  buffer_cell gate122 (
    .in (net281),
    .out (net282)
  );
  mux_cell mux20 (
    .a (net78),
    .b (net265),
    .sel (net283),
    .out (net77)
  );
  buffer_cell gate123 (
    .in (net282),
    .out (net283)
  );
  mux_cell mux21 (
    .a (net88),
    .b (net266),
    .sel (net284),
    .out (net87)
  );
  buffer_cell gate124 (
    .in (net283),
    .out (net284)
  );
  mux_cell mux22 (
    .a (net100),
    .b (net268),
    .sel (net285),
    .out (net99)
  );
  buffer_cell gate125 (
    .in (net286),
    .out (net285)
  );
  and_cell and18 (
    .a (net2),
    .b (net176),
    .out (net286)
  );
  mux_cell mux23 (
    .a (net107),
    .b (net269),
    .sel (net287),
    .out (net106)
  );
  buffer_cell gate116 (
    .in (net285),
    .out (net287)
  );
  mux_cell mux24 (
    .a (net117),
    .b (net270),
    .sel (net288),
    .out (net116)
  );
  buffer_cell gate126 (
    .in (net287),
    .out (net288)
  );
  mux_cell mux25 (
    .a (net127),
    .b (net271),
    .sel (net289),
    .out (net126)
  );
  buffer_cell gate127 (
    .in (net288),
    .out (net289)
  );
  mux_cell mux26 (
    .a (net137),
    .b (net272),
    .sel (net290),
    .out (net136)
  );
  buffer_cell gate128 (
    .in (net289),
    .out (net290)
  );
  mux_cell mux27 (
    .a (net147),
    .b (net273),
    .sel (net291),
    .out (net146)
  );
  buffer_cell gate129 (
    .in (net290),
    .out (net291)
  );
  mux_cell mux28 (
    .a (net157),
    .b (net274),
    .sel (net292),
    .out (net156)
  );
  buffer_cell gate208 (
    .in (net291),
    .out (net292)
  );
  mux_cell mux29 (
    .a (net167),
    .b (net275),
    .sel (net293),
    .out (net166)
  );
  buffer_cell gate209 (
    .in (net292),
    .out (net293)
  );
endmodule
