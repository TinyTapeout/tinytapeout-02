VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_tto
  CLASS BLOCK ;
  FOREIGN top_tto ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 120.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 2.000 4.040 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.000 11.520 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.000 19.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.000 26.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.000 33.960 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.000 41.440 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.000 48.920 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.000 56.400 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 2.000 63.880 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 2.000 71.360 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.000 78.840 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.000 86.320 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.000 93.800 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.000 101.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 2.000 108.760 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.000 116.240 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.590 5.200 16.190 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.330 5.200 35.930 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.070 5.200 55.670 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.810 5.200 75.410 114.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.460 5.200 26.060 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.200 5.200 45.800 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.940 5.200 65.540 114.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 84.180 114.325 ;
      LAYER met1 ;
        RECT 0.070 4.460 85.030 114.480 ;
      LAYER met2 ;
        RECT 0.100 3.555 85.010 116.125 ;
      LAYER met3 ;
        RECT 2.400 115.240 85.035 116.105 ;
        RECT 1.445 109.160 85.035 115.240 ;
        RECT 2.400 107.760 85.035 109.160 ;
        RECT 1.445 101.680 85.035 107.760 ;
        RECT 2.400 100.280 85.035 101.680 ;
        RECT 1.445 94.200 85.035 100.280 ;
        RECT 2.400 92.800 85.035 94.200 ;
        RECT 1.445 86.720 85.035 92.800 ;
        RECT 2.400 85.320 85.035 86.720 ;
        RECT 1.445 79.240 85.035 85.320 ;
        RECT 2.400 77.840 85.035 79.240 ;
        RECT 1.445 71.760 85.035 77.840 ;
        RECT 2.400 70.360 85.035 71.760 ;
        RECT 1.445 64.280 85.035 70.360 ;
        RECT 2.400 62.880 85.035 64.280 ;
        RECT 1.445 56.800 85.035 62.880 ;
        RECT 2.400 55.400 85.035 56.800 ;
        RECT 1.445 49.320 85.035 55.400 ;
        RECT 2.400 47.920 85.035 49.320 ;
        RECT 1.445 41.840 85.035 47.920 ;
        RECT 2.400 40.440 85.035 41.840 ;
        RECT 1.445 34.360 85.035 40.440 ;
        RECT 2.400 32.960 85.035 34.360 ;
        RECT 1.445 26.880 85.035 32.960 ;
        RECT 2.400 25.480 85.035 26.880 ;
        RECT 1.445 19.400 85.035 25.480 ;
        RECT 2.400 18.000 85.035 19.400 ;
        RECT 1.445 11.920 85.035 18.000 ;
        RECT 2.400 10.520 85.035 11.920 ;
        RECT 1.445 4.440 85.035 10.520 ;
        RECT 2.400 3.040 85.035 4.440 ;
        RECT 1.445 2.900 85.035 3.040 ;
      LAYER met4 ;
        RECT 3.055 4.800 14.190 112.705 ;
        RECT 16.590 4.800 24.060 112.705 ;
        RECT 26.460 4.800 33.930 112.705 ;
        RECT 36.330 4.800 43.800 112.705 ;
        RECT 46.200 4.800 53.670 112.705 ;
        RECT 56.070 4.800 63.540 112.705 ;
        RECT 65.940 4.800 73.410 112.705 ;
        RECT 75.810 4.800 83.425 112.705 ;
        RECT 3.055 2.895 83.425 4.800 ;
  END
END top_tto
END LIBRARY

