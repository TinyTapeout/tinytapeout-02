module secretFile (
    input [7:0] io_in,
    output reg [7:0] io_out
);

wire clk = io_in[0];

reg [8:0] index;

always@(posedge clk) begin
//	if(index == 9'd487)
//		index <= 9'd0;
//	else
	index <= index + 1'd1;
	case(index)
		9'b000000000: io_out <= 8'b01000111;
		9'b000000001: io_out <= 8'b01001001;
		9'b000000010: io_out <= 8'b01000110;
		9'b000000011: io_out <= 8'b00111000;
		9'b000000100: io_out <= 8'b00111001;
		9'b000000101: io_out <= 8'b01100001;
		9'b000000110: io_out <= 8'b00100000;
		9'b000001000: io_out <= 8'b00100000;
		9'b000001010: io_out <= 8'b11110001;
		9'b000001101: io_out <= 8'b01000001;
		9'b000001110: io_out <= 8'b00111000;
		9'b000001111: io_out <= 8'b00101110;
		9'b000010000: io_out <= 8'b10010111;
		9'b000010001: io_out <= 8'b01101000;
		9'b000010010: io_out <= 8'b01100110;
		9'b000010011: io_out <= 8'b10100001;
		9'b000010100: io_out <= 8'b10100010;
		9'b000010101: io_out <= 8'b10110010;
		9'b000011001: io_out <= 8'b00100001;
		9'b000011010: io_out <= 8'b11111111;
		9'b000011011: io_out <= 8'b00001011;
		9'b000011100: io_out <= 8'b01001110;
		9'b000011101: io_out <= 8'b01000101;
		9'b000011110: io_out <= 8'b01010100;
		9'b000011111: io_out <= 8'b01010011;
		9'b000100000: io_out <= 8'b01000011;
		9'b000100001: io_out <= 8'b01000001;
		9'b000100010: io_out <= 8'b01010000;
		9'b000100011: io_out <= 8'b01000101;
		9'b000100100: io_out <= 8'b00110010;
		9'b000100101: io_out <= 8'b00101110;
		9'b000100110: io_out <= 8'b00110000;
		9'b000100111: io_out <= 8'b00000011;
		9'b000101000: io_out <= 8'b00000001;
		9'b000101100: io_out <= 8'b00100001;
		9'b000101101: io_out <= 8'b11111001;
		9'b000101110: io_out <= 8'b00000100;
		9'b000101111: io_out <= 8'b00000100;
		9'b000110000: io_out <= 8'b00011110;
		9'b000110010: io_out <= 8'b11111111;
		9'b000110100: io_out <= 8'b00101100;
		9'b000111001: io_out <= 8'b00100000;
		9'b000111011: io_out <= 8'b00100000;
		9'b000111110: io_out <= 8'b00000010;
		9'b000111111: io_out <= 8'b01110001;
		9'b001000000: io_out <= 8'b10010100;
		9'b001000001: io_out <= 8'b10001111;
		9'b001000010: io_out <= 8'b10101001;
		9'b001000011: io_out <= 8'b11001011;
		9'b001000100: io_out <= 8'b11101101;
		9'b001000101: io_out <= 8'b00001111;
		9'b001000110: io_out <= 8'b10100011;
		9'b001000111: io_out <= 8'b10011100;
		9'b001001000: io_out <= 8'b00110100;
		9'b001001001: io_out <= 8'b10000001;
		9'b001001010: io_out <= 8'b00001011;
		9'b001001011: io_out <= 8'b01000010;
		9'b001001100: io_out <= 8'b01110101;
		9'b001001101: io_out <= 8'b00011000;
		9'b001001110: io_out <= 8'b11101111;
		9'b001001111: io_out <= 8'b00010101;
		9'b001010000: io_out <= 8'b01100100;
		9'b001010001: io_out <= 8'b01000001;
		9'b001010010: io_out <= 8'b00001000;
		9'b001010011: io_out <= 8'b01111100;
		9'b001010100: io_out <= 8'b11001010;
		9'b001010101: io_out <= 8'b10001000;
		9'b001010110: io_out <= 8'b10001110;
		9'b001010111: io_out <= 8'b11100110;
		9'b001011000: io_out <= 8'b10011001;
		9'b001011001: io_out <= 8'b01101010;
		9'b001011010: io_out <= 8'b00101011;
		9'b001011011: io_out <= 8'b11010010;
		9'b001011100: io_out <= 8'b10111010;
		9'b001011101: io_out <= 8'b10101111;
		9'b001011110: io_out <= 8'b00010001;
		9'b001011111: io_out <= 8'b11001111;
		9'b001100000: io_out <= 8'b01000111;
		9'b001100001: io_out <= 8'b01101011;
		9'b001100010: io_out <= 8'b11011111;
		9'b001100011: io_out <= 8'b01101001;
		9'b001100100: io_out <= 8'b10101110;
		9'b001100101: io_out <= 8'b10101011;
		9'b001100110: io_out <= 8'b01111100;
		9'b001100111: io_out <= 8'b11101100;
		9'b001101000: io_out <= 8'b00110011;
		9'b001101001: io_out <= 8'b10000101;
		9'b001101010: io_out <= 8'b01110000;
		9'b001101011: io_out <= 8'b00011101;
		9'b001101100: io_out <= 8'b10011001;
		9'b001101101: io_out <= 8'b10000100;
		9'b001101110: io_out <= 8'b10010100;
		9'b001101111: io_out <= 8'b00010001;
		9'b001110000: io_out <= 8'b11111000;
		9'b001110001: io_out <= 8'b00111010;
		9'b001110010: io_out <= 8'b00010111;
		9'b001110011: io_out <= 8'b01100011;
		9'b001110100: io_out <= 8'b01100011;
		9'b001110101: io_out <= 8'b01010100;
		9'b001110110: io_out <= 8'b01010100;
		9'b001110111: io_out <= 8'b11010010;
		9'b001111000: io_out <= 8'b10011000;
		9'b001111001: io_out <= 8'b01001001;
		9'b001111010: io_out <= 8'b00001000;
		9'b001111011: io_out <= 8'b10110101;
		9'b001111100: io_out <= 8'b00001001;
		9'b001111101: io_out <= 8'b10111101;
		9'b001111110: io_out <= 8'b01000110;
		9'b001111111: io_out <= 8'b10101110;
		9'b010000000: io_out <= 8'b00100010;
		9'b010000001: io_out <= 8'b01101110;
		9'b010000010: io_out <= 8'b11001001;
		9'b010000011: io_out <= 8'b01111010;
		9'b010000100: io_out <= 8'b11001101;
		9'b010000101: io_out <= 8'b01101010;
		9'b010000110: io_out <= 8'b11000001;
		9'b010000111: io_out <= 8'b01010100;
		9'b010001000: io_out <= 8'b00010010;
		9'b010001001: io_out <= 8'b10001010;
		9'b010001010: io_out <= 8'b10111001;
		9'b010001011: io_out <= 8'b11100101;
		9'b010001100: io_out <= 8'b00001110;
		9'b010001101: io_out <= 8'b11000101;
		9'b010001110: io_out <= 8'b10010111;
		9'b010001111: io_out <= 8'b10110100;
		9'b010010000: io_out <= 8'b11110111;
		9'b010010001: io_out <= 8'b11011100;
		9'b010010010: io_out <= 8'b01110001;
		9'b010010011: io_out <= 8'b10111111;
		9'b010010100: io_out <= 8'b10010001;
		9'b010010101: io_out <= 8'b01001101;
		9'b010010110: io_out <= 8'b10110010;
		9'b010010111: io_out <= 8'b10010111;
		9'b010011000: io_out <= 8'b11111011;
		9'b010011001: io_out <= 8'b01100000;
		9'b010011010: io_out <= 8'b11011111;
		9'b010011011: io_out <= 8'b10011001;
		9'b010011100: io_out <= 8'b11001110;
		9'b010011101: io_out <= 8'b00000100;
		9'b010011110: io_out <= 8'b01111100;
		9'b010011111: io_out <= 8'b10001111;
		9'b010100000: io_out <= 8'b11110110;
		9'b010100001: io_out <= 8'b11110100;
		9'b010100010: io_out <= 8'b00000111;
		9'b010100011: io_out <= 8'b01011000;
		9'b010100100: io_out <= 8'b11100111;
		9'b010100101: io_out <= 8'b10100000;
		9'b010100110: io_out <= 8'b00000111;
		9'b010100111: io_out <= 8'b11011000;
		9'b010101000: io_out <= 8'b01110111;
		9'b010101001: io_out <= 8'b01000010;
		9'b010101010: io_out <= 8'b01011000;
		9'b010101011: io_out <= 8'b01111000;
		9'b010101100: io_out <= 8'b10100100;
		9'b010101101: io_out <= 8'b11000110;
		9'b010101110: io_out <= 8'b11010111;
		9'b010101111: io_out <= 8'b01010000;
		9'b010110010: io_out <= 8'b00100001;
		9'b010110011: io_out <= 8'b11111001;
		9'b010110100: io_out <= 8'b00000100;
		9'b010110101: io_out <= 8'b00000101;
		9'b010110110: io_out <= 8'b00011110;
		9'b010111000: io_out <= 8'b00000011;
		9'b010111010: io_out <= 8'b00101100;
		9'b010111011: io_out <= 8'b00000101;
		9'b010111101: io_out <= 8'b00000011;
		9'b010111111: io_out <= 8'b00011000;
		9'b011000001: io_out <= 8'b00011101;
		9'b011000100: io_out <= 8'b00000010;
		9'b011000101: io_out <= 8'b01100010;
		9'b011000110: io_out <= 8'b10010100;
		9'b011000111: io_out <= 8'b10001111;
		9'b011001000: io_out <= 8'b00010010;
		9'b011001010: io_out <= 8'b11101001;
		9'b011001011: io_out <= 8'b10101111;
		9'b011001100: io_out <= 8'b00011000;
		9'b011001101: io_out <= 8'b00001011;
		9'b011001110: io_out <= 8'b10110000;
		9'b011001111: io_out <= 8'b00001010;
		9'b011010000: io_out <= 8'b10111001;
		9'b011010001: io_out <= 8'b10011010;
		9'b011010010: io_out <= 8'b01111101;
		9'b011010011: io_out <= 8'b00100000;
		9'b011010100: io_out <= 8'b01111000;
		9'b011010101: io_out <= 8'b10111111;
		9'b011010110: io_out <= 8'b00111001;
		9'b011010111: io_out <= 8'b11011111;
		9'b011011000: io_out <= 8'b00011000;
		9'b011011001: io_out <= 8'b10001010;
		9'b011011010: io_out <= 8'b00100011;
		9'b011011011: io_out <= 8'b01010101;
		9'b011011100: io_out <= 8'b00100010;
		9'b011011101: io_out <= 8'b00100111;
		9'b011011110: io_out <= 8'b10011010;
		9'b011011111: io_out <= 8'b00011010;
		9'b011100000: io_out <= 8'b01101011;
		9'b011100001: io_out <= 8'b10101011;
		9'b011100010: io_out <= 8'b01111110;
		9'b011100011: io_out <= 8'b01110000;
		9'b011100100: io_out <= 8'b00101100;
		9'b011100101: io_out <= 8'b11001111;
		9'b011100110: io_out <= 8'b11101110;
		9'b011100111: io_out <= 8'b01101001;
		9'b011101000: io_out <= 8'b11001011;
		9'b011101001: io_out <= 8'b01011001;
		9'b011101010: io_out <= 8'b11000111;
		9'b011101011: io_out <= 8'b01010110;
		9'b011101100: io_out <= 8'b10010100;
		9'b011101101: io_out <= 8'b00101110;
		9'b011101110: io_out <= 8'b11000001;
		9'b011101111: io_out <= 8'b11111000;
		9'b011110000: io_out <= 8'b01111110;
		9'b011110001: io_out <= 8'b10100000;
		9'b011110010: io_out <= 8'b01100000;
		9'b011110011: io_out <= 8'b00010000;
		9'b011110100: io_out <= 8'b10010010;
		9'b011110101: io_out <= 8'b00011001;
		9'b011110110: io_out <= 8'b00011001;
		9'b011110111: io_out <= 8'b10001111;
		9'b011111000: io_out <= 8'b10001001;
		9'b011111001: io_out <= 8'b00011101;
		9'b011111010: io_out <= 8'b11001111;
		9'b011111011: io_out <= 8'b10110011;
		9'b011111100: io_out <= 8'b10010100;
		9'b011111101: io_out <= 8'b10001000;
		9'b011111110: io_out <= 8'b10001100;
		9'b011111111: io_out <= 8'b10011111;
		9'b100000000: io_out <= 8'b00101000;
		9'b100000001: io_out <= 8'b01100011;
		9'b100000010: io_out <= 8'b00011010;
		9'b100000011: io_out <= 8'b01110100;
		9'b100000100: io_out <= 8'b01000110;
		9'b100000101: io_out <= 8'b10110001;
		9'b100000110: io_out <= 8'b01011001;
		9'b100000111: io_out <= 8'b11101011;
		9'b100001000: io_out <= 8'b10100100;
		9'b100001001: io_out <= 8'b10111001;
		9'b100001010: io_out <= 8'b11010100;
		9'b100001011: io_out <= 8'b01010010;
		9'b100001100: io_out <= 8'b11000001;
		9'b100001101: io_out <= 8'b01011101;
		9'b100001110: io_out <= 8'b11101111;
		9'b100001111: io_out <= 8'b00110101;
		9'b100010000: io_out <= 8'b01100001;
		9'b100010001: io_out <= 8'b10110110;
		9'b100010010: io_out <= 8'b00110110;
		9'b100010011: io_out <= 8'b11000101;
		9'b100010100: io_out <= 8'b01101001;
		9'b100010101: io_out <= 8'b01110010;
		9'b100010110: io_out <= 8'b11011010;
		9'b100010111: io_out <= 8'b11101000;
		9'b100011000: io_out <= 8'b01111110;
		9'b100011001: io_out <= 8'b01001011;
		9'b100011010: io_out <= 8'b00001111;
		9'b100011011: io_out <= 8'b01010101;
		9'b100011100: io_out <= 8'b11111001;
		9'b100011101: io_out <= 8'b11111100;
		9'b100011110: io_out <= 8'b11000110;
		9'b100011111: io_out <= 8'b00110110;
		9'b100100000: io_out <= 8'b11010011;
		9'b100100001: io_out <= 8'b10101000;
		9'b100100010: io_out <= 8'b11100110;
		9'b100100011: io_out <= 8'b01011110;
		9'b100100100: io_out <= 8'b00111110;
		9'b100100101: io_out <= 8'b11011111;
		9'b100100110: io_out <= 8'b01010001;
		9'b100101001: io_out <= 8'b00100001;
		9'b100101010: io_out <= 8'b11111001;
		9'b100101011: io_out <= 8'b00000100;
		9'b100101100: io_out <= 8'b00000101;
		9'b100101101: io_out <= 8'b00011110;
		9'b100101111: io_out <= 8'b00000011;
		9'b100110001: io_out <= 8'b00101100;
		9'b100110110: io_out <= 8'b00011101;
		9'b100111000: io_out <= 8'b00100000;
		9'b100111011: io_out <= 8'b00000010;
		9'b100111100: io_out <= 8'b01111101;
		9'b100111101: io_out <= 8'b10010100;
		9'b100111110: io_out <= 8'b10001111;
		9'b100111111: io_out <= 8'b00010110;
		9'b101000000: io_out <= 8'b00011011;
		9'b101000001: io_out <= 8'b11101001;
		9'b101000010: io_out <= 8'b11101111;
		9'b101000011: io_out <= 8'b00000010;
		9'b101000100: io_out <= 8'b10011000;
		9'b101000101: io_out <= 8'b10100000;
		9'b101000110: io_out <= 8'b11000001;
		9'b101000111: io_out <= 8'b10001011;
		9'b101001000: io_out <= 8'b00100100;
		9'b101001001: io_out <= 8'b10011101;
		9'b101001010: io_out <= 8'b10111000;
		9'b101001011: io_out <= 8'b10001011;
		9'b101001100: io_out <= 8'b11001101;
		9'b101001101: io_out <= 8'b01111000;
		9'b101001110: io_out <= 8'b10010111;
		9'b101001111: io_out <= 8'b11000110;
		9'b101010000: io_out <= 8'b00101100;
		9'b101010001: io_out <= 8'b00100010;
		9'b101010010: io_out <= 8'b01000100;
		9'b101010011: io_out <= 8'b10010101;
		9'b101010100: io_out <= 8'b11010110;
		9'b101010101: io_out <= 8'b10011001;
		9'b101010110: io_out <= 8'b10010000;
		9'b101010111: io_out <= 8'b00100101;
		9'b101011000: io_out <= 8'b00011011;
		9'b101011001: io_out <= 8'b10101001;
		9'b101011010: io_out <= 8'b00100110;
		9'b101011011: io_out <= 8'b11011100;
		9'b101011100: io_out <= 8'b11001010;
		9'b101011101: io_out <= 8'b01110100;
		9'b101011110: io_out <= 8'b10101101;
		9'b101011111: io_out <= 8'b11011110;
		9'b101100000: io_out <= 8'b10000111;
		9'b101100001: io_out <= 8'b10111100;
		9'b101100010: io_out <= 8'b11011110;
		9'b101100011: io_out <= 8'b10010010;
		9'b101100100: io_out <= 8'b01001101;
		9'b101100101: io_out <= 8'b11010011;
		9'b101100110: io_out <= 8'b01001100;
		9'b101100111: io_out <= 8'b01111000;
		9'b101101000: io_out <= 8'b01000011;
		9'b101101001: io_out <= 8'b10001111;
		9'b101101010: io_out <= 8'b01110000;
		9'b101101011: io_out <= 8'b00100011;
		9'b101101100: io_out <= 8'b00110000;
		9'b101101101: io_out <= 8'b00101101;
		9'b101101110: io_out <= 8'b01010010;
		9'b101101111: io_out <= 8'b10011101;
		9'b101110000: io_out <= 8'b00001101;
		9'b101110001: io_out <= 8'b00110010;
		9'b101110010: io_out <= 8'b10011001;
		9'b101110011: io_out <= 8'b00010100;
		9'b101110100: io_out <= 8'b11110110;
		9'b101110101: io_out <= 8'b00100010;
		9'b101110110: io_out <= 8'b11001110;
		9'b101110111: io_out <= 8'b11010100;
		9'b101111000: io_out <= 8'b10110010;
		9'b101111001: io_out <= 8'b11110010;
		9'b101111010: io_out <= 8'b01000100;
		9'b101111011: io_out <= 8'b01010101;
		9'b101111100: io_out <= 8'b10101101;
		9'b101111101: io_out <= 8'b11000011;
		9'b101111110: io_out <= 8'b11101100;
		9'b101111111: io_out <= 8'b01100011;
		9'b110000000: io_out <= 8'b11001011;
		9'b110000001: io_out <= 8'b00000101;
		9'b110000010: io_out <= 8'b01111100;
		9'b110000011: io_out <= 8'b00101000;
		9'b110000100: io_out <= 8'b00100011;
		9'b110000101: io_out <= 8'b11110000;
		9'b110000110: io_out <= 8'b11110000;
		9'b110000111: io_out <= 8'b01001000;
		9'b110001000: io_out <= 8'b10000110;
		9'b110001001: io_out <= 8'b10100000;
		9'b110001010: io_out <= 8'b10101011;
		9'b110001011: io_out <= 8'b01101011;
		9'b110001100: io_out <= 8'b10110001;
		9'b110001101: io_out <= 8'b11010110;
		9'b110001110: io_out <= 8'b01101100;
		9'b110001111: io_out <= 8'b10111110;
		9'b110010000: io_out <= 8'b11000000;
		9'b110010001: io_out <= 8'b11100001;
		9'b110010010: io_out <= 8'b11010011;
		9'b110010011: io_out <= 8'b11000011;
		9'b110010100: io_out <= 8'b00011100;
		9'b110010101: io_out <= 8'b10111011;
		9'b110010110: io_out <= 8'b00001101;
		9'b110010111: io_out <= 8'b00100001;
		9'b110011000: io_out <= 8'b11100110;
		9'b110011001: io_out <= 8'b10001100;
		9'b110011010: io_out <= 8'b11111100;
		9'b110011011: io_out <= 8'b01001100;
		9'b110011100: io_out <= 8'b11000001;
		9'b110011101: io_out <= 8'b01110111;
		9'b110011110: io_out <= 8'b11000101;
		9'b110011111: io_out <= 8'b00110110;
		9'b110100000: io_out <= 8'b01110101;
		9'b110100001: io_out <= 8'b11010111;
		9'b110100010: io_out <= 8'b01110110;
		9'b110100011: io_out <= 8'b00000110;
		9'b110100100: io_out <= 8'b00000101;
		9'b110100101: io_out <= 8'b01111000;
		9'b110100110: io_out <= 8'b00000111;
		9'b110100111: io_out <= 8'b10100110;
		9'b110101000: io_out <= 8'b10110111;
		9'b110101001: io_out <= 8'b10100011;
		9'b110101010: io_out <= 8'b01001000;
		9'b110101011: io_out <= 8'b10010110;
		9'b110101100: io_out <= 8'b11110011;
		9'b110101101: io_out <= 8'b11100101;
		9'b110101110: io_out <= 8'b01111000;
		9'b110101111: io_out <= 8'b11100010;
		9'b110110000: io_out <= 8'b01011000;
		9'b110110001: io_out <= 8'b00100001;
		9'b110110010: io_out <= 8'b01000010;
		9'b110110011: io_out <= 8'b01011001;
		9'b110110100: io_out <= 8'b01000111;
		9'b110110101: io_out <= 8'b11100101;
		9'b110110110: io_out <= 8'b10001000;
		9'b110110111: io_out <= 8'b01101001;
		9'b110111000: io_out <= 8'b01010000;
		9'b110111011: io_out <= 8'b00111011;
		9'b110111100: io_out <= 8'b01100010;
		9'b110111101: io_out <= 8'b01101001;
		9'b110111110: io_out <= 8'b01110100;
		9'b110111111: io_out <= 8'b01101100;
		9'b111000000: io_out <= 8'b01110101;
		9'b111000001: io_out <= 8'b01101110;
		9'b111000010: io_out <= 8'b01101001;
		default: io_out <= 8'b00000000;
	endcase;
end

endmodule
