magic
tech sky130B
magscale 1 2
timestamp 1669905304
<< viali >>
rect 17693 17289 17727 17323
rect 20913 17289 20947 17323
rect 31033 17289 31067 17323
rect 40877 17289 40911 17323
rect 44097 17289 44131 17323
rect 2973 17221 3007 17255
rect 3985 17221 4019 17255
rect 38853 17221 38887 17255
rect 2237 17153 2271 17187
rect 4629 17153 4663 17187
rect 6745 17153 6779 17187
rect 8033 17153 8067 17187
rect 9965 17153 9999 17187
rect 11529 17153 11563 17187
rect 13185 17153 13219 17187
rect 14473 17153 14507 17187
rect 16681 17153 16715 17187
rect 17509 17153 17543 17187
rect 19625 17153 19659 17187
rect 20729 17153 20763 17187
rect 22845 17153 22879 17187
rect 24593 17153 24627 17187
rect 26065 17153 26099 17187
rect 27997 17153 28031 17187
rect 29745 17153 29779 17187
rect 31217 17153 31251 17187
rect 32321 17153 32355 17187
rect 34897 17153 34931 17187
rect 35725 17153 35759 17187
rect 37657 17153 37691 17187
rect 40693 17153 40727 17187
rect 42625 17153 42659 17187
rect 43913 17153 43947 17187
rect 2421 17085 2455 17119
rect 4905 17085 4939 17119
rect 11805 17085 11839 17119
rect 32597 17085 32631 17119
rect 43453 17085 43487 17119
rect 4169 17017 4203 17051
rect 3065 16949 3099 16983
rect 9781 16949 9815 16983
rect 16865 16949 16899 16983
rect 24409 16949 24443 16983
rect 34713 16949 34747 16983
rect 38945 16949 38979 16983
rect 3985 16745 4019 16779
rect 43453 16745 43487 16779
rect 44097 16745 44131 16779
rect 2053 16677 2087 16711
rect 1869 16541 1903 16575
rect 16497 16541 16531 16575
rect 17141 16541 17175 16575
rect 40049 16541 40083 16575
rect 16313 16405 16347 16439
rect 16957 16405 16991 16439
rect 39865 16405 39899 16439
rect 44189 15861 44223 15895
rect 1409 15453 1443 15487
rect 18521 15453 18555 15487
rect 19533 15453 19567 15487
rect 34897 15453 34931 15487
rect 19257 15385 19291 15419
rect 19441 15385 19475 15419
rect 1593 15317 1627 15351
rect 18337 15317 18371 15351
rect 19533 15317 19567 15351
rect 34713 15317 34747 15351
rect 20085 15113 20119 15147
rect 18061 15045 18095 15079
rect 18981 15045 19015 15079
rect 8769 14977 8803 15011
rect 12449 14977 12483 15011
rect 12909 14977 12943 15011
rect 13093 14977 13127 15011
rect 13737 14977 13771 15011
rect 16865 14977 16899 15011
rect 17877 14977 17911 15011
rect 18889 14977 18923 15011
rect 19073 14977 19107 15011
rect 19901 14977 19935 15011
rect 20177 14977 20211 15011
rect 8585 14909 8619 14943
rect 22845 14909 22879 14943
rect 23121 14909 23155 14943
rect 18705 14841 18739 14875
rect 8953 14773 8987 14807
rect 12265 14773 12299 14807
rect 13001 14773 13035 14807
rect 13553 14773 13587 14807
rect 16681 14773 16715 14807
rect 18245 14773 18279 14807
rect 19257 14773 19291 14807
rect 19717 14773 19751 14807
rect 9137 14569 9171 14603
rect 20545 14569 20579 14603
rect 23857 14569 23891 14603
rect 9321 14501 9355 14535
rect 21741 14501 21775 14535
rect 19717 14433 19751 14467
rect 19809 14433 19843 14467
rect 7573 14365 7607 14399
rect 8217 14365 8251 14399
rect 11989 14365 12023 14399
rect 12173 14365 12207 14399
rect 13093 14365 13127 14399
rect 13185 14365 13219 14399
rect 13277 14365 13311 14399
rect 13461 14365 13495 14399
rect 15485 14365 15519 14399
rect 17325 14365 17359 14399
rect 19533 14365 19567 14399
rect 19625 14365 19659 14399
rect 21925 14365 21959 14399
rect 22477 14365 22511 14399
rect 42993 14365 43027 14399
rect 43913 14365 43947 14399
rect 8953 14297 8987 14331
rect 9153 14297 9187 14331
rect 15752 14297 15786 14331
rect 17592 14297 17626 14331
rect 20361 14297 20395 14331
rect 20561 14297 20595 14331
rect 22722 14297 22756 14331
rect 7389 14229 7423 14263
rect 8033 14229 8067 14263
rect 12357 14229 12391 14263
rect 12817 14229 12851 14263
rect 16865 14229 16899 14263
rect 18705 14229 18739 14263
rect 19349 14229 19383 14263
rect 20729 14229 20763 14263
rect 42809 14229 42843 14263
rect 44097 14229 44131 14263
rect 3157 14025 3191 14059
rect 12265 14025 12299 14059
rect 14657 14025 14691 14059
rect 16129 14025 16163 14059
rect 17601 14025 17635 14059
rect 20177 14025 20211 14059
rect 21097 14025 21131 14059
rect 23397 14025 23431 14059
rect 33333 14025 33367 14059
rect 7634 13957 7668 13991
rect 9597 13957 9631 13991
rect 10425 13957 10459 13991
rect 11897 13957 11931 13991
rect 12113 13957 12147 13991
rect 18245 13957 18279 13991
rect 18461 13957 18495 13991
rect 19993 13957 20027 13991
rect 22262 13957 22296 13991
rect 24869 13957 24903 13991
rect 33701 13957 33735 13991
rect 3341 13889 3375 13923
rect 3985 13889 4019 13923
rect 4252 13889 4286 13923
rect 10241 13889 10275 13923
rect 12725 13889 12759 13923
rect 12981 13889 13015 13923
rect 14565 13889 14599 13923
rect 15945 13889 15979 13923
rect 16681 13889 16715 13923
rect 17785 13889 17819 13923
rect 19625 13889 19659 13923
rect 21281 13889 21315 13923
rect 24041 13889 24075 13923
rect 25053 13889 25087 13923
rect 1593 13821 1627 13855
rect 7389 13821 7423 13855
rect 15761 13821 15795 13855
rect 16773 13821 16807 13855
rect 22017 13821 22051 13855
rect 23949 13821 23983 13855
rect 25237 13821 25271 13855
rect 33793 13821 33827 13855
rect 33885 13821 33919 13855
rect 9229 13753 9263 13787
rect 10609 13753 10643 13787
rect 14105 13753 14139 13787
rect 5365 13685 5399 13719
rect 8769 13685 8803 13719
rect 9597 13685 9631 13719
rect 9781 13685 9815 13719
rect 12081 13685 12115 13719
rect 18429 13685 18463 13719
rect 18613 13685 18647 13719
rect 19993 13685 20027 13719
rect 24409 13685 24443 13719
rect 8401 13481 8435 13515
rect 9321 13481 9355 13515
rect 9505 13481 9539 13515
rect 8953 13413 8987 13447
rect 14197 13413 14231 13447
rect 14841 13413 14875 13447
rect 17969 13413 18003 13447
rect 18613 13413 18647 13447
rect 19257 13413 19291 13447
rect 40325 13413 40359 13447
rect 41061 13413 41095 13447
rect 17693 13345 17727 13379
rect 21465 13345 21499 13379
rect 23213 13345 23247 13379
rect 37289 13345 37323 13379
rect 37749 13345 37783 13379
rect 7021 13277 7055 13311
rect 10517 13277 10551 13311
rect 11161 13277 11195 13311
rect 11805 13277 11839 13311
rect 12061 13277 12095 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 15022 13277 15056 13311
rect 15393 13277 15427 13311
rect 15485 13277 15519 13311
rect 15945 13277 15979 13311
rect 16313 13277 16347 13311
rect 17601 13277 17635 13311
rect 18521 13277 18555 13311
rect 18705 13277 18739 13311
rect 19441 13277 19475 13311
rect 21005 13277 21039 13311
rect 23673 13277 23707 13311
rect 23857 13277 23891 13311
rect 26341 13277 26375 13311
rect 26801 13277 26835 13311
rect 30297 13277 30331 13311
rect 32781 13277 32815 13311
rect 37381 13277 37415 13311
rect 38301 13277 38335 13311
rect 38393 13277 38427 13311
rect 39129 13277 39163 13311
rect 40601 13277 40635 13311
rect 41337 13277 41371 13311
rect 7288 13209 7322 13243
rect 9321 13209 9355 13243
rect 16129 13209 16163 13243
rect 16221 13209 16255 13243
rect 21741 13209 21775 13243
rect 27077 13209 27111 13243
rect 33048 13209 33082 13243
rect 40325 13209 40359 13243
rect 41061 13209 41095 13243
rect 10609 13141 10643 13175
rect 11253 13141 11287 13175
rect 13185 13141 13219 13175
rect 15025 13141 15059 13175
rect 16497 13141 16531 13175
rect 20821 13141 20855 13175
rect 23765 13141 23799 13175
rect 26157 13141 26191 13175
rect 28549 13141 28583 13175
rect 30389 13141 30423 13175
rect 34161 13141 34195 13175
rect 38577 13141 38611 13175
rect 39221 13141 39255 13175
rect 40509 13141 40543 13175
rect 41245 13141 41279 13175
rect 22293 12937 22327 12971
rect 22385 12937 22419 12971
rect 23305 12937 23339 12971
rect 23857 12937 23891 12971
rect 24041 12937 24075 12971
rect 33517 12937 33551 12971
rect 34437 12937 34471 12971
rect 35633 12937 35667 12971
rect 38669 12937 38703 12971
rect 39421 12937 39455 12971
rect 4712 12869 4746 12903
rect 8677 12869 8711 12903
rect 9045 12869 9079 12903
rect 13645 12869 13679 12903
rect 13829 12869 13863 12903
rect 25237 12869 25271 12903
rect 25437 12869 25471 12903
rect 39221 12869 39255 12903
rect 3157 12801 3191 12835
rect 4445 12801 4479 12835
rect 8861 12801 8895 12835
rect 9873 12801 9907 12835
rect 10701 12801 10735 12835
rect 11989 12801 12023 12835
rect 13001 12801 13035 12835
rect 13461 12801 13495 12835
rect 14473 12801 14507 12835
rect 14657 12801 14691 12835
rect 14749 12801 14783 12835
rect 15209 12801 15243 12835
rect 15393 12801 15427 12835
rect 15485 12801 15519 12835
rect 15761 12801 15795 12835
rect 16681 12801 16715 12835
rect 18475 12801 18509 12835
rect 19901 12801 19935 12835
rect 20913 12801 20947 12835
rect 23121 12801 23155 12835
rect 23397 12801 23431 12835
rect 23982 12801 24016 12835
rect 26249 12801 26283 12835
rect 31585 12801 31619 12835
rect 32137 12801 32171 12835
rect 32393 12801 32427 12835
rect 34345 12801 34379 12835
rect 35541 12801 35575 12835
rect 37556 12801 37590 12835
rect 40509 12801 40543 12835
rect 40776 12801 40810 12835
rect 9781 12733 9815 12767
rect 15577 12733 15611 12767
rect 17049 12733 17083 12767
rect 20269 12733 20303 12767
rect 21005 12733 21039 12767
rect 21097 12733 21131 12767
rect 22477 12733 22511 12767
rect 24501 12733 24535 12767
rect 26065 12733 26099 12767
rect 26985 12733 27019 12767
rect 27261 12733 27295 12767
rect 29193 12733 29227 12767
rect 29469 12733 29503 12767
rect 34529 12733 34563 12767
rect 35725 12733 35759 12767
rect 37289 12733 37323 12767
rect 10241 12665 10275 12699
rect 19717 12665 19751 12699
rect 20545 12665 20579 12699
rect 21925 12665 21959 12699
rect 25605 12665 25639 12699
rect 31401 12665 31435 12699
rect 33977 12665 34011 12699
rect 2973 12597 3007 12631
rect 5825 12597 5859 12631
rect 10885 12597 10919 12631
rect 12081 12597 12115 12631
rect 12817 12597 12851 12631
rect 14473 12597 14507 12631
rect 15945 12597 15979 12631
rect 23121 12597 23155 12631
rect 24409 12597 24443 12631
rect 25421 12597 25455 12631
rect 26433 12597 26467 12631
rect 28733 12597 28767 12631
rect 30941 12597 30975 12631
rect 35173 12597 35207 12631
rect 39405 12597 39439 12631
rect 39589 12597 39623 12631
rect 41889 12597 41923 12631
rect 44189 12597 44223 12631
rect 6101 12393 6135 12427
rect 14197 12393 14231 12427
rect 14933 12393 14967 12427
rect 22339 12393 22373 12427
rect 23673 12393 23707 12427
rect 24593 12393 24627 12427
rect 25237 12393 25271 12427
rect 25697 12393 25731 12427
rect 26433 12393 26467 12427
rect 27813 12393 27847 12427
rect 28825 12393 28859 12427
rect 29561 12393 29595 12427
rect 33241 12393 33275 12427
rect 42901 12393 42935 12427
rect 16957 12325 16991 12359
rect 29009 12325 29043 12359
rect 4721 12257 4755 12291
rect 9965 12257 9999 12291
rect 11069 12257 11103 12291
rect 12541 12257 12575 12291
rect 15761 12257 15795 12291
rect 16037 12257 16071 12291
rect 16246 12257 16280 12291
rect 18153 12257 18187 12291
rect 19809 12257 19843 12291
rect 20913 12257 20947 12291
rect 27077 12257 27111 12291
rect 33885 12257 33919 12291
rect 36185 12257 36219 12291
rect 36553 12257 36587 12291
rect 40326 12257 40360 12291
rect 40509 12257 40543 12291
rect 41061 12257 41095 12291
rect 2605 12189 2639 12223
rect 4169 12189 4203 12223
rect 6653 12189 6687 12223
rect 8401 12189 8435 12223
rect 10793 12189 10827 12223
rect 13001 12189 13035 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 14841 12189 14875 12223
rect 16129 12189 16163 12223
rect 16865 12189 16899 12223
rect 17877 12189 17911 12223
rect 19625 12189 19659 12223
rect 20545 12189 20579 12223
rect 23213 12189 23247 12223
rect 23857 12189 23891 12223
rect 25421 12189 25455 12223
rect 25513 12189 25547 12223
rect 26893 12189 26927 12223
rect 27721 12189 27755 12223
rect 28641 12189 28675 12223
rect 28733 12189 28767 12223
rect 29745 12189 29779 12223
rect 30021 12189 30055 12223
rect 31033 12189 31067 12223
rect 33609 12189 33643 12223
rect 33701 12189 33735 12223
rect 36369 12189 36403 12223
rect 37013 12189 37047 12223
rect 39037 12189 39071 12223
rect 39221 12189 39255 12223
rect 39313 12189 39347 12223
rect 40234 12189 40268 12223
rect 40417 12189 40451 12223
rect 42901 12189 42935 12223
rect 43085 12189 43119 12223
rect 4988 12121 5022 12155
rect 9781 12121 9815 12155
rect 24409 12121 24443 12155
rect 25237 12121 25271 12155
rect 31309 12121 31343 12155
rect 37280 12121 37314 12155
rect 38853 12121 38887 12155
rect 41306 12121 41340 12155
rect 3249 12053 3283 12087
rect 3985 12053 4019 12087
rect 7205 12053 7239 12087
rect 8217 12053 8251 12087
rect 9413 12053 9447 12087
rect 9873 12053 9907 12087
rect 13185 12053 13219 12087
rect 16405 12053 16439 12087
rect 17509 12053 17543 12087
rect 17969 12053 18003 12087
rect 19257 12053 19291 12087
rect 19717 12053 19751 12087
rect 23029 12053 23063 12087
rect 24609 12053 24643 12087
rect 24777 12053 24811 12087
rect 26801 12053 26835 12087
rect 29929 12053 29963 12087
rect 32781 12053 32815 12087
rect 38393 12053 38427 12087
rect 40049 12053 40083 12087
rect 42441 12053 42475 12087
rect 4445 11849 4479 11883
rect 5089 11849 5123 11883
rect 5457 11849 5491 11883
rect 5549 11849 5583 11883
rect 13461 11849 13495 11883
rect 17049 11849 17083 11883
rect 19625 11849 19659 11883
rect 20453 11849 20487 11883
rect 21189 11849 21223 11883
rect 22661 11849 22695 11883
rect 26985 11849 27019 11883
rect 28365 11849 28399 11883
rect 29929 11849 29963 11883
rect 30665 11849 30699 11883
rect 33241 11849 33275 11883
rect 33977 11849 34011 11883
rect 34713 11849 34747 11883
rect 37289 11849 37323 11883
rect 38307 11849 38341 11883
rect 9229 11781 9263 11815
rect 11989 11781 12023 11815
rect 23857 11781 23891 11815
rect 24073 11781 24107 11815
rect 29653 11781 29687 11815
rect 39313 11781 39347 11815
rect 40233 11781 40267 11815
rect 3065 11713 3099 11747
rect 3332 11713 3366 11747
rect 6745 11713 6779 11747
rect 12081 11713 12115 11747
rect 14381 11713 14415 11747
rect 15209 11713 15243 11747
rect 17233 11713 17267 11747
rect 20361 11713 20395 11747
rect 21097 11713 21131 11747
rect 21833 11713 21867 11747
rect 22569 11713 22603 11747
rect 23213 11713 23247 11747
rect 23397 11713 23431 11747
rect 24685 11713 24719 11747
rect 27169 11713 27203 11747
rect 27629 11713 27663 11747
rect 28273 11713 28307 11747
rect 29377 11713 29411 11747
rect 29561 11713 29595 11747
rect 29745 11713 29779 11747
rect 30941 11713 30975 11747
rect 32597 11713 32631 11747
rect 33425 11713 33459 11747
rect 33885 11713 33919 11747
rect 34621 11713 34655 11747
rect 36553 11713 36587 11747
rect 36737 11713 36771 11747
rect 37473 11713 37507 11747
rect 37749 11713 37783 11747
rect 38209 11713 38243 11747
rect 38393 11713 38427 11747
rect 38485 11713 38519 11747
rect 38945 11713 38979 11747
rect 39038 11713 39072 11747
rect 39221 11713 39255 11747
rect 39410 11713 39444 11747
rect 40325 11713 40359 11747
rect 40417 11713 40451 11747
rect 40601 11713 40635 11747
rect 41061 11713 41095 11747
rect 5733 11645 5767 11679
rect 7481 11645 7515 11679
rect 8953 11645 8987 11679
rect 10701 11645 10735 11679
rect 12265 11645 12299 11679
rect 12817 11645 12851 11679
rect 15301 11645 15335 11679
rect 15485 11645 15519 11679
rect 17877 11645 17911 11679
rect 18153 11645 18187 11679
rect 24961 11645 24995 11679
rect 26433 11645 26467 11679
rect 27721 11645 27755 11679
rect 30849 11645 30883 11679
rect 31217 11645 31251 11679
rect 31309 11645 31343 11679
rect 36645 11645 36679 11679
rect 42441 11645 42475 11679
rect 42717 11645 42751 11679
rect 6561 11577 6595 11611
rect 11621 11577 11655 11611
rect 14841 11577 14875 11611
rect 24225 11577 24259 11611
rect 40049 11577 40083 11611
rect 8033 11509 8067 11543
rect 14197 11509 14231 11543
rect 22017 11509 22051 11543
rect 23305 11509 23339 11543
rect 24041 11509 24075 11543
rect 32689 11509 32723 11543
rect 37657 11509 37691 11543
rect 39589 11509 39623 11543
rect 41153 11509 41187 11543
rect 41521 11509 41555 11543
rect 2513 11305 2547 11339
rect 8217 11305 8251 11339
rect 10333 11305 10367 11339
rect 12817 11305 12851 11339
rect 15945 11305 15979 11339
rect 17877 11305 17911 11339
rect 18613 11305 18647 11339
rect 20729 11305 20763 11339
rect 26157 11305 26191 11339
rect 30665 11305 30699 11339
rect 31033 11305 31067 11339
rect 41061 11305 41095 11339
rect 42073 11305 42107 11339
rect 7757 11237 7791 11271
rect 10793 11237 10827 11271
rect 12357 11237 12391 11271
rect 27261 11237 27295 11271
rect 31493 11237 31527 11271
rect 37197 11237 37231 11271
rect 39313 11237 39347 11271
rect 2973 11169 3007 11203
rect 3157 11169 3191 11203
rect 11437 11169 11471 11203
rect 13461 11169 13495 11203
rect 14197 11169 14231 11203
rect 22661 11169 22695 11203
rect 26341 11169 26375 11203
rect 26709 11169 26743 11203
rect 34115 11169 34149 11203
rect 34713 11169 34747 11203
rect 37933 11169 37967 11203
rect 41521 11169 41555 11203
rect 4353 11101 4387 11135
rect 4620 11101 4654 11135
rect 6377 11101 6411 11135
rect 8401 11101 8435 11135
rect 8953 11101 8987 11135
rect 11161 11101 11195 11135
rect 12173 11101 12207 11135
rect 13277 11101 13311 11135
rect 16681 11101 16715 11135
rect 18061 11101 18095 11135
rect 18521 11101 18555 11135
rect 19349 11101 19383 11135
rect 22477 11101 22511 11135
rect 22569 11101 22603 11135
rect 23857 11101 23891 11135
rect 24961 11101 24995 11135
rect 25237 11101 25271 11135
rect 26433 11101 26467 11135
rect 27445 11101 27479 11135
rect 30021 11101 30055 11135
rect 30665 11101 30699 11135
rect 30757 11101 30791 11135
rect 31493 11101 31527 11135
rect 32321 11101 32355 11135
rect 32689 11101 32723 11135
rect 34989 11101 35023 11135
rect 36553 11101 36587 11135
rect 36737 11101 36771 11135
rect 37473 11101 37507 11135
rect 39865 11101 39899 11135
rect 40049 11101 40083 11135
rect 40141 11101 40175 11135
rect 40233 11101 40267 11135
rect 40417 11101 40451 11135
rect 41245 11101 41279 11135
rect 41429 11101 41463 11135
rect 41981 11101 42015 11135
rect 42809 11101 42843 11135
rect 43453 11101 43487 11135
rect 43637 11101 43671 11135
rect 2881 11033 2915 11067
rect 6644 11033 6678 11067
rect 9198 11033 9232 11067
rect 11253 11033 11287 11067
rect 13185 11033 13219 11067
rect 14473 11033 14507 11067
rect 19616 11033 19650 11067
rect 26801 11033 26835 11067
rect 30113 11033 30147 11067
rect 37197 11033 37231 11067
rect 37381 11033 37415 11067
rect 38178 11033 38212 11067
rect 42625 11033 42659 11067
rect 5733 10965 5767 10999
rect 16497 10965 16531 10999
rect 22109 10965 22143 10999
rect 23673 10965 23707 10999
rect 24777 10965 24811 10999
rect 25145 10965 25179 10999
rect 36737 10965 36771 10999
rect 40601 10965 40635 10999
rect 42993 10965 43027 10999
rect 43545 10965 43579 10999
rect 3249 10761 3283 10795
rect 7113 10761 7147 10795
rect 14841 10761 14875 10795
rect 15393 10761 15427 10795
rect 22201 10761 22235 10795
rect 26249 10761 26283 10795
rect 35081 10761 35115 10795
rect 7021 10693 7055 10727
rect 13369 10693 13403 10727
rect 24777 10693 24811 10727
rect 33793 10693 33827 10727
rect 38301 10693 38335 10727
rect 42901 10693 42935 10727
rect 1409 10625 1443 10659
rect 2421 10625 2455 10659
rect 3065 10625 3099 10659
rect 3801 10625 3835 10659
rect 4057 10625 4091 10659
rect 7849 10625 7883 10659
rect 10793 10625 10827 10659
rect 11989 10625 12023 10659
rect 13093 10625 13127 10659
rect 15301 10625 15335 10659
rect 16129 10625 16163 10659
rect 17693 10625 17727 10659
rect 21005 10625 21039 10659
rect 23029 10625 23063 10659
rect 24501 10625 24535 10659
rect 28641 10625 28675 10659
rect 30849 10625 30883 10659
rect 32597 10625 32631 10659
rect 32781 10625 32815 10659
rect 32965 10625 32999 10659
rect 33057 10625 33091 10659
rect 36001 10625 36035 10659
rect 37381 10647 37415 10681
rect 38117 10625 38151 10659
rect 38945 10625 38979 10659
rect 40785 10625 40819 10659
rect 40969 10625 41003 10659
rect 41613 10625 41647 10659
rect 42625 10625 42659 10659
rect 42809 10625 42843 10659
rect 42993 10625 43027 10659
rect 44189 10625 44223 10659
rect 2881 10557 2915 10591
rect 7297 10557 7331 10591
rect 10609 10557 10643 10591
rect 11805 10557 11839 10591
rect 12173 10557 12207 10591
rect 22293 10557 22327 10591
rect 22477 10557 22511 10591
rect 30297 10557 30331 10591
rect 37473 10557 37507 10591
rect 37657 10557 37691 10591
rect 39221 10557 39255 10591
rect 40877 10557 40911 10591
rect 41061 10557 41095 10591
rect 10977 10489 11011 10523
rect 21189 10489 21223 10523
rect 36093 10489 36127 10523
rect 37381 10489 37415 10523
rect 43177 10489 43211 10523
rect 1593 10421 1627 10455
rect 2237 10421 2271 10455
rect 5181 10421 5215 10455
rect 6653 10421 6687 10455
rect 9321 10421 9355 10455
rect 15945 10421 15979 10455
rect 17785 10421 17819 10455
rect 21833 10421 21867 10455
rect 23121 10421 23155 10455
rect 30941 10421 30975 10455
rect 38485 10421 38519 10455
rect 40601 10421 40635 10455
rect 41705 10421 41739 10455
rect 5181 10217 5215 10251
rect 8953 10217 8987 10251
rect 11069 10217 11103 10251
rect 14473 10217 14507 10251
rect 15025 10217 15059 10251
rect 19717 10217 19751 10251
rect 22017 10217 22051 10251
rect 22661 10217 22695 10251
rect 23765 10217 23799 10251
rect 25605 10217 25639 10251
rect 33517 10217 33551 10251
rect 35633 10217 35667 10251
rect 36277 10217 36311 10251
rect 39313 10217 39347 10251
rect 40325 10217 40359 10251
rect 40509 10217 40543 10251
rect 43361 10217 43395 10251
rect 41613 10149 41647 10183
rect 9689 10081 9723 10115
rect 12725 10081 12759 10115
rect 14105 10081 14139 10115
rect 15761 10081 15795 10115
rect 17509 10081 17543 10115
rect 20637 10081 20671 10115
rect 29561 10081 29595 10115
rect 31769 10081 31803 10115
rect 37933 10081 37967 10115
rect 2697 10013 2731 10047
rect 3801 10013 3835 10047
rect 6101 10013 6135 10047
rect 9137 10013 9171 10047
rect 11529 10013 11563 10047
rect 12909 10013 12943 10047
rect 14289 10013 14323 10047
rect 14933 10013 14967 10047
rect 18521 10013 18555 10047
rect 19901 10013 19935 10047
rect 22477 10013 22511 10047
rect 23673 10013 23707 10047
rect 24777 10013 24811 10047
rect 25421 10013 25455 10047
rect 26709 10013 26743 10047
rect 26985 10013 27019 10047
rect 27445 10013 27479 10047
rect 28457 10013 28491 10047
rect 34713 10013 34747 10047
rect 34897 10013 34931 10047
rect 35541 10013 35575 10047
rect 36185 10013 36219 10047
rect 37289 10013 37323 10047
rect 37473 10013 37507 10047
rect 40141 10013 40175 10047
rect 40325 10013 40359 10047
rect 40958 10013 40992 10047
rect 41117 10013 41151 10047
rect 41245 10013 41279 10047
rect 41337 10013 41371 10047
rect 41475 10013 41509 10047
rect 42165 10013 42199 10047
rect 42257 10013 42291 10047
rect 42349 10013 42383 10047
rect 42993 10013 43027 10047
rect 4046 9945 4080 9979
rect 9934 9945 9968 9979
rect 16037 9945 16071 9979
rect 20904 9945 20938 9979
rect 26893 9945 26927 9979
rect 29837 9945 29871 9979
rect 32045 9945 32079 9979
rect 38200 9945 38234 9979
rect 39865 9945 39899 9979
rect 42533 9945 42567 9979
rect 43177 9945 43211 9979
rect 3249 9877 3283 9911
rect 7389 9877 7423 9911
rect 12173 9877 12207 9911
rect 13093 9877 13127 9911
rect 18613 9877 18647 9911
rect 24869 9877 24903 9911
rect 26525 9877 26559 9911
rect 27537 9877 27571 9911
rect 28549 9877 28583 9911
rect 31309 9877 31343 9911
rect 35081 9877 35115 9911
rect 37381 9877 37415 9911
rect 5089 9673 5123 9707
rect 11989 9673 12023 9707
rect 20177 9673 20211 9707
rect 25145 9673 25179 9707
rect 25789 9673 25823 9707
rect 31033 9673 31067 9707
rect 32603 9673 32637 9707
rect 33977 9673 34011 9707
rect 38853 9673 38887 9707
rect 41245 9673 41279 9707
rect 42441 9673 42475 9707
rect 3976 9605 4010 9639
rect 9772 9605 9806 9639
rect 11897 9605 11931 9639
rect 14749 9605 14783 9639
rect 23673 9605 23707 9639
rect 35633 9605 35667 9639
rect 38301 9605 38335 9639
rect 38669 9605 38703 9639
rect 40877 9605 40911 9639
rect 43545 9605 43579 9639
rect 1869 9537 1903 9571
rect 2136 9537 2170 9571
rect 5733 9537 5767 9571
rect 6745 9537 6779 9571
rect 6837 9537 6871 9571
rect 7573 9537 7607 9571
rect 8861 9537 8895 9571
rect 9505 9537 9539 9571
rect 13001 9537 13035 9571
rect 15761 9537 15795 9571
rect 16681 9537 16715 9571
rect 17509 9537 17543 9571
rect 20821 9537 20855 9571
rect 25605 9537 25639 9571
rect 29920 9537 29954 9571
rect 32689 9537 32723 9571
rect 32781 9537 32815 9571
rect 33057 9537 33091 9571
rect 33885 9537 33919 9571
rect 34897 9537 34931 9571
rect 35817 9537 35851 9571
rect 35909 9537 35943 9571
rect 36369 9537 36403 9571
rect 36553 9537 36587 9571
rect 38485 9537 38519 9571
rect 38577 9537 38611 9571
rect 40601 9537 40635 9571
rect 40694 9537 40728 9571
rect 40969 9537 41003 9571
rect 41107 9537 41141 9571
rect 41705 9537 41739 9571
rect 41889 9537 41923 9571
rect 42625 9537 42659 9571
rect 42717 9537 42751 9571
rect 42993 9537 43027 9571
rect 43453 9537 43487 9571
rect 43637 9537 43671 9571
rect 3709 9469 3743 9503
rect 6929 9469 6963 9503
rect 12081 9469 12115 9503
rect 15853 9469 15887 9503
rect 15945 9469 15979 9503
rect 17785 9469 17819 9503
rect 19717 9469 19751 9503
rect 20637 9469 20671 9503
rect 21833 9469 21867 9503
rect 22109 9469 22143 9503
rect 23397 9469 23431 9503
rect 27445 9469 27479 9503
rect 27721 9469 27755 9503
rect 29653 9469 29687 9503
rect 32965 9469 32999 9503
rect 34069 9469 34103 9503
rect 35173 9469 35207 9503
rect 36461 9469 36495 9503
rect 39313 9469 39347 9503
rect 42901 9469 42935 9503
rect 3249 9401 3283 9435
rect 6377 9401 6411 9435
rect 15393 9401 15427 9435
rect 19257 9401 19291 9435
rect 19993 9401 20027 9435
rect 33517 9401 33551 9435
rect 39543 9401 39577 9435
rect 5549 9333 5583 9367
rect 8217 9333 8251 9367
rect 8677 9333 8711 9367
rect 10885 9333 10919 9367
rect 11529 9333 11563 9367
rect 16773 9333 16807 9367
rect 21005 9333 21039 9367
rect 29193 9333 29227 9367
rect 32321 9333 32355 9367
rect 34713 9333 34747 9367
rect 35081 9333 35115 9367
rect 35909 9333 35943 9367
rect 41705 9333 41739 9367
rect 5825 9129 5859 9163
rect 11989 9129 12023 9163
rect 27813 9129 27847 9163
rect 30389 9129 30423 9163
rect 35081 9129 35115 9163
rect 37381 9129 37415 9163
rect 38209 9129 38243 9163
rect 38853 9129 38887 9163
rect 40233 9129 40267 9163
rect 42993 9129 43027 9163
rect 43453 9129 43487 9163
rect 6285 9061 6319 9095
rect 17049 9061 17083 9095
rect 21189 9061 21223 9095
rect 31769 9061 31803 9095
rect 38393 9061 38427 9095
rect 39221 9061 39255 9095
rect 42165 9061 42199 9095
rect 3157 8993 3191 9027
rect 6745 8993 6779 9027
rect 6837 8993 6871 9027
rect 9137 8993 9171 9027
rect 13461 8993 13495 9027
rect 14657 8993 14691 9027
rect 15301 8993 15335 9027
rect 19717 8993 19751 9027
rect 23857 8993 23891 9027
rect 30665 8993 30699 9027
rect 31861 8993 31895 9027
rect 32781 8993 32815 9027
rect 35173 8993 35207 9027
rect 40785 8993 40819 9027
rect 2881 8925 2915 8959
rect 3985 8925 4019 8959
rect 4445 8925 4479 8959
rect 6653 8925 6687 8959
rect 7665 8925 7699 8959
rect 7849 8925 7883 8959
rect 9413 8925 9447 8959
rect 10609 8925 10643 8959
rect 13185 8925 13219 8959
rect 14565 8925 14599 8959
rect 19441 8925 19475 8959
rect 24409 8925 24443 8959
rect 24593 8925 24627 8959
rect 24777 8925 24811 8959
rect 25421 8925 25455 8959
rect 26065 8925 26099 8959
rect 28825 8925 28859 8959
rect 29009 8925 29043 8959
rect 29745 8925 29779 8959
rect 30573 8925 30607 8959
rect 30757 8925 30791 8959
rect 30849 8925 30883 8959
rect 31585 8925 31619 8959
rect 33048 8925 33082 8959
rect 34897 8925 34931 8959
rect 37565 8925 37599 8959
rect 39037 8925 39071 8959
rect 39313 8925 39347 8959
rect 40049 8925 40083 8959
rect 40325 8925 40359 8959
rect 42625 8925 42659 8959
rect 42809 8925 42843 8959
rect 43637 8925 43671 8959
rect 4690 8857 4724 8891
rect 10876 8857 10910 8891
rect 14473 8857 14507 8891
rect 15577 8857 15611 8891
rect 22109 8857 22143 8891
rect 26341 8857 26375 8891
rect 31401 8857 31435 8891
rect 38025 8857 38059 8891
rect 38241 8857 38275 8891
rect 41030 8857 41064 8891
rect 2513 8789 2547 8823
rect 2973 8789 3007 8823
rect 3801 8789 3835 8823
rect 8033 8789 8067 8823
rect 12817 8789 12851 8823
rect 13277 8789 13311 8823
rect 14105 8789 14139 8823
rect 25237 8789 25271 8823
rect 28917 8789 28951 8823
rect 29837 8789 29871 8823
rect 34161 8789 34195 8823
rect 34713 8789 34747 8823
rect 39865 8789 39899 8823
rect 1409 8585 1443 8619
rect 3065 8585 3099 8619
rect 4905 8585 4939 8619
rect 7527 8585 7561 8619
rect 10609 8585 10643 8619
rect 13093 8585 13127 8619
rect 13553 8585 13587 8619
rect 13921 8585 13955 8619
rect 16129 8585 16163 8619
rect 19441 8585 19475 8619
rect 25881 8585 25915 8619
rect 27445 8585 27479 8619
rect 38485 8585 38519 8619
rect 40417 8585 40451 8619
rect 44005 8585 44039 8619
rect 14013 8517 14047 8551
rect 22109 8517 22143 8551
rect 28273 8517 28307 8551
rect 28457 8517 28491 8551
rect 42809 8517 42843 8551
rect 1593 8449 1627 8483
rect 2513 8449 2547 8483
rect 3781 8449 3815 8483
rect 5641 8449 5675 8483
rect 6561 8449 6595 8483
rect 7297 8449 7331 8483
rect 8769 8449 8803 8483
rect 9229 8449 9263 8483
rect 9485 8449 9519 8483
rect 11713 8449 11747 8483
rect 11969 8449 12003 8483
rect 14749 8449 14783 8483
rect 15016 8449 15050 8483
rect 18317 8449 18351 8483
rect 20269 8449 20303 8483
rect 21281 8449 21315 8483
rect 24757 8449 24791 8483
rect 27353 8449 27387 8483
rect 29009 8449 29043 8483
rect 29745 8449 29779 8483
rect 29883 8449 29917 8483
rect 30021 8449 30055 8483
rect 30137 8449 30171 8483
rect 31401 8449 31435 8483
rect 32413 8449 32447 8483
rect 33609 8449 33643 8483
rect 33876 8449 33910 8483
rect 37381 8449 37415 8483
rect 38393 8449 38427 8483
rect 38577 8449 38611 8483
rect 39037 8449 39071 8483
rect 39304 8449 39338 8483
rect 40877 8449 40911 8483
rect 42625 8449 42659 8483
rect 43269 8449 43303 8483
rect 44189 8449 44223 8483
rect 3525 8381 3559 8415
rect 5457 8381 5491 8415
rect 6377 8381 6411 8415
rect 14197 8381 14231 8415
rect 18061 8381 18095 8415
rect 20361 8381 20395 8415
rect 20499 8381 20533 8415
rect 21833 8381 21867 8415
rect 23581 8381 23615 8415
rect 24501 8381 24535 8415
rect 27537 8381 27571 8415
rect 29193 8381 29227 8415
rect 31217 8381 31251 8415
rect 32229 8381 32263 8415
rect 41153 8381 41187 8415
rect 42441 8381 42475 8415
rect 43361 8381 43395 8415
rect 5825 8313 5859 8347
rect 6745 8313 6779 8347
rect 21097 8313 21131 8347
rect 31585 8313 31619 8347
rect 32597 8313 32631 8347
rect 34989 8313 35023 8347
rect 37473 8313 37507 8347
rect 8585 8245 8619 8279
rect 19901 8245 19935 8279
rect 26985 8245 27019 8279
rect 30297 8245 30331 8279
rect 5365 8041 5399 8075
rect 7849 8041 7883 8075
rect 10793 8041 10827 8075
rect 15577 8041 15611 8075
rect 21097 8041 21131 8075
rect 23857 8041 23891 8075
rect 33977 8041 34011 8075
rect 39129 8041 39163 8075
rect 41245 8041 41279 8075
rect 44005 8041 44039 8075
rect 16037 7973 16071 8007
rect 35357 7973 35391 8007
rect 11897 7905 11931 7939
rect 16589 7905 16623 7939
rect 21741 7905 21775 7939
rect 26433 7905 26467 7939
rect 28825 7905 28859 7939
rect 39865 7905 39899 7939
rect 41705 7905 41739 7939
rect 3985 7837 4019 7871
rect 6469 7837 6503 7871
rect 8953 7837 8987 7871
rect 10977 7837 11011 7871
rect 14197 7837 14231 7871
rect 16497 7837 16531 7871
rect 17417 7837 17451 7871
rect 18705 7837 18739 7871
rect 19257 7837 19291 7871
rect 22477 7837 22511 7871
rect 22744 7837 22778 7871
rect 24593 7837 24627 7871
rect 24860 7837 24894 7871
rect 29745 7837 29779 7871
rect 30012 7837 30046 7871
rect 32137 7837 32171 7871
rect 32404 7837 32438 7871
rect 33977 7837 34011 7871
rect 34161 7837 34195 7871
rect 34897 7837 34931 7871
rect 35541 7837 35575 7871
rect 39129 7837 39163 7871
rect 39313 7837 39347 7871
rect 41889 7837 41923 7871
rect 44189 7837 44223 7871
rect 4252 7769 4286 7803
rect 6714 7769 6748 7803
rect 9198 7769 9232 7803
rect 12142 7769 12176 7803
rect 14464 7769 14498 7803
rect 19502 7769 19536 7803
rect 26678 7769 26712 7803
rect 28641 7769 28675 7803
rect 40110 7769 40144 7803
rect 10333 7701 10367 7735
rect 13277 7701 13311 7735
rect 16405 7701 16439 7735
rect 17233 7701 17267 7735
rect 18521 7701 18555 7735
rect 20637 7701 20671 7735
rect 21465 7701 21499 7735
rect 21557 7701 21591 7735
rect 25973 7701 26007 7735
rect 27813 7701 27847 7735
rect 28273 7701 28307 7735
rect 28733 7701 28767 7735
rect 31125 7701 31159 7735
rect 33517 7701 33551 7735
rect 34713 7701 34747 7735
rect 42073 7701 42107 7735
rect 3893 7497 3927 7531
rect 10609 7497 10643 7531
rect 12081 7497 12115 7531
rect 14749 7497 14783 7531
rect 15577 7497 15611 7531
rect 17325 7497 17359 7531
rect 19441 7497 19475 7531
rect 22201 7497 22235 7531
rect 22661 7497 22695 7531
rect 24133 7497 24167 7531
rect 26157 7497 26191 7531
rect 27169 7497 27203 7531
rect 27537 7497 27571 7531
rect 29929 7497 29963 7531
rect 39865 7497 39899 7531
rect 40785 7497 40819 7531
rect 2605 7429 2639 7463
rect 7849 7429 7883 7463
rect 9505 7429 9539 7463
rect 10425 7429 10459 7463
rect 10701 7429 10735 7463
rect 12173 7429 12207 7463
rect 17233 7429 17267 7463
rect 26065 7429 26099 7463
rect 13369 7361 13403 7395
rect 13636 7361 13670 7395
rect 18328 7361 18362 7395
rect 19901 7361 19935 7395
rect 20168 7361 20202 7395
rect 22569 7361 22603 7395
rect 23581 7361 23615 7395
rect 24041 7361 24075 7395
rect 25237 7361 25271 7395
rect 27629 7361 27663 7395
rect 28641 7361 28675 7395
rect 30941 7361 30975 7395
rect 32137 7361 32171 7395
rect 33057 7361 33091 7395
rect 39221 7361 39255 7395
rect 39405 7361 39439 7395
rect 40049 7361 40083 7395
rect 40325 7361 40359 7395
rect 40969 7361 41003 7395
rect 41153 7361 41187 7395
rect 41245 7361 41279 7395
rect 12357 7293 12391 7327
rect 15669 7293 15703 7327
rect 15853 7293 15887 7327
rect 17509 7293 17543 7327
rect 18061 7293 18095 7327
rect 22845 7293 22879 7327
rect 26249 7293 26283 7327
rect 27721 7293 27755 7327
rect 33333 7293 33367 7327
rect 39313 7293 39347 7327
rect 15209 7225 15243 7259
rect 25053 7225 25087 7259
rect 40233 7225 40267 7259
rect 1593 7157 1627 7191
rect 10149 7157 10183 7191
rect 11713 7157 11747 7191
rect 16865 7157 16899 7191
rect 21281 7157 21315 7191
rect 23397 7157 23431 7191
rect 25697 7157 25731 7191
rect 31033 7157 31067 7191
rect 32321 7157 32355 7191
rect 34805 7157 34839 7191
rect 16037 6953 16071 6987
rect 18521 6953 18555 6987
rect 23305 6953 23339 6987
rect 26433 6953 26467 6987
rect 28365 6953 28399 6987
rect 30100 6953 30134 6987
rect 40049 6953 40083 6987
rect 8401 6885 8435 6919
rect 9229 6885 9263 6919
rect 7021 6817 7055 6851
rect 13277 6817 13311 6851
rect 13461 6817 13495 6851
rect 19257 6817 19291 6851
rect 21189 6817 21223 6851
rect 21373 6817 21407 6851
rect 26985 6817 27019 6851
rect 29837 6817 29871 6851
rect 32689 6817 32723 6851
rect 6561 6749 6595 6783
rect 9873 6749 9907 6783
rect 10057 6749 10091 6783
rect 10793 6749 10827 6783
rect 14657 6749 14691 6783
rect 16681 6749 16715 6783
rect 18705 6749 18739 6783
rect 19441 6749 19475 6783
rect 21925 6749 21959 6783
rect 25789 6749 25823 6783
rect 27241 6749 27275 6783
rect 32037 6759 32071 6793
rect 32956 6749 32990 6783
rect 40049 6749 40083 6783
rect 40233 6749 40267 6783
rect 7288 6681 7322 6715
rect 8953 6681 8987 6715
rect 10241 6681 10275 6715
rect 11038 6681 11072 6715
rect 13185 6681 13219 6715
rect 14924 6681 14958 6715
rect 19625 6681 19659 6715
rect 22192 6681 22226 6715
rect 26341 6681 26375 6715
rect 6377 6613 6411 6647
rect 9413 6613 9447 6647
rect 12173 6613 12207 6647
rect 12817 6613 12851 6647
rect 16497 6613 16531 6647
rect 20729 6613 20763 6647
rect 21097 6613 21131 6647
rect 25605 6613 25639 6647
rect 31585 6613 31619 6647
rect 32137 6613 32171 6647
rect 34069 6613 34103 6647
rect 8217 6409 8251 6443
rect 8953 6409 8987 6443
rect 11529 6409 11563 6443
rect 17509 6409 17543 6443
rect 17969 6409 18003 6443
rect 21097 6409 21131 6443
rect 30849 6409 30883 6443
rect 31217 6409 31251 6443
rect 34713 6409 34747 6443
rect 35909 6409 35943 6443
rect 12510 6341 12544 6375
rect 14832 6341 14866 6375
rect 26341 6341 26375 6375
rect 35265 6341 35299 6375
rect 6377 6273 6411 6307
rect 6633 6273 6667 6307
rect 8401 6273 8435 6307
rect 9137 6273 9171 6307
rect 9597 6273 9631 6307
rect 9864 6273 9898 6307
rect 11713 6273 11747 6307
rect 12265 6273 12299 6307
rect 14565 6273 14599 6307
rect 17049 6273 17083 6307
rect 17877 6273 17911 6307
rect 21281 6273 21315 6307
rect 21833 6273 21867 6307
rect 22089 6273 22123 6307
rect 23857 6273 23891 6307
rect 26249 6273 26283 6307
rect 26985 6273 27019 6307
rect 29561 6273 29595 6307
rect 31309 6273 31343 6307
rect 32137 6273 32171 6307
rect 32321 6273 32355 6307
rect 32965 6273 32999 6307
rect 35173 6273 35207 6307
rect 35817 6273 35851 6307
rect 18061 6205 18095 6239
rect 23765 6205 23799 6239
rect 27261 6205 27295 6239
rect 29837 6205 29871 6239
rect 31401 6205 31435 6239
rect 33241 6205 33275 6239
rect 7757 6137 7791 6171
rect 10977 6069 11011 6103
rect 13645 6069 13679 6103
rect 15945 6069 15979 6103
rect 16865 6069 16899 6103
rect 23213 6069 23247 6103
rect 24225 6069 24259 6103
rect 28733 6069 28767 6103
rect 32505 6069 32539 6103
rect 8309 5865 8343 5899
rect 11713 5865 11747 5899
rect 15761 5865 15795 5899
rect 18337 5865 18371 5899
rect 24409 5865 24443 5899
rect 26893 5865 26927 5899
rect 34713 5865 34747 5899
rect 35357 5865 35391 5899
rect 9781 5797 9815 5831
rect 12817 5797 12851 5831
rect 14749 5797 14783 5831
rect 13369 5729 13403 5763
rect 15393 5729 15427 5763
rect 19349 5729 19383 5763
rect 19809 5729 19843 5763
rect 22937 5729 22971 5763
rect 23397 5729 23431 5763
rect 24501 5729 24535 5763
rect 29745 5729 29779 5763
rect 32781 5729 32815 5763
rect 6929 5661 6963 5695
rect 9137 5661 9171 5695
rect 9965 5661 9999 5695
rect 10425 5661 10459 5695
rect 13185 5661 13219 5695
rect 15577 5661 15611 5695
rect 16957 5661 16991 5695
rect 19441 5661 19475 5695
rect 21833 5661 21867 5695
rect 23029 5661 23063 5695
rect 24409 5661 24443 5695
rect 24685 5661 24719 5695
rect 26433 5661 26467 5695
rect 27077 5661 27111 5695
rect 27721 5661 27755 5695
rect 27813 5661 27847 5695
rect 28457 5661 28491 5695
rect 28733 5661 28767 5695
rect 29837 5661 29871 5695
rect 29929 5661 29963 5695
rect 30021 5661 30055 5695
rect 31217 5661 31251 5695
rect 33425 5661 33459 5695
rect 33609 5661 33643 5695
rect 34897 5661 34931 5695
rect 35541 5661 35575 5695
rect 36185 5661 36219 5695
rect 43913 5661 43947 5695
rect 7196 5593 7230 5627
rect 14565 5593 14599 5627
rect 17202 5593 17236 5627
rect 27537 5593 27571 5627
rect 8953 5525 8987 5559
rect 13277 5525 13311 5559
rect 22017 5525 22051 5559
rect 24869 5525 24903 5559
rect 26249 5525 26283 5559
rect 27813 5525 27847 5559
rect 28273 5525 28307 5559
rect 28641 5525 28675 5559
rect 29561 5525 29595 5559
rect 33517 5525 33551 5559
rect 36001 5525 36035 5559
rect 44097 5525 44131 5559
rect 10977 5321 11011 5355
rect 11805 5321 11839 5355
rect 12265 5321 12299 5355
rect 18797 5321 18831 5355
rect 19625 5321 19659 5355
rect 19717 5321 19751 5355
rect 8024 5253 8058 5287
rect 13001 5253 13035 5287
rect 17684 5253 17718 5287
rect 23949 5253 23983 5287
rect 25421 5253 25455 5287
rect 27997 5253 28031 5287
rect 28457 5253 28491 5287
rect 28657 5253 28691 5287
rect 30573 5253 30607 5287
rect 30849 5253 30883 5287
rect 30941 5253 30975 5287
rect 31125 5253 31159 5287
rect 32321 5253 32355 5287
rect 35817 5253 35851 5287
rect 7757 5185 7791 5219
rect 10149 5185 10183 5219
rect 10793 5185 10827 5219
rect 12173 5185 12207 5219
rect 15393 5185 15427 5219
rect 17417 5185 17451 5219
rect 20453 5185 20487 5219
rect 20729 5185 20763 5219
rect 22109 5185 22143 5219
rect 23121 5185 23155 5219
rect 24133 5185 24167 5219
rect 25053 5185 25087 5219
rect 25145 5185 25179 5219
rect 25329 5185 25363 5219
rect 25513 5185 25547 5219
rect 27077 5185 27111 5219
rect 27261 5185 27295 5219
rect 27813 5185 27847 5219
rect 30757 5185 30791 5219
rect 32137 5185 32171 5219
rect 33425 5185 33459 5219
rect 35725 5185 35759 5219
rect 42993 5185 43027 5219
rect 43269 5185 43303 5219
rect 1409 5117 1443 5151
rect 1685 5117 1719 5151
rect 10609 5117 10643 5151
rect 12357 5117 12391 5151
rect 14749 5117 14783 5151
rect 19901 5117 19935 5151
rect 20545 5117 20579 5151
rect 22201 5117 22235 5151
rect 23029 5117 23063 5151
rect 23489 5117 23523 5151
rect 27169 5117 27203 5151
rect 29285 5117 29319 5151
rect 29561 5117 29595 5151
rect 33701 5117 33735 5151
rect 9965 5049 9999 5083
rect 22477 5049 22511 5083
rect 28825 5049 28859 5083
rect 9137 4981 9171 5015
rect 15209 4981 15243 5015
rect 19257 4981 19291 5015
rect 20453 4981 20487 5015
rect 20913 4981 20947 5015
rect 24317 4981 24351 5015
rect 25053 4981 25087 5015
rect 28641 4981 28675 5015
rect 32505 4981 32539 5015
rect 35173 4981 35207 5015
rect 42809 4981 42843 5015
rect 14105 4777 14139 4811
rect 17509 4777 17543 4811
rect 19809 4777 19843 4811
rect 22096 4777 22130 4811
rect 24869 4777 24903 4811
rect 25053 4777 25087 4811
rect 25605 4777 25639 4811
rect 26801 4777 26835 4811
rect 28641 4777 28675 4811
rect 31309 4777 31343 4811
rect 31953 4777 31987 4811
rect 32137 4777 32171 4811
rect 32781 4777 32815 4811
rect 32965 4777 32999 4811
rect 33609 4777 33643 4811
rect 33793 4777 33827 4811
rect 10333 4709 10367 4743
rect 18705 4709 18739 4743
rect 11529 4641 11563 4675
rect 12173 4641 12207 4675
rect 14749 4641 14783 4675
rect 18245 4641 18279 4675
rect 19349 4641 19383 4675
rect 21833 4641 21867 4675
rect 29561 4641 29595 4675
rect 10517 4573 10551 4607
rect 14289 4573 14323 4607
rect 15016 4573 15050 4607
rect 17693 4573 17727 4607
rect 18337 4573 18371 4607
rect 19441 4573 19475 4607
rect 25513 4573 25547 4607
rect 27445 4573 27479 4607
rect 43913 4573 43947 4607
rect 11345 4505 11379 4539
rect 12440 4505 12474 4539
rect 24685 4505 24719 4539
rect 24901 4505 24935 4539
rect 26617 4505 26651 4539
rect 26833 4505 26867 4539
rect 27629 4505 27663 4539
rect 28457 4505 28491 4539
rect 28673 4505 28707 4539
rect 29837 4505 29871 4539
rect 31769 4505 31803 4539
rect 31969 4505 32003 4539
rect 32597 4505 32631 4539
rect 33425 4505 33459 4539
rect 33625 4505 33659 4539
rect 10977 4437 11011 4471
rect 11437 4437 11471 4471
rect 13553 4437 13587 4471
rect 16129 4437 16163 4471
rect 23581 4437 23615 4471
rect 26985 4437 27019 4471
rect 27813 4437 27847 4471
rect 28825 4437 28859 4471
rect 32797 4437 32831 4471
rect 44097 4437 44131 4471
rect 14749 4233 14783 4267
rect 15117 4233 15151 4267
rect 15209 4233 15243 4267
rect 26157 4233 26191 4267
rect 29929 4233 29963 4267
rect 11897 4097 11931 4131
rect 12153 4097 12187 4131
rect 17417 4097 17451 4131
rect 18245 4097 18279 4131
rect 19073 4097 19107 4131
rect 24317 4097 24351 4131
rect 24501 4097 24535 4131
rect 24961 4097 24995 4131
rect 25145 4097 25179 4131
rect 26065 4097 26099 4131
rect 26249 4097 26283 4131
rect 27261 4097 27295 4131
rect 29745 4097 29779 4131
rect 30021 4097 30055 4131
rect 31217 4097 31251 4131
rect 32137 4097 32171 4131
rect 15393 4029 15427 4063
rect 18153 4029 18187 4063
rect 18613 4029 18647 4063
rect 22109 4029 22143 4063
rect 22385 4029 22419 4063
rect 27537 4029 27571 4063
rect 29009 4029 29043 4063
rect 31125 4029 31159 4063
rect 32413 4029 32447 4063
rect 13277 3961 13311 3995
rect 31585 3961 31619 3995
rect 16957 3893 16991 3927
rect 17509 3893 17543 3927
rect 19165 3893 19199 3927
rect 23857 3893 23891 3927
rect 24317 3893 24351 3927
rect 25053 3893 25087 3927
rect 29561 3893 29595 3927
rect 33885 3893 33919 3927
rect 11529 3689 11563 3723
rect 23581 3689 23615 3723
rect 23765 3689 23799 3723
rect 24501 3689 24535 3723
rect 27261 3689 27295 3723
rect 28089 3689 28123 3723
rect 28825 3689 28859 3723
rect 29561 3689 29595 3723
rect 30297 3689 30331 3723
rect 31033 3689 31067 3723
rect 31861 3689 31895 3723
rect 12173 3621 12207 3655
rect 29009 3621 29043 3655
rect 12633 3553 12667 3587
rect 12725 3553 12759 3587
rect 16773 3553 16807 3587
rect 19257 3553 19291 3587
rect 1593 3485 1627 3519
rect 11713 3485 11747 3519
rect 12541 3485 12575 3519
rect 15761 3485 15795 3519
rect 15853 3485 15887 3519
rect 16405 3485 16439 3519
rect 19625 3485 19659 3519
rect 21051 3485 21085 3519
rect 22201 3485 22235 3519
rect 24409 3485 24443 3519
rect 27445 3485 27479 3519
rect 27997 3485 28031 3519
rect 29561 3485 29595 3519
rect 30473 3481 30507 3515
rect 30941 3485 30975 3519
rect 31769 3485 31803 3519
rect 31953 3485 31987 3519
rect 44189 3485 44223 3519
rect 23397 3417 23431 3451
rect 23613 3417 23647 3451
rect 28641 3417 28675 3451
rect 28846 3417 28880 3451
rect 18199 3349 18233 3383
rect 22385 3349 22419 3383
rect 16037 3145 16071 3179
rect 17233 3145 17267 3179
rect 19579 3145 19613 3179
rect 20177 3145 20211 3179
rect 23029 3145 23063 3179
rect 23581 3145 23615 3179
rect 31401 3145 31435 3179
rect 34069 3145 34103 3179
rect 43269 3145 43303 3179
rect 43913 3145 43947 3179
rect 6561 3009 6595 3043
rect 12909 3009 12943 3043
rect 15945 3009 15979 3043
rect 17141 3009 17175 3043
rect 17785 3009 17819 3043
rect 18153 3009 18187 3043
rect 20085 3009 20119 3043
rect 22109 3009 22143 3043
rect 22937 3009 22971 3043
rect 23765 3009 23799 3043
rect 31309 3009 31343 3043
rect 34529 3009 34563 3043
rect 43453 3009 43487 3043
rect 44097 3009 44131 3043
rect 1593 2805 1627 2839
rect 6377 2805 6411 2839
rect 13093 2805 13127 2839
rect 21925 2805 21959 2839
rect 34345 2805 34379 2839
rect 13001 2601 13035 2635
rect 25881 2601 25915 2635
rect 37289 2601 37323 2635
rect 43085 2533 43119 2567
rect 2237 2465 2271 2499
rect 17785 2465 17819 2499
rect 1593 2397 1627 2431
rect 3985 2397 4019 2431
rect 4813 2397 4847 2431
rect 6561 2397 6595 2431
rect 8033 2397 8067 2431
rect 9781 2397 9815 2431
rect 11713 2397 11747 2431
rect 13185 2397 13219 2431
rect 14473 2397 14507 2431
rect 15485 2397 15519 2431
rect 17509 2397 17543 2431
rect 19625 2397 19659 2431
rect 20913 2397 20947 2431
rect 22661 2397 22695 2431
rect 24593 2397 24627 2431
rect 26065 2397 26099 2431
rect 27169 2397 27203 2431
rect 29745 2397 29779 2431
rect 30573 2397 30607 2431
rect 35541 2397 35575 2431
rect 37473 2397 37507 2431
rect 38945 2397 38979 2431
rect 40233 2397 40267 2431
rect 43913 2397 43947 2431
rect 32597 2329 32631 2363
rect 42901 2329 42935 2363
rect 6745 2261 6779 2295
rect 9965 2261 9999 2295
rect 14289 2261 14323 2295
rect 22845 2261 22879 2295
rect 27353 2261 27387 2295
rect 32689 2261 32723 2295
rect 35725 2261 35759 2295
rect 44097 2261 44131 2295
<< metal1 >>
rect 1104 17434 45056 17456
rect 1104 17382 11898 17434
rect 11950 17382 11962 17434
rect 12014 17382 12026 17434
rect 12078 17382 12090 17434
rect 12142 17382 12154 17434
rect 12206 17382 22846 17434
rect 22898 17382 22910 17434
rect 22962 17382 22974 17434
rect 23026 17382 23038 17434
rect 23090 17382 23102 17434
rect 23154 17382 33794 17434
rect 33846 17382 33858 17434
rect 33910 17382 33922 17434
rect 33974 17382 33986 17434
rect 34038 17382 34050 17434
rect 34102 17382 44742 17434
rect 44794 17382 44806 17434
rect 44858 17382 44870 17434
rect 44922 17382 44934 17434
rect 44986 17382 44998 17434
rect 45050 17382 45056 17434
rect 1104 17360 45056 17382
rect 17402 17280 17408 17332
rect 17460 17320 17466 17332
rect 17681 17323 17739 17329
rect 17681 17320 17693 17323
rect 17460 17292 17693 17320
rect 17460 17280 17466 17292
rect 17681 17289 17693 17292
rect 17727 17289 17739 17323
rect 17681 17283 17739 17289
rect 20714 17280 20720 17332
rect 20772 17320 20778 17332
rect 20901 17323 20959 17329
rect 20901 17320 20913 17323
rect 20772 17292 20913 17320
rect 20772 17280 20778 17292
rect 20901 17289 20913 17292
rect 20947 17289 20959 17323
rect 20901 17283 20959 17289
rect 31021 17323 31079 17329
rect 31021 17289 31033 17323
rect 31067 17320 31079 17323
rect 37274 17320 37280 17332
rect 31067 17292 37280 17320
rect 31067 17289 31079 17292
rect 31021 17283 31079 17289
rect 37274 17280 37280 17292
rect 37332 17280 37338 17332
rect 40586 17280 40592 17332
rect 40644 17320 40650 17332
rect 40865 17323 40923 17329
rect 40865 17320 40877 17323
rect 40644 17292 40877 17320
rect 40644 17280 40650 17292
rect 40865 17289 40877 17292
rect 40911 17289 40923 17323
rect 44082 17320 44088 17332
rect 44043 17292 44088 17320
rect 40865 17283 40923 17289
rect 44082 17280 44088 17292
rect 44140 17280 44146 17332
rect 1302 17212 1308 17264
rect 1360 17252 1366 17264
rect 2961 17255 3019 17261
rect 2961 17252 2973 17255
rect 1360 17224 2973 17252
rect 1360 17212 1366 17224
rect 2961 17221 2973 17224
rect 3007 17221 3019 17255
rect 2961 17215 3019 17221
rect 3234 17212 3240 17264
rect 3292 17252 3298 17264
rect 3973 17255 4031 17261
rect 3973 17252 3985 17255
rect 3292 17224 3985 17252
rect 3292 17212 3298 17224
rect 3973 17221 3985 17224
rect 4019 17221 4031 17255
rect 3973 17215 4031 17221
rect 38654 17212 38660 17264
rect 38712 17252 38718 17264
rect 38841 17255 38899 17261
rect 38841 17252 38853 17255
rect 38712 17224 38853 17252
rect 38712 17212 38718 17224
rect 38841 17221 38853 17224
rect 38887 17221 38899 17255
rect 38841 17215 38899 17221
rect 2222 17184 2228 17196
rect 2183 17156 2228 17184
rect 2222 17144 2228 17156
rect 2280 17144 2286 17196
rect 4522 17144 4528 17196
rect 4580 17184 4586 17196
rect 4617 17187 4675 17193
rect 4617 17184 4629 17187
rect 4580 17156 4629 17184
rect 4580 17144 4586 17156
rect 4617 17153 4629 17156
rect 4663 17153 4675 17187
rect 4617 17147 4675 17153
rect 6454 17144 6460 17196
rect 6512 17184 6518 17196
rect 6733 17187 6791 17193
rect 6733 17184 6745 17187
rect 6512 17156 6745 17184
rect 6512 17144 6518 17156
rect 6733 17153 6745 17156
rect 6779 17153 6791 17187
rect 6733 17147 6791 17153
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7800 17156 8033 17184
rect 7800 17144 7806 17156
rect 8021 17153 8033 17156
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9732 17156 9965 17184
rect 9732 17144 9738 17156
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 11112 17156 11529 17184
rect 11112 17144 11118 17156
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 12894 17144 12900 17196
rect 12952 17184 12958 17196
rect 13173 17187 13231 17193
rect 13173 17184 13185 17187
rect 12952 17156 13185 17184
rect 12952 17144 12958 17156
rect 13173 17153 13185 17156
rect 13219 17153 13231 17187
rect 13173 17147 13231 17153
rect 14182 17144 14188 17196
rect 14240 17184 14246 17196
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14240 17156 14473 17184
rect 14240 17144 14246 17156
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 14461 17147 14519 17153
rect 16114 17144 16120 17196
rect 16172 17184 16178 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 16172 17156 16681 17184
rect 16172 17144 16178 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 16758 17144 16764 17196
rect 16816 17184 16822 17196
rect 17497 17187 17555 17193
rect 17497 17184 17509 17187
rect 16816 17156 17509 17184
rect 16816 17144 16822 17156
rect 17497 17153 17509 17156
rect 17543 17153 17555 17187
rect 17497 17147 17555 17153
rect 19334 17144 19340 17196
rect 19392 17184 19398 17196
rect 19613 17187 19671 17193
rect 19613 17184 19625 17187
rect 19392 17156 19625 17184
rect 19392 17144 19398 17156
rect 19613 17153 19625 17156
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17153 20775 17187
rect 20717 17147 20775 17153
rect 2409 17119 2467 17125
rect 2409 17085 2421 17119
rect 2455 17116 2467 17119
rect 4890 17116 4896 17128
rect 2455 17088 4660 17116
rect 4851 17088 4896 17116
rect 2455 17085 2467 17088
rect 2409 17079 2467 17085
rect 4154 17048 4160 17060
rect 4115 17020 4160 17048
rect 4154 17008 4160 17020
rect 4212 17008 4218 17060
rect 4632 17048 4660 17088
rect 4890 17076 4896 17088
rect 4948 17076 4954 17128
rect 11793 17119 11851 17125
rect 11793 17085 11805 17119
rect 11839 17116 11851 17119
rect 17218 17116 17224 17128
rect 11839 17088 17224 17116
rect 11839 17085 11851 17088
rect 11793 17079 11851 17085
rect 17218 17076 17224 17088
rect 17276 17076 17282 17128
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 20732 17116 20760 17147
rect 22554 17144 22560 17196
rect 22612 17184 22618 17196
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 22612 17156 22845 17184
rect 22612 17144 22618 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 23842 17144 23848 17196
rect 23900 17184 23906 17196
rect 24581 17187 24639 17193
rect 24581 17184 24593 17187
rect 23900 17156 24593 17184
rect 23900 17144 23906 17156
rect 24581 17153 24593 17156
rect 24627 17153 24639 17187
rect 24581 17147 24639 17153
rect 25774 17144 25780 17196
rect 25832 17184 25838 17196
rect 26053 17187 26111 17193
rect 26053 17184 26065 17187
rect 25832 17156 26065 17184
rect 25832 17144 25838 17156
rect 26053 17153 26065 17156
rect 26099 17153 26111 17187
rect 26053 17147 26111 17153
rect 27706 17144 27712 17196
rect 27764 17184 27770 17196
rect 27985 17187 28043 17193
rect 27985 17184 27997 17187
rect 27764 17156 27997 17184
rect 27764 17144 27770 17156
rect 27985 17153 27997 17156
rect 28031 17153 28043 17187
rect 27985 17147 28043 17153
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 29733 17187 29791 17193
rect 29733 17184 29745 17187
rect 29052 17156 29745 17184
rect 29052 17144 29058 17156
rect 29733 17153 29745 17156
rect 29779 17153 29791 17187
rect 29733 17147 29791 17153
rect 30926 17144 30932 17196
rect 30984 17184 30990 17196
rect 31205 17187 31263 17193
rect 31205 17184 31217 17187
rect 30984 17156 31217 17184
rect 30984 17144 30990 17156
rect 31205 17153 31217 17156
rect 31251 17153 31263 17187
rect 31205 17147 31263 17153
rect 32214 17144 32220 17196
rect 32272 17184 32278 17196
rect 32309 17187 32367 17193
rect 32309 17184 32321 17187
rect 32272 17156 32321 17184
rect 32272 17144 32278 17156
rect 32309 17153 32321 17156
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 34146 17144 34152 17196
rect 34204 17184 34210 17196
rect 34885 17187 34943 17193
rect 34885 17184 34897 17187
rect 34204 17156 34897 17184
rect 34204 17144 34210 17156
rect 34885 17153 34897 17156
rect 34931 17153 34943 17187
rect 34885 17147 34943 17153
rect 35434 17144 35440 17196
rect 35492 17184 35498 17196
rect 35713 17187 35771 17193
rect 35713 17184 35725 17187
rect 35492 17156 35725 17184
rect 35492 17144 35498 17156
rect 35713 17153 35725 17156
rect 35759 17153 35771 17187
rect 35713 17147 35771 17153
rect 37366 17144 37372 17196
rect 37424 17184 37430 17196
rect 37645 17187 37703 17193
rect 37645 17184 37657 17187
rect 37424 17156 37657 17184
rect 37424 17144 37430 17156
rect 37645 17153 37657 17156
rect 37691 17153 37703 17187
rect 40678 17184 40684 17196
rect 40639 17156 40684 17184
rect 37645 17147 37703 17153
rect 40678 17144 40684 17156
rect 40736 17144 40742 17196
rect 41874 17144 41880 17196
rect 41932 17184 41938 17196
rect 42613 17187 42671 17193
rect 42613 17184 42625 17187
rect 41932 17156 42625 17184
rect 41932 17144 41938 17156
rect 42613 17153 42625 17156
rect 42659 17153 42671 17187
rect 43898 17184 43904 17196
rect 43859 17156 43904 17184
rect 42613 17147 42671 17153
rect 43898 17144 43904 17156
rect 43956 17144 43962 17196
rect 32582 17116 32588 17128
rect 18012 17088 20760 17116
rect 32543 17088 32588 17116
rect 18012 17076 18018 17088
rect 32582 17076 32588 17088
rect 32640 17076 32646 17128
rect 43441 17119 43499 17125
rect 43441 17085 43453 17119
rect 43487 17116 43499 17119
rect 45094 17116 45100 17128
rect 43487 17088 45100 17116
rect 43487 17085 43499 17088
rect 43441 17079 43499 17085
rect 45094 17076 45100 17088
rect 45152 17076 45158 17128
rect 42518 17048 42524 17060
rect 4632 17020 42524 17048
rect 42518 17008 42524 17020
rect 42576 17008 42582 17060
rect 3050 16980 3056 16992
rect 3011 16952 3056 16980
rect 3050 16940 3056 16952
rect 3108 16940 3114 16992
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 9769 16983 9827 16989
rect 9769 16980 9781 16983
rect 9732 16952 9781 16980
rect 9732 16940 9738 16952
rect 9769 16949 9781 16952
rect 9815 16949 9827 16983
rect 16850 16980 16856 16992
rect 16811 16952 16856 16980
rect 9769 16943 9827 16949
rect 16850 16940 16856 16952
rect 16908 16940 16914 16992
rect 23566 16940 23572 16992
rect 23624 16980 23630 16992
rect 24397 16983 24455 16989
rect 24397 16980 24409 16983
rect 23624 16952 24409 16980
rect 23624 16940 23630 16952
rect 24397 16949 24409 16952
rect 24443 16949 24455 16983
rect 24397 16943 24455 16949
rect 34146 16940 34152 16992
rect 34204 16980 34210 16992
rect 34701 16983 34759 16989
rect 34701 16980 34713 16983
rect 34204 16952 34713 16980
rect 34204 16940 34210 16952
rect 34701 16949 34713 16952
rect 34747 16949 34759 16983
rect 38930 16980 38936 16992
rect 38891 16952 38936 16980
rect 34701 16943 34759 16949
rect 38930 16940 38936 16952
rect 38988 16940 38994 16992
rect 1104 16890 44896 16912
rect 1104 16838 6424 16890
rect 6476 16838 6488 16890
rect 6540 16838 6552 16890
rect 6604 16838 6616 16890
rect 6668 16838 6680 16890
rect 6732 16838 17372 16890
rect 17424 16838 17436 16890
rect 17488 16838 17500 16890
rect 17552 16838 17564 16890
rect 17616 16838 17628 16890
rect 17680 16838 28320 16890
rect 28372 16838 28384 16890
rect 28436 16838 28448 16890
rect 28500 16838 28512 16890
rect 28564 16838 28576 16890
rect 28628 16838 39268 16890
rect 39320 16838 39332 16890
rect 39384 16838 39396 16890
rect 39448 16838 39460 16890
rect 39512 16838 39524 16890
rect 39576 16838 44896 16890
rect 1104 16816 44896 16838
rect 3970 16776 3976 16788
rect 3931 16748 3976 16776
rect 3970 16736 3976 16748
rect 4028 16736 4034 16788
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 11698 16776 11704 16788
rect 4948 16748 11704 16776
rect 4948 16736 4954 16748
rect 11698 16736 11704 16748
rect 11756 16736 11762 16788
rect 16850 16736 16856 16788
rect 16908 16776 16914 16788
rect 33686 16776 33692 16788
rect 16908 16748 33692 16776
rect 16908 16736 16914 16748
rect 33686 16736 33692 16748
rect 33744 16736 33750 16788
rect 43438 16776 43444 16788
rect 43399 16748 43444 16776
rect 43438 16736 43444 16748
rect 43496 16736 43502 16788
rect 43806 16736 43812 16788
rect 43864 16776 43870 16788
rect 44085 16779 44143 16785
rect 44085 16776 44097 16779
rect 43864 16748 44097 16776
rect 43864 16736 43870 16748
rect 44085 16745 44097 16748
rect 44131 16745 44143 16779
rect 44085 16739 44143 16745
rect 2041 16711 2099 16717
rect 2041 16677 2053 16711
rect 2087 16708 2099 16711
rect 10686 16708 10692 16720
rect 2087 16680 10692 16708
rect 2087 16677 2099 16680
rect 2041 16671 2099 16677
rect 10686 16668 10692 16680
rect 10744 16668 10750 16720
rect 14 16532 20 16584
rect 72 16572 78 16584
rect 1857 16575 1915 16581
rect 1857 16572 1869 16575
rect 72 16544 1869 16572
rect 72 16532 78 16544
rect 1857 16541 1869 16544
rect 1903 16541 1915 16575
rect 1857 16535 1915 16541
rect 15654 16532 15660 16584
rect 15712 16572 15718 16584
rect 16485 16575 16543 16581
rect 16485 16572 16497 16575
rect 15712 16544 16497 16572
rect 15712 16532 15718 16544
rect 16485 16541 16497 16544
rect 16531 16541 16543 16575
rect 17126 16572 17132 16584
rect 17087 16544 17132 16572
rect 16485 16535 16543 16541
rect 17126 16532 17132 16544
rect 17184 16532 17190 16584
rect 40034 16572 40040 16584
rect 39995 16544 40040 16572
rect 40034 16532 40040 16544
rect 40092 16532 40098 16584
rect 16301 16439 16359 16445
rect 16301 16405 16313 16439
rect 16347 16436 16359 16439
rect 16758 16436 16764 16448
rect 16347 16408 16764 16436
rect 16347 16405 16359 16408
rect 16301 16399 16359 16405
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 16945 16439 17003 16445
rect 16945 16405 16957 16439
rect 16991 16436 17003 16439
rect 17954 16436 17960 16448
rect 16991 16408 17960 16436
rect 16991 16405 17003 16408
rect 16945 16399 17003 16405
rect 17954 16396 17960 16408
rect 18012 16396 18018 16448
rect 39853 16439 39911 16445
rect 39853 16405 39865 16439
rect 39899 16436 39911 16439
rect 40678 16436 40684 16448
rect 39899 16408 40684 16436
rect 39899 16405 39911 16408
rect 39853 16399 39911 16405
rect 40678 16396 40684 16408
rect 40736 16396 40742 16448
rect 1104 16346 45056 16368
rect 1104 16294 11898 16346
rect 11950 16294 11962 16346
rect 12014 16294 12026 16346
rect 12078 16294 12090 16346
rect 12142 16294 12154 16346
rect 12206 16294 22846 16346
rect 22898 16294 22910 16346
rect 22962 16294 22974 16346
rect 23026 16294 23038 16346
rect 23090 16294 23102 16346
rect 23154 16294 33794 16346
rect 33846 16294 33858 16346
rect 33910 16294 33922 16346
rect 33974 16294 33986 16346
rect 34038 16294 34050 16346
rect 34102 16294 44742 16346
rect 44794 16294 44806 16346
rect 44858 16294 44870 16346
rect 44922 16294 44934 16346
rect 44986 16294 44998 16346
rect 45050 16294 45056 16346
rect 1104 16272 45056 16294
rect 44174 15892 44180 15904
rect 44135 15864 44180 15892
rect 44174 15852 44180 15864
rect 44232 15852 44238 15904
rect 1104 15802 44896 15824
rect 1104 15750 6424 15802
rect 6476 15750 6488 15802
rect 6540 15750 6552 15802
rect 6604 15750 6616 15802
rect 6668 15750 6680 15802
rect 6732 15750 17372 15802
rect 17424 15750 17436 15802
rect 17488 15750 17500 15802
rect 17552 15750 17564 15802
rect 17616 15750 17628 15802
rect 17680 15750 28320 15802
rect 28372 15750 28384 15802
rect 28436 15750 28448 15802
rect 28500 15750 28512 15802
rect 28564 15750 28576 15802
rect 28628 15750 39268 15802
rect 39320 15750 39332 15802
rect 39384 15750 39396 15802
rect 39448 15750 39460 15802
rect 39512 15750 39524 15802
rect 39576 15750 44896 15802
rect 1104 15728 44896 15750
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15484 1455 15487
rect 3142 15484 3148 15496
rect 1443 15456 3148 15484
rect 1443 15453 1455 15456
rect 1397 15447 1455 15453
rect 3142 15444 3148 15456
rect 3200 15444 3206 15496
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15484 18567 15487
rect 18598 15484 18604 15496
rect 18555 15456 18604 15484
rect 18555 15453 18567 15456
rect 18509 15447 18567 15453
rect 18598 15444 18604 15456
rect 18656 15444 18662 15496
rect 19150 15444 19156 15496
rect 19208 15484 19214 15496
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 19208 15456 19533 15484
rect 19208 15444 19214 15456
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 34882 15484 34888 15496
rect 34843 15456 34888 15484
rect 19521 15447 19579 15453
rect 34882 15444 34888 15456
rect 34940 15444 34946 15496
rect 19242 15416 19248 15428
rect 19203 15388 19248 15416
rect 19242 15376 19248 15388
rect 19300 15376 19306 15428
rect 19426 15416 19432 15428
rect 19387 15388 19432 15416
rect 19426 15376 19432 15388
rect 19484 15376 19490 15428
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 18046 15308 18052 15360
rect 18104 15348 18110 15360
rect 18325 15351 18383 15357
rect 18325 15348 18337 15351
rect 18104 15320 18337 15348
rect 18104 15308 18110 15320
rect 18325 15317 18337 15320
rect 18371 15348 18383 15351
rect 19150 15348 19156 15360
rect 18371 15320 19156 15348
rect 18371 15317 18383 15320
rect 18325 15311 18383 15317
rect 19150 15308 19156 15320
rect 19208 15308 19214 15360
rect 19518 15348 19524 15360
rect 19479 15320 19524 15348
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 34701 15351 34759 15357
rect 34701 15317 34713 15351
rect 34747 15348 34759 15351
rect 43898 15348 43904 15360
rect 34747 15320 43904 15348
rect 34747 15317 34759 15320
rect 34701 15311 34759 15317
rect 43898 15308 43904 15320
rect 43956 15308 43962 15360
rect 1104 15258 45056 15280
rect 1104 15206 11898 15258
rect 11950 15206 11962 15258
rect 12014 15206 12026 15258
rect 12078 15206 12090 15258
rect 12142 15206 12154 15258
rect 12206 15206 22846 15258
rect 22898 15206 22910 15258
rect 22962 15206 22974 15258
rect 23026 15206 23038 15258
rect 23090 15206 23102 15258
rect 23154 15206 33794 15258
rect 33846 15206 33858 15258
rect 33910 15206 33922 15258
rect 33974 15206 33986 15258
rect 34038 15206 34050 15258
rect 34102 15206 44742 15258
rect 44794 15206 44806 15258
rect 44858 15206 44870 15258
rect 44922 15206 44934 15258
rect 44986 15206 44998 15258
rect 45050 15206 45056 15258
rect 1104 15184 45056 15206
rect 18690 15144 18696 15156
rect 16040 15116 18696 15144
rect 12820 15048 13768 15076
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 15008 8815 15011
rect 8803 14980 8892 15008
rect 8803 14977 8815 14980
rect 8757 14971 8815 14977
rect 8573 14943 8631 14949
rect 8573 14909 8585 14943
rect 8619 14909 8631 14943
rect 8573 14903 8631 14909
rect 8588 14872 8616 14903
rect 8754 14872 8760 14884
rect 8588 14844 8760 14872
rect 8754 14832 8760 14844
rect 8812 14832 8818 14884
rect 8864 14872 8892 14980
rect 12250 14968 12256 15020
rect 12308 15008 12314 15020
rect 12437 15011 12495 15017
rect 12437 15008 12449 15011
rect 12308 14980 12449 15008
rect 12308 14968 12314 14980
rect 12437 14977 12449 14980
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 9582 14900 9588 14952
rect 9640 14940 9646 14952
rect 12820 14940 12848 15048
rect 12894 14968 12900 15020
rect 12952 15008 12958 15020
rect 13078 15008 13084 15020
rect 12952 14980 12997 15008
rect 13039 14980 13084 15008
rect 12952 14968 12958 14980
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 13740 15017 13768 15048
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 15008 13783 15011
rect 16040 15008 16068 15116
rect 18690 15104 18696 15116
rect 18748 15104 18754 15156
rect 19150 15104 19156 15156
rect 19208 15144 19214 15156
rect 20073 15147 20131 15153
rect 20073 15144 20085 15147
rect 19208 15116 20085 15144
rect 19208 15104 19214 15116
rect 20073 15113 20085 15116
rect 20119 15113 20131 15147
rect 20073 15107 20131 15113
rect 18046 15076 18052 15088
rect 18007 15048 18052 15076
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 18969 15079 19027 15085
rect 18969 15045 18981 15079
rect 19015 15076 19027 15079
rect 19242 15076 19248 15088
rect 19015 15048 19248 15076
rect 19015 15045 19027 15048
rect 18969 15039 19027 15045
rect 19242 15036 19248 15048
rect 19300 15076 19306 15088
rect 19300 15048 23152 15076
rect 19300 15036 19306 15048
rect 13771 14980 16068 15008
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 16114 14968 16120 15020
rect 16172 15008 16178 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16172 14980 16865 15008
rect 16172 14968 16178 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 17865 15011 17923 15017
rect 17865 14977 17877 15011
rect 17911 14977 17923 15011
rect 17865 14971 17923 14977
rect 9640 14912 12848 14940
rect 17880 14940 17908 14971
rect 18782 14968 18788 15020
rect 18840 15008 18846 15020
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 18840 14980 18889 15008
rect 18840 14968 18846 14980
rect 18877 14977 18889 14980
rect 18923 14977 18935 15011
rect 18877 14971 18935 14977
rect 19061 15011 19119 15017
rect 19061 14977 19073 15011
rect 19107 15008 19119 15011
rect 19794 15008 19800 15020
rect 19107 14980 19800 15008
rect 19107 14977 19119 14980
rect 19061 14971 19119 14977
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 19904 15017 19932 15048
rect 19889 15011 19947 15017
rect 19889 14977 19901 15011
rect 19935 14977 19947 15011
rect 19889 14971 19947 14977
rect 20165 15011 20223 15017
rect 20165 14977 20177 15011
rect 20211 14977 20223 15011
rect 20165 14971 20223 14977
rect 19426 14940 19432 14952
rect 17880 14912 19432 14940
rect 9640 14900 9646 14912
rect 19426 14900 19432 14912
rect 19484 14940 19490 14952
rect 20180 14940 20208 14971
rect 23124 14949 23152 15048
rect 19484 14912 20208 14940
rect 22833 14943 22891 14949
rect 19484 14900 19490 14912
rect 22833 14909 22845 14943
rect 22879 14909 22891 14943
rect 22833 14903 22891 14909
rect 23109 14943 23167 14949
rect 23109 14909 23121 14943
rect 23155 14940 23167 14943
rect 23290 14940 23296 14952
rect 23155 14912 23296 14940
rect 23155 14909 23167 14912
rect 23109 14903 23167 14909
rect 9122 14872 9128 14884
rect 8864 14844 9128 14872
rect 9122 14832 9128 14844
rect 9180 14872 9186 14884
rect 9180 14844 18552 14872
rect 9180 14832 9186 14844
rect 8938 14804 8944 14816
rect 8899 14776 8944 14804
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 12253 14807 12311 14813
rect 12253 14804 12265 14807
rect 11848 14776 12265 14804
rect 11848 14764 11854 14776
rect 12253 14773 12265 14776
rect 12299 14773 12311 14807
rect 12253 14767 12311 14773
rect 12989 14807 13047 14813
rect 12989 14773 13001 14807
rect 13035 14804 13047 14807
rect 13262 14804 13268 14816
rect 13035 14776 13268 14804
rect 13035 14773 13047 14776
rect 12989 14767 13047 14773
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 13538 14804 13544 14816
rect 13499 14776 13544 14804
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 16669 14807 16727 14813
rect 16669 14804 16681 14807
rect 15804 14776 16681 14804
rect 15804 14764 15810 14776
rect 16669 14773 16681 14776
rect 16715 14773 16727 14807
rect 16669 14767 16727 14773
rect 18233 14807 18291 14813
rect 18233 14773 18245 14807
rect 18279 14804 18291 14807
rect 18414 14804 18420 14816
rect 18279 14776 18420 14804
rect 18279 14773 18291 14776
rect 18233 14767 18291 14773
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 18524 14804 18552 14844
rect 18598 14832 18604 14884
rect 18656 14872 18662 14884
rect 18693 14875 18751 14881
rect 18693 14872 18705 14875
rect 18656 14844 18705 14872
rect 18656 14832 18662 14844
rect 18693 14841 18705 14844
rect 18739 14841 18751 14875
rect 22848 14872 22876 14903
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 23382 14872 23388 14884
rect 22848 14844 23388 14872
rect 18693 14835 18751 14841
rect 23382 14832 23388 14844
rect 23440 14832 23446 14884
rect 19245 14807 19303 14813
rect 19245 14804 19257 14807
rect 18524 14776 19257 14804
rect 19245 14773 19257 14776
rect 19291 14804 19303 14807
rect 19334 14804 19340 14816
rect 19291 14776 19340 14804
rect 19291 14773 19303 14776
rect 19245 14767 19303 14773
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 19705 14807 19763 14813
rect 19705 14773 19717 14807
rect 19751 14804 19763 14807
rect 20530 14804 20536 14816
rect 19751 14776 20536 14804
rect 19751 14773 19763 14776
rect 19705 14767 19763 14773
rect 20530 14764 20536 14776
rect 20588 14764 20594 14816
rect 1104 14714 44896 14736
rect 1104 14662 6424 14714
rect 6476 14662 6488 14714
rect 6540 14662 6552 14714
rect 6604 14662 6616 14714
rect 6668 14662 6680 14714
rect 6732 14662 17372 14714
rect 17424 14662 17436 14714
rect 17488 14662 17500 14714
rect 17552 14662 17564 14714
rect 17616 14662 17628 14714
rect 17680 14662 28320 14714
rect 28372 14662 28384 14714
rect 28436 14662 28448 14714
rect 28500 14662 28512 14714
rect 28564 14662 28576 14714
rect 28628 14662 39268 14714
rect 39320 14662 39332 14714
rect 39384 14662 39396 14714
rect 39448 14662 39460 14714
rect 39512 14662 39524 14714
rect 39576 14662 44896 14714
rect 1104 14640 44896 14662
rect 8386 14560 8392 14612
rect 8444 14600 8450 14612
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 8444 14572 9137 14600
rect 8444 14560 8450 14572
rect 9125 14569 9137 14572
rect 9171 14569 9183 14603
rect 9125 14563 9183 14569
rect 19518 14560 19524 14612
rect 19576 14600 19582 14612
rect 20533 14603 20591 14609
rect 20533 14600 20545 14603
rect 19576 14572 20545 14600
rect 19576 14560 19582 14572
rect 20533 14569 20545 14572
rect 20579 14569 20591 14603
rect 23845 14603 23903 14609
rect 23845 14600 23857 14603
rect 20533 14563 20591 14569
rect 20640 14572 23857 14600
rect 9214 14492 9220 14544
rect 9272 14532 9278 14544
rect 9309 14535 9367 14541
rect 9309 14532 9321 14535
rect 9272 14504 9321 14532
rect 9272 14492 9278 14504
rect 9309 14501 9321 14504
rect 9355 14532 9367 14535
rect 9355 14504 12020 14532
rect 9355 14501 9367 14504
rect 9309 14495 9367 14501
rect 9490 14464 9496 14476
rect 7576 14436 9496 14464
rect 7576 14405 7604 14436
rect 9490 14424 9496 14436
rect 9548 14424 9554 14476
rect 11992 14464 12020 14504
rect 19150 14492 19156 14544
rect 19208 14532 19214 14544
rect 19208 14504 19748 14532
rect 19208 14492 19214 14504
rect 12526 14464 12532 14476
rect 11992 14436 12532 14464
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 8205 14399 8263 14405
rect 8205 14365 8217 14399
rect 8251 14396 8263 14399
rect 9766 14396 9772 14408
rect 8251 14368 9772 14396
rect 8251 14365 8263 14368
rect 8205 14359 8263 14365
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 11992 14405 12020 14436
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 12710 14424 12716 14476
rect 12768 14464 12774 14476
rect 19720 14473 19748 14504
rect 19705 14467 19763 14473
rect 12768 14436 13216 14464
rect 12768 14424 12774 14436
rect 11977 14399 12035 14405
rect 11977 14365 11989 14399
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14396 12219 14399
rect 12894 14396 12900 14408
rect 12207 14368 12900 14396
rect 12207 14365 12219 14368
rect 12161 14359 12219 14365
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 13078 14396 13084 14408
rect 13039 14368 13084 14396
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 13188 14405 13216 14436
rect 19705 14433 19717 14467
rect 19751 14433 19763 14467
rect 19705 14427 19763 14433
rect 19794 14424 19800 14476
rect 19852 14464 19858 14476
rect 20640 14464 20668 14572
rect 23845 14569 23857 14572
rect 23891 14600 23903 14603
rect 23934 14600 23940 14612
rect 23891 14572 23940 14600
rect 23891 14569 23903 14572
rect 23845 14563 23903 14569
rect 23934 14560 23940 14572
rect 23992 14560 23998 14612
rect 21729 14535 21787 14541
rect 21729 14501 21741 14535
rect 21775 14532 21787 14535
rect 21775 14504 22094 14532
rect 21775 14501 21787 14504
rect 21729 14495 21787 14501
rect 19852 14436 20668 14464
rect 19852 14424 19858 14436
rect 13173 14399 13231 14405
rect 13173 14365 13185 14399
rect 13219 14365 13231 14399
rect 13173 14359 13231 14365
rect 13262 14356 13268 14408
rect 13320 14396 13326 14408
rect 13449 14399 13507 14405
rect 13320 14368 13365 14396
rect 13320 14356 13326 14368
rect 13449 14365 13461 14399
rect 13495 14396 13507 14399
rect 13538 14396 13544 14408
rect 13495 14368 13544 14396
rect 13495 14365 13507 14368
rect 13449 14359 13507 14365
rect 8754 14288 8760 14340
rect 8812 14328 8818 14340
rect 8941 14331 8999 14337
rect 8941 14328 8953 14331
rect 8812 14300 8953 14328
rect 8812 14288 8818 14300
rect 8941 14297 8953 14300
rect 8987 14297 8999 14331
rect 8941 14291 8999 14297
rect 9122 14288 9128 14340
rect 9180 14337 9186 14340
rect 9180 14331 9199 14337
rect 9187 14297 9199 14331
rect 9180 14291 9199 14297
rect 9180 14288 9186 14291
rect 12618 14288 12624 14340
rect 12676 14328 12682 14340
rect 13464 14328 13492 14359
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 15470 14396 15476 14408
rect 15431 14368 15476 14396
rect 15470 14356 15476 14368
rect 15528 14396 15534 14408
rect 16666 14396 16672 14408
rect 15528 14368 16672 14396
rect 15528 14356 15534 14368
rect 16666 14356 16672 14368
rect 16724 14396 16730 14408
rect 17313 14399 17371 14405
rect 17313 14396 17325 14399
rect 16724 14368 17325 14396
rect 16724 14356 16730 14368
rect 17313 14365 17325 14368
rect 17359 14365 17371 14399
rect 17313 14359 17371 14365
rect 19242 14356 19248 14408
rect 19300 14396 19306 14408
rect 19521 14399 19579 14405
rect 19521 14396 19533 14399
rect 19300 14368 19533 14396
rect 19300 14356 19306 14368
rect 19521 14365 19533 14368
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 19610 14356 19616 14408
rect 19668 14396 19674 14408
rect 19668 14368 19713 14396
rect 19668 14356 19674 14368
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 21913 14399 21971 14405
rect 21913 14396 21925 14399
rect 20220 14368 21925 14396
rect 20220 14356 20226 14368
rect 21913 14365 21925 14368
rect 21959 14365 21971 14399
rect 21913 14359 21971 14365
rect 15562 14328 15568 14340
rect 12676 14300 15568 14328
rect 12676 14288 12682 14300
rect 15562 14288 15568 14300
rect 15620 14288 15626 14340
rect 15746 14337 15752 14340
rect 15740 14328 15752 14337
rect 15707 14300 15752 14328
rect 15740 14291 15752 14300
rect 15746 14288 15752 14291
rect 15804 14288 15810 14340
rect 17586 14337 17592 14340
rect 17580 14291 17592 14337
rect 17644 14328 17650 14340
rect 17644 14300 17680 14328
rect 17586 14288 17592 14291
rect 17644 14288 17650 14300
rect 19794 14288 19800 14340
rect 19852 14328 19858 14340
rect 20349 14331 20407 14337
rect 20349 14328 20361 14331
rect 19852 14300 20361 14328
rect 19852 14288 19858 14300
rect 20349 14297 20361 14300
rect 20395 14297 20407 14331
rect 20349 14291 20407 14297
rect 20530 14288 20536 14340
rect 20588 14337 20594 14340
rect 20588 14331 20607 14337
rect 20595 14297 20607 14331
rect 22066 14328 22094 14504
rect 22465 14399 22523 14405
rect 22465 14365 22477 14399
rect 22511 14396 22523 14399
rect 24670 14396 24676 14408
rect 22511 14368 24676 14396
rect 22511 14365 22523 14368
rect 22465 14359 22523 14365
rect 24670 14356 24676 14368
rect 24728 14356 24734 14408
rect 42978 14396 42984 14408
rect 42939 14368 42984 14396
rect 42978 14356 42984 14368
rect 43036 14356 43042 14408
rect 43901 14399 43959 14405
rect 43901 14365 43913 14399
rect 43947 14365 43959 14399
rect 43901 14359 43959 14365
rect 22710 14331 22768 14337
rect 22710 14328 22722 14331
rect 22066 14300 22722 14328
rect 20588 14291 20607 14297
rect 22710 14297 22722 14300
rect 22756 14297 22768 14331
rect 43916 14328 43944 14359
rect 22710 14291 22768 14297
rect 42812 14300 43944 14328
rect 20588 14288 20594 14291
rect 7374 14260 7380 14272
rect 7335 14232 7380 14260
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 8018 14260 8024 14272
rect 7979 14232 8024 14260
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 8570 14220 8576 14272
rect 8628 14260 8634 14272
rect 9140 14260 9168 14288
rect 12342 14260 12348 14272
rect 8628 14232 9168 14260
rect 12303 14232 12348 14260
rect 8628 14220 8634 14232
rect 12342 14220 12348 14232
rect 12400 14220 12406 14272
rect 12802 14260 12808 14272
rect 12763 14232 12808 14260
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 16850 14260 16856 14272
rect 16811 14232 16856 14260
rect 16850 14220 16856 14232
rect 16908 14260 16914 14272
rect 18598 14260 18604 14272
rect 16908 14232 18604 14260
rect 16908 14220 16914 14232
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 18693 14263 18751 14269
rect 18693 14229 18705 14263
rect 18739 14260 18751 14263
rect 18782 14260 18788 14272
rect 18739 14232 18788 14260
rect 18739 14229 18751 14232
rect 18693 14223 18751 14229
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 19337 14263 19395 14269
rect 19337 14229 19349 14263
rect 19383 14260 19395 14263
rect 19978 14260 19984 14272
rect 19383 14232 19984 14260
rect 19383 14229 19395 14232
rect 19337 14223 19395 14229
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 20717 14263 20775 14269
rect 20717 14229 20729 14263
rect 20763 14260 20775 14263
rect 21266 14260 21272 14272
rect 20763 14232 21272 14260
rect 20763 14229 20775 14232
rect 20717 14223 20775 14229
rect 21266 14220 21272 14232
rect 21324 14220 21330 14272
rect 21358 14220 21364 14272
rect 21416 14260 21422 14272
rect 23842 14260 23848 14272
rect 21416 14232 23848 14260
rect 21416 14220 21422 14232
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 42812 14269 42840 14300
rect 42797 14263 42855 14269
rect 42797 14229 42809 14263
rect 42843 14229 42855 14263
rect 44082 14260 44088 14272
rect 44043 14232 44088 14260
rect 42797 14223 42855 14229
rect 44082 14220 44088 14232
rect 44140 14220 44146 14272
rect 1104 14170 45056 14192
rect 1104 14118 11898 14170
rect 11950 14118 11962 14170
rect 12014 14118 12026 14170
rect 12078 14118 12090 14170
rect 12142 14118 12154 14170
rect 12206 14118 22846 14170
rect 22898 14118 22910 14170
rect 22962 14118 22974 14170
rect 23026 14118 23038 14170
rect 23090 14118 23102 14170
rect 23154 14118 33794 14170
rect 33846 14118 33858 14170
rect 33910 14118 33922 14170
rect 33974 14118 33986 14170
rect 34038 14118 34050 14170
rect 34102 14118 44742 14170
rect 44794 14118 44806 14170
rect 44858 14118 44870 14170
rect 44922 14118 44934 14170
rect 44986 14118 44998 14170
rect 45050 14118 45056 14170
rect 1104 14096 45056 14118
rect 3142 14056 3148 14068
rect 3103 14028 3148 14056
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 8386 14016 8392 14068
rect 8444 14056 8450 14068
rect 12250 14056 12256 14068
rect 8444 14028 9720 14056
rect 12211 14028 12256 14056
rect 8444 14016 8450 14028
rect 4430 13988 4436 14000
rect 3988 13960 4436 13988
rect 3326 13920 3332 13932
rect 3287 13892 3332 13920
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 3988 13929 4016 13960
rect 4430 13948 4436 13960
rect 4488 13948 4494 14000
rect 7374 13948 7380 14000
rect 7432 13988 7438 14000
rect 7622 13991 7680 13997
rect 7622 13988 7634 13991
rect 7432 13960 7634 13988
rect 7432 13948 7438 13960
rect 7622 13957 7634 13960
rect 7668 13957 7680 13991
rect 9582 13988 9588 14000
rect 9543 13960 9588 13988
rect 7622 13951 7680 13957
rect 9582 13948 9588 13960
rect 9640 13948 9646 14000
rect 9692 13988 9720 14028
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 12710 14056 12716 14068
rect 12406 14028 12716 14056
rect 10413 13991 10471 13997
rect 10413 13988 10425 13991
rect 9692 13960 10425 13988
rect 10413 13957 10425 13960
rect 10459 13957 10471 13991
rect 10413 13951 10471 13957
rect 11885 13991 11943 13997
rect 11885 13957 11897 13991
rect 11931 13957 11943 13991
rect 11885 13951 11943 13957
rect 12101 13991 12159 13997
rect 12101 13957 12113 13991
rect 12147 13988 12159 13991
rect 12406 13988 12434 14028
rect 12710 14016 12716 14028
rect 12768 14056 12774 14068
rect 12986 14056 12992 14068
rect 12768 14028 12992 14056
rect 12768 14016 12774 14028
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 14645 14059 14703 14065
rect 14645 14056 14657 14059
rect 13136 14028 14657 14056
rect 13136 14016 13142 14028
rect 14645 14025 14657 14028
rect 14691 14056 14703 14059
rect 15010 14056 15016 14068
rect 14691 14028 15016 14056
rect 14691 14025 14703 14028
rect 14645 14019 14703 14025
rect 15010 14016 15016 14028
rect 15068 14016 15074 14068
rect 16114 14056 16120 14068
rect 16075 14028 16120 14056
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 17586 14056 17592 14068
rect 17547 14028 17592 14056
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 19794 14056 19800 14068
rect 18248 14028 19800 14056
rect 15470 13988 15476 14000
rect 12147 13960 12434 13988
rect 12728 13960 15476 13988
rect 12147 13957 12159 13960
rect 12101 13951 12159 13957
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 4240 13923 4298 13929
rect 4240 13889 4252 13923
rect 4286 13920 4298 13923
rect 4286 13892 8432 13920
rect 4286 13889 4298 13892
rect 4240 13883 4298 13889
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7377 13855 7435 13861
rect 7377 13852 7389 13855
rect 7156 13824 7389 13852
rect 7156 13812 7162 13824
rect 7377 13821 7389 13824
rect 7423 13821 7435 13855
rect 8404 13852 8432 13892
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 8996 13892 10241 13920
rect 8996 13880 9002 13892
rect 10229 13889 10241 13892
rect 10275 13889 10287 13923
rect 11900 13920 11928 13951
rect 12618 13920 12624 13932
rect 11900 13892 12624 13920
rect 10229 13883 10287 13889
rect 12618 13880 12624 13892
rect 12676 13880 12682 13932
rect 12728 13929 12756 13960
rect 15470 13948 15476 13960
rect 15528 13948 15534 14000
rect 15562 13948 15568 14000
rect 15620 13988 15626 14000
rect 18248 13997 18276 14028
rect 19794 14016 19800 14028
rect 19852 14016 19858 14068
rect 20162 14056 20168 14068
rect 20123 14028 20168 14056
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 21085 14059 21143 14065
rect 21085 14025 21097 14059
rect 21131 14056 21143 14059
rect 23382 14056 23388 14068
rect 21131 14028 22094 14056
rect 23343 14028 23388 14056
rect 21131 14025 21143 14028
rect 21085 14019 21143 14025
rect 18506 13997 18512 14000
rect 18233 13991 18291 13997
rect 18233 13988 18245 13991
rect 15620 13960 18245 13988
rect 15620 13948 15626 13960
rect 12713 13923 12771 13929
rect 12713 13889 12725 13923
rect 12759 13889 12771 13923
rect 12713 13883 12771 13889
rect 12802 13880 12808 13932
rect 12860 13920 12866 13932
rect 15948 13929 15976 13960
rect 18233 13957 18245 13960
rect 18279 13957 18291 13991
rect 18233 13951 18291 13957
rect 18449 13991 18512 13997
rect 18449 13957 18461 13991
rect 18495 13957 18512 13991
rect 18449 13951 18512 13957
rect 18506 13948 18512 13951
rect 18564 13948 18570 14000
rect 18690 13948 18696 14000
rect 18748 13988 18754 14000
rect 19981 13991 20039 13997
rect 19981 13988 19993 13991
rect 18748 13960 19993 13988
rect 18748 13948 18754 13960
rect 19981 13957 19993 13960
rect 20027 13988 20039 13991
rect 21358 13988 21364 14000
rect 20027 13960 21364 13988
rect 20027 13957 20039 13960
rect 19981 13951 20039 13957
rect 21358 13948 21364 13960
rect 21416 13948 21422 14000
rect 22066 13988 22094 14028
rect 23382 14016 23388 14028
rect 23440 14056 23446 14068
rect 33321 14059 33379 14065
rect 23440 14028 24900 14056
rect 23440 14016 23446 14028
rect 24872 13997 24900 14028
rect 33321 14025 33333 14059
rect 33367 14056 33379 14059
rect 34882 14056 34888 14068
rect 33367 14028 34888 14056
rect 33367 14025 33379 14028
rect 33321 14019 33379 14025
rect 34882 14016 34888 14028
rect 34940 14016 34946 14068
rect 22250 13991 22308 13997
rect 22250 13988 22262 13991
rect 22066 13960 22262 13988
rect 22250 13957 22262 13960
rect 22296 13957 22308 13991
rect 24857 13991 24915 13997
rect 22250 13951 22308 13957
rect 23400 13960 24164 13988
rect 23400 13932 23428 13960
rect 12969 13923 13027 13929
rect 12969 13920 12981 13923
rect 12860 13892 12981 13920
rect 12860 13880 12866 13892
rect 12969 13889 12981 13892
rect 13015 13889 13027 13923
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 12969 13883 13027 13889
rect 14108 13892 14565 13920
rect 9674 13852 9680 13864
rect 8404 13824 9680 13852
rect 7377 13815 7435 13821
rect 9674 13812 9680 13824
rect 9732 13812 9738 13864
rect 11992 13824 12434 13852
rect 9214 13784 9220 13796
rect 4908 13756 6914 13784
rect 9175 13756 9220 13784
rect 3050 13676 3056 13728
rect 3108 13716 3114 13728
rect 4908 13716 4936 13756
rect 5350 13716 5356 13728
rect 3108 13688 4936 13716
rect 5311 13688 5356 13716
rect 3108 13676 3114 13688
rect 5350 13676 5356 13688
rect 5408 13676 5414 13728
rect 6886 13716 6914 13756
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 10597 13787 10655 13793
rect 10597 13784 10609 13787
rect 9600 13756 10609 13784
rect 8662 13716 8668 13728
rect 6886 13688 8668 13716
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 9600 13725 9628 13756
rect 10597 13753 10609 13756
rect 10643 13753 10655 13787
rect 10597 13747 10655 13753
rect 11146 13744 11152 13796
rect 11204 13784 11210 13796
rect 11992 13784 12020 13824
rect 11204 13756 12020 13784
rect 12406 13784 12434 13824
rect 14108 13793 14136 13892
rect 14553 13889 14565 13892
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13889 15991 13923
rect 15933 13883 15991 13889
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13920 16727 13923
rect 16850 13920 16856 13932
rect 16715 13892 16856 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 17773 13923 17831 13929
rect 17773 13889 17785 13923
rect 17819 13920 17831 13923
rect 18598 13920 18604 13932
rect 17819 13892 18604 13920
rect 17819 13889 17831 13892
rect 17773 13883 17831 13889
rect 18598 13880 18604 13892
rect 18656 13880 18662 13932
rect 19334 13880 19340 13932
rect 19392 13920 19398 13932
rect 19613 13923 19671 13929
rect 19613 13920 19625 13923
rect 19392 13892 19625 13920
rect 19392 13880 19398 13892
rect 19613 13889 19625 13892
rect 19659 13889 19671 13923
rect 21266 13920 21272 13932
rect 21227 13892 21272 13920
rect 19613 13883 19671 13889
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 23382 13880 23388 13932
rect 23440 13880 23446 13932
rect 24029 13923 24087 13929
rect 24029 13920 24041 13923
rect 23492 13892 24041 13920
rect 15749 13855 15807 13861
rect 15749 13821 15761 13855
rect 15795 13852 15807 13855
rect 16298 13852 16304 13864
rect 15795 13824 16304 13852
rect 15795 13821 15807 13824
rect 15749 13815 15807 13821
rect 16298 13812 16304 13824
rect 16356 13852 16362 13864
rect 16761 13855 16819 13861
rect 16761 13852 16773 13855
rect 16356 13824 16773 13852
rect 16356 13812 16362 13824
rect 16761 13821 16773 13824
rect 16807 13821 16819 13855
rect 16761 13815 16819 13821
rect 20622 13812 20628 13864
rect 20680 13852 20686 13864
rect 22005 13855 22063 13861
rect 22005 13852 22017 13855
rect 20680 13824 22017 13852
rect 20680 13812 20686 13824
rect 22005 13821 22017 13824
rect 22051 13821 22063 13855
rect 22005 13815 22063 13821
rect 23198 13812 23204 13864
rect 23256 13852 23262 13864
rect 23492 13852 23520 13892
rect 24029 13889 24041 13892
rect 24075 13889 24087 13923
rect 24029 13883 24087 13889
rect 23934 13852 23940 13864
rect 23256 13824 23520 13852
rect 23895 13824 23940 13852
rect 23256 13812 23262 13824
rect 23934 13812 23940 13824
rect 23992 13812 23998 13864
rect 24136 13852 24164 13960
rect 24857 13957 24869 13991
rect 24903 13957 24915 13991
rect 33686 13988 33692 14000
rect 33599 13960 33692 13988
rect 24857 13951 24915 13957
rect 33686 13948 33692 13960
rect 33744 13988 33750 14000
rect 42978 13988 42984 14000
rect 33744 13960 42984 13988
rect 33744 13948 33750 13960
rect 42978 13948 42984 13960
rect 43036 13948 43042 14000
rect 24210 13880 24216 13932
rect 24268 13920 24274 13932
rect 25041 13923 25099 13929
rect 25041 13920 25053 13923
rect 24268 13892 25053 13920
rect 24268 13880 24274 13892
rect 25041 13889 25053 13892
rect 25087 13889 25099 13923
rect 25041 13883 25099 13889
rect 33226 13880 33232 13932
rect 33284 13920 33290 13932
rect 33284 13892 33916 13920
rect 33284 13880 33290 13892
rect 33888 13861 33916 13892
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 24136 13824 25237 13852
rect 25225 13821 25237 13824
rect 25271 13821 25283 13855
rect 33781 13855 33839 13861
rect 33781 13852 33793 13855
rect 25225 13815 25283 13821
rect 28966 13824 33364 13852
rect 14093 13787 14151 13793
rect 12406 13756 12480 13784
rect 11204 13744 11210 13756
rect 9585 13719 9643 13725
rect 8812 13688 8857 13716
rect 8812 13676 8818 13688
rect 9585 13685 9597 13719
rect 9631 13685 9643 13719
rect 9766 13716 9772 13728
rect 9727 13688 9772 13716
rect 9585 13679 9643 13685
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 12069 13719 12127 13725
rect 12069 13685 12081 13719
rect 12115 13716 12127 13719
rect 12342 13716 12348 13728
rect 12115 13688 12348 13716
rect 12115 13685 12127 13688
rect 12069 13679 12127 13685
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 12452 13716 12480 13756
rect 14093 13753 14105 13787
rect 14139 13753 14151 13787
rect 14093 13747 14151 13753
rect 16390 13744 16396 13796
rect 16448 13784 16454 13796
rect 16448 13756 20116 13784
rect 16448 13744 16454 13756
rect 16850 13716 16856 13728
rect 12452 13688 16856 13716
rect 16850 13676 16856 13688
rect 16908 13676 16914 13728
rect 18414 13716 18420 13728
rect 18375 13688 18420 13716
rect 18414 13676 18420 13688
rect 18472 13676 18478 13728
rect 18598 13716 18604 13728
rect 18559 13688 18604 13716
rect 18598 13676 18604 13688
rect 18656 13676 18662 13728
rect 19978 13716 19984 13728
rect 19939 13688 19984 13716
rect 19978 13676 19984 13688
rect 20036 13676 20042 13728
rect 20088 13716 20116 13756
rect 23308 13756 25360 13784
rect 23308 13716 23336 13756
rect 20088 13688 23336 13716
rect 23474 13676 23480 13728
rect 23532 13716 23538 13728
rect 24397 13719 24455 13725
rect 24397 13716 24409 13719
rect 23532 13688 24409 13716
rect 23532 13676 23538 13688
rect 24397 13685 24409 13688
rect 24443 13685 24455 13719
rect 25332 13716 25360 13756
rect 25406 13744 25412 13796
rect 25464 13784 25470 13796
rect 28966 13784 28994 13824
rect 25464 13756 28994 13784
rect 25464 13744 25470 13756
rect 33226 13716 33232 13728
rect 25332 13688 33232 13716
rect 24397 13679 24455 13685
rect 33226 13676 33232 13688
rect 33284 13676 33290 13728
rect 33336 13716 33364 13824
rect 33704 13824 33793 13852
rect 33704 13796 33732 13824
rect 33781 13821 33793 13824
rect 33827 13821 33839 13855
rect 33781 13815 33839 13821
rect 33873 13855 33931 13861
rect 33873 13821 33885 13855
rect 33919 13852 33931 13855
rect 34514 13852 34520 13864
rect 33919 13824 34520 13852
rect 33919 13821 33931 13824
rect 33873 13815 33931 13821
rect 34514 13812 34520 13824
rect 34572 13812 34578 13864
rect 33686 13744 33692 13796
rect 33744 13744 33750 13796
rect 38930 13716 38936 13728
rect 33336 13688 38936 13716
rect 38930 13676 38936 13688
rect 38988 13676 38994 13728
rect 1104 13626 44896 13648
rect 1104 13574 6424 13626
rect 6476 13574 6488 13626
rect 6540 13574 6552 13626
rect 6604 13574 6616 13626
rect 6668 13574 6680 13626
rect 6732 13574 17372 13626
rect 17424 13574 17436 13626
rect 17488 13574 17500 13626
rect 17552 13574 17564 13626
rect 17616 13574 17628 13626
rect 17680 13574 28320 13626
rect 28372 13574 28384 13626
rect 28436 13574 28448 13626
rect 28500 13574 28512 13626
rect 28564 13574 28576 13626
rect 28628 13574 39268 13626
rect 39320 13574 39332 13626
rect 39384 13574 39396 13626
rect 39448 13574 39460 13626
rect 39512 13574 39524 13626
rect 39576 13574 44896 13626
rect 1104 13552 44896 13574
rect 8386 13512 8392 13524
rect 8347 13484 8392 13512
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 9030 13472 9036 13524
rect 9088 13512 9094 13524
rect 9309 13515 9367 13521
rect 9309 13512 9321 13515
rect 9088 13484 9321 13512
rect 9088 13472 9094 13484
rect 9309 13481 9321 13484
rect 9355 13481 9367 13515
rect 9490 13512 9496 13524
rect 9451 13484 9496 13512
rect 9309 13475 9367 13481
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 9600 13484 39160 13512
rect 8938 13444 8944 13456
rect 8899 13416 8944 13444
rect 8938 13404 8944 13416
rect 8996 13404 9002 13456
rect 8662 13336 8668 13388
rect 8720 13376 8726 13388
rect 9600 13376 9628 13484
rect 12986 13404 12992 13456
rect 13044 13444 13050 13456
rect 14185 13447 14243 13453
rect 14185 13444 14197 13447
rect 13044 13416 14197 13444
rect 13044 13404 13050 13416
rect 14185 13413 14197 13416
rect 14231 13413 14243 13447
rect 14185 13407 14243 13413
rect 14829 13447 14887 13453
rect 14829 13413 14841 13447
rect 14875 13444 14887 13447
rect 16022 13444 16028 13456
rect 14875 13416 16028 13444
rect 14875 13413 14887 13416
rect 14829 13407 14887 13413
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 17957 13447 18015 13453
rect 17957 13444 17969 13447
rect 16132 13416 17969 13444
rect 8720 13348 9628 13376
rect 8720 13336 8726 13348
rect 14458 13336 14464 13388
rect 14516 13376 14522 13388
rect 16132 13376 16160 13416
rect 17957 13413 17969 13416
rect 18003 13413 18015 13447
rect 17957 13407 18015 13413
rect 18506 13404 18512 13456
rect 18564 13444 18570 13456
rect 18601 13447 18659 13453
rect 18601 13444 18613 13447
rect 18564 13416 18613 13444
rect 18564 13404 18570 13416
rect 18601 13413 18613 13416
rect 18647 13413 18659 13447
rect 18601 13407 18659 13413
rect 19245 13447 19303 13453
rect 19245 13413 19257 13447
rect 19291 13444 19303 13447
rect 19426 13444 19432 13456
rect 19291 13416 19432 13444
rect 19291 13413 19303 13416
rect 19245 13407 19303 13413
rect 19426 13404 19432 13416
rect 19484 13404 19490 13456
rect 20254 13404 20260 13456
rect 20312 13444 20318 13456
rect 20990 13444 20996 13456
rect 20312 13416 20996 13444
rect 20312 13404 20318 13416
rect 20990 13404 20996 13416
rect 21048 13444 21054 13456
rect 21048 13416 21588 13444
rect 21048 13404 21054 13416
rect 14516 13348 16160 13376
rect 17681 13379 17739 13385
rect 14516 13336 14522 13348
rect 17681 13345 17693 13379
rect 17727 13376 17739 13379
rect 18782 13376 18788 13388
rect 17727 13348 18788 13376
rect 17727 13345 17739 13348
rect 17681 13339 17739 13345
rect 18782 13336 18788 13348
rect 18840 13376 18846 13388
rect 18840 13348 19472 13376
rect 18840 13336 18846 13348
rect 4430 13268 4436 13320
rect 4488 13308 4494 13320
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 4488 13280 7021 13308
rect 4488 13268 4494 13280
rect 7009 13277 7021 13280
rect 7055 13308 7067 13311
rect 7098 13308 7104 13320
rect 7055 13280 7104 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 7098 13268 7104 13280
rect 7156 13308 7162 13320
rect 8846 13308 8852 13320
rect 7156 13280 8852 13308
rect 7156 13268 7162 13280
rect 8846 13268 8852 13280
rect 8904 13268 8910 13320
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13308 10563 13311
rect 11146 13308 11152 13320
rect 10551 13280 11152 13308
rect 10551 13277 10563 13280
rect 10505 13271 10563 13277
rect 11146 13268 11152 13280
rect 11204 13268 11210 13320
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 7276 13243 7334 13249
rect 7276 13209 7288 13243
rect 7322 13240 7334 13243
rect 8018 13240 8024 13252
rect 7322 13212 8024 13240
rect 7322 13209 7334 13212
rect 7276 13203 7334 13209
rect 8018 13200 8024 13212
rect 8076 13200 8082 13252
rect 9309 13243 9367 13249
rect 9309 13209 9321 13243
rect 9355 13240 9367 13243
rect 9582 13240 9588 13252
rect 9355 13212 9588 13240
rect 9355 13209 9367 13212
rect 9309 13203 9367 13209
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 10778 13200 10784 13252
rect 10836 13240 10842 13252
rect 11808 13240 11836 13271
rect 11882 13268 11888 13320
rect 11940 13308 11946 13320
rect 12049 13311 12107 13317
rect 12049 13308 12061 13311
rect 11940 13280 12061 13308
rect 11940 13268 11946 13280
rect 12049 13277 12061 13280
rect 12095 13277 12107 13311
rect 12049 13271 12107 13277
rect 12526 13268 12532 13320
rect 12584 13308 12590 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 12584 13280 14105 13308
rect 12584 13268 12590 13280
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 15010 13311 15068 13317
rect 15010 13277 15022 13311
rect 15056 13308 15068 13311
rect 15286 13308 15292 13320
rect 15056 13280 15292 13308
rect 15056 13277 15068 13280
rect 15010 13271 15068 13277
rect 14292 13240 14320 13271
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 15381 13311 15439 13317
rect 15381 13277 15393 13311
rect 15427 13277 15439 13311
rect 15381 13271 15439 13277
rect 15396 13240 15424 13271
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 15933 13311 15991 13317
rect 15933 13308 15945 13311
rect 15528 13280 15945 13308
rect 15528 13268 15534 13280
rect 15933 13277 15945 13280
rect 15979 13277 15991 13311
rect 16298 13308 16304 13320
rect 16259 13280 16304 13308
rect 15933 13271 15991 13277
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 17589 13311 17647 13317
rect 17589 13277 17601 13311
rect 17635 13308 17647 13311
rect 17862 13308 17868 13320
rect 17635 13280 17868 13308
rect 17635 13277 17647 13280
rect 17589 13271 17647 13277
rect 17862 13268 17868 13280
rect 17920 13268 17926 13320
rect 18509 13311 18567 13317
rect 18509 13277 18521 13311
rect 18555 13277 18567 13311
rect 18509 13271 18567 13277
rect 18693 13311 18751 13317
rect 18693 13277 18705 13311
rect 18739 13308 18751 13311
rect 19150 13308 19156 13320
rect 18739 13280 19156 13308
rect 18739 13277 18751 13280
rect 18693 13271 18751 13277
rect 16117 13243 16175 13249
rect 16117 13240 16129 13243
rect 10836 13212 11836 13240
rect 13188 13212 16129 13240
rect 10836 13200 10842 13212
rect 10594 13172 10600 13184
rect 10555 13144 10600 13172
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 11241 13175 11299 13181
rect 11241 13141 11253 13175
rect 11287 13172 11299 13175
rect 11514 13172 11520 13184
rect 11287 13144 11520 13172
rect 11287 13141 11299 13144
rect 11241 13135 11299 13141
rect 11514 13132 11520 13144
rect 11572 13132 11578 13184
rect 12894 13132 12900 13184
rect 12952 13172 12958 13184
rect 13188 13181 13216 13212
rect 16117 13209 16129 13212
rect 16163 13209 16175 13243
rect 16117 13203 16175 13209
rect 16206 13200 16212 13252
rect 16264 13240 16270 13252
rect 18414 13240 18420 13252
rect 16264 13212 18420 13240
rect 16264 13200 16270 13212
rect 18414 13200 18420 13212
rect 18472 13200 18478 13252
rect 18524 13240 18552 13271
rect 19150 13268 19156 13280
rect 19208 13268 19214 13320
rect 19444 13317 19472 13348
rect 20622 13336 20628 13388
rect 20680 13376 20686 13388
rect 21453 13379 21511 13385
rect 21453 13376 21465 13379
rect 20680 13348 21465 13376
rect 20680 13336 20686 13348
rect 21453 13345 21465 13348
rect 21499 13345 21511 13379
rect 21560 13376 21588 13416
rect 22738 13404 22744 13456
rect 22796 13444 22802 13456
rect 25406 13444 25412 13456
rect 22796 13416 25412 13444
rect 22796 13404 22802 13416
rect 25406 13404 25412 13416
rect 25464 13404 25470 13456
rect 22186 13376 22192 13388
rect 21560 13348 22192 13376
rect 21453 13339 21511 13345
rect 22186 13336 22192 13348
rect 22244 13336 22250 13388
rect 22278 13336 22284 13388
rect 22336 13376 22342 13388
rect 23201 13379 23259 13385
rect 23201 13376 23213 13379
rect 22336 13348 23213 13376
rect 22336 13336 22342 13348
rect 23201 13345 23213 13348
rect 23247 13376 23259 13379
rect 32582 13376 32588 13388
rect 23247 13348 23888 13376
rect 23247 13345 23259 13348
rect 23201 13339 23259 13345
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13308 21051 13311
rect 21358 13308 21364 13320
rect 21039 13280 21364 13308
rect 21039 13277 21051 13280
rect 20993 13271 21051 13277
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 23290 13268 23296 13320
rect 23348 13308 23354 13320
rect 23860 13317 23888 13348
rect 24504 13348 32588 13376
rect 23661 13311 23719 13317
rect 23661 13308 23673 13311
rect 23348 13280 23673 13308
rect 23348 13268 23354 13280
rect 23661 13277 23673 13280
rect 23707 13277 23719 13311
rect 23661 13271 23719 13277
rect 23845 13311 23903 13317
rect 23845 13277 23857 13311
rect 23891 13308 23903 13311
rect 24210 13308 24216 13320
rect 23891 13280 24216 13308
rect 23891 13277 23903 13280
rect 23845 13271 23903 13277
rect 24210 13268 24216 13280
rect 24268 13268 24274 13320
rect 19334 13240 19340 13252
rect 18524 13212 19340 13240
rect 19334 13200 19340 13212
rect 19392 13200 19398 13252
rect 21729 13243 21787 13249
rect 21729 13240 21741 13243
rect 20824 13212 21741 13240
rect 13173 13175 13231 13181
rect 13173 13172 13185 13175
rect 12952 13144 13185 13172
rect 12952 13132 12958 13144
rect 13173 13141 13185 13144
rect 13219 13141 13231 13175
rect 15010 13172 15016 13184
rect 14971 13144 15016 13172
rect 13173 13135 13231 13141
rect 15010 13132 15016 13144
rect 15068 13132 15074 13184
rect 16482 13172 16488 13184
rect 16443 13144 16488 13172
rect 16482 13132 16488 13144
rect 16540 13132 16546 13184
rect 20824 13181 20852 13212
rect 21729 13209 21741 13212
rect 21775 13209 21787 13243
rect 21729 13203 21787 13209
rect 22738 13200 22744 13252
rect 22796 13200 22802 13252
rect 24504 13240 24532 13348
rect 32582 13336 32588 13348
rect 32640 13376 32646 13388
rect 37274 13376 37280 13388
rect 32640 13348 32904 13376
rect 37235 13348 37280 13376
rect 32640 13336 32646 13348
rect 26326 13308 26332 13320
rect 26287 13280 26332 13308
rect 26326 13268 26332 13280
rect 26384 13268 26390 13320
rect 26786 13308 26792 13320
rect 26747 13280 26792 13308
rect 26786 13268 26792 13280
rect 26844 13268 26850 13320
rect 30282 13308 30288 13320
rect 30243 13280 30288 13308
rect 30282 13268 30288 13280
rect 30340 13268 30346 13320
rect 32306 13268 32312 13320
rect 32364 13308 32370 13320
rect 32769 13311 32827 13317
rect 32769 13308 32781 13311
rect 32364 13280 32781 13308
rect 32364 13268 32370 13280
rect 32769 13277 32781 13280
rect 32815 13277 32827 13311
rect 32876 13308 32904 13348
rect 37274 13336 37280 13348
rect 37332 13336 37338 13388
rect 37737 13379 37795 13385
rect 37737 13345 37749 13379
rect 37783 13376 37795 13379
rect 38930 13376 38936 13388
rect 37783 13348 38936 13376
rect 37783 13345 37795 13348
rect 37737 13339 37795 13345
rect 38930 13336 38936 13348
rect 38988 13336 38994 13388
rect 33318 13308 33324 13320
rect 32876 13280 33324 13308
rect 32769 13271 32827 13277
rect 33318 13268 33324 13280
rect 33376 13268 33382 13320
rect 37369 13311 37427 13317
rect 37369 13277 37381 13311
rect 37415 13308 37427 13311
rect 37642 13308 37648 13320
rect 37415 13280 37648 13308
rect 37415 13277 37427 13280
rect 37369 13271 37427 13277
rect 37642 13268 37648 13280
rect 37700 13268 37706 13320
rect 38286 13308 38292 13320
rect 38247 13280 38292 13308
rect 38286 13268 38292 13280
rect 38344 13268 38350 13320
rect 38378 13268 38384 13320
rect 38436 13308 38442 13320
rect 39132 13317 39160 13484
rect 40313 13447 40371 13453
rect 40313 13413 40325 13447
rect 40359 13444 40371 13447
rect 40954 13444 40960 13456
rect 40359 13416 40960 13444
rect 40359 13413 40371 13416
rect 40313 13407 40371 13413
rect 40954 13404 40960 13416
rect 41012 13404 41018 13456
rect 41049 13447 41107 13453
rect 41049 13413 41061 13447
rect 41095 13444 41107 13447
rect 42610 13444 42616 13456
rect 41095 13416 42616 13444
rect 41095 13413 41107 13416
rect 41049 13407 41107 13413
rect 42610 13404 42616 13416
rect 42668 13404 42674 13456
rect 39117 13311 39175 13317
rect 38436 13280 38529 13308
rect 38436 13268 38442 13280
rect 39117 13277 39129 13311
rect 39163 13277 39175 13311
rect 39117 13271 39175 13277
rect 39666 13268 39672 13320
rect 39724 13308 39730 13320
rect 40589 13311 40647 13317
rect 40589 13308 40601 13311
rect 39724 13280 40601 13308
rect 39724 13268 39730 13280
rect 40589 13277 40601 13280
rect 40635 13308 40647 13311
rect 41325 13311 41383 13317
rect 41325 13308 41337 13311
rect 40635 13280 41337 13308
rect 40635 13277 40647 13280
rect 40589 13271 40647 13277
rect 41325 13277 41337 13280
rect 41371 13277 41383 13311
rect 41325 13271 41383 13277
rect 23032 13212 24532 13240
rect 27065 13243 27123 13249
rect 20809 13175 20867 13181
rect 20809 13141 20821 13175
rect 20855 13141 20867 13175
rect 20809 13135 20867 13141
rect 22370 13132 22376 13184
rect 22428 13172 22434 13184
rect 22646 13172 22652 13184
rect 22428 13144 22652 13172
rect 22428 13132 22434 13144
rect 22646 13132 22652 13144
rect 22704 13172 22710 13184
rect 23032 13172 23060 13212
rect 27065 13209 27077 13243
rect 27111 13209 27123 13243
rect 27065 13203 27123 13209
rect 22704 13144 23060 13172
rect 22704 13132 22710 13144
rect 23290 13132 23296 13184
rect 23348 13172 23354 13184
rect 23753 13175 23811 13181
rect 23753 13172 23765 13175
rect 23348 13144 23765 13172
rect 23348 13132 23354 13144
rect 23753 13141 23765 13144
rect 23799 13141 23811 13175
rect 23753 13135 23811 13141
rect 26145 13175 26203 13181
rect 26145 13141 26157 13175
rect 26191 13172 26203 13175
rect 27080 13172 27108 13203
rect 27798 13200 27804 13252
rect 27856 13200 27862 13252
rect 33036 13243 33094 13249
rect 33036 13209 33048 13243
rect 33082 13240 33094 13243
rect 33226 13240 33232 13252
rect 33082 13212 33232 13240
rect 33082 13209 33094 13212
rect 33036 13203 33094 13209
rect 33226 13200 33232 13212
rect 33284 13200 33290 13252
rect 37660 13240 37688 13268
rect 38396 13240 38424 13268
rect 37660 13212 38424 13240
rect 38470 13200 38476 13252
rect 38528 13240 38534 13252
rect 40313 13243 40371 13249
rect 40313 13240 40325 13243
rect 38528 13212 40325 13240
rect 38528 13200 38534 13212
rect 40313 13209 40325 13212
rect 40359 13209 40371 13243
rect 40313 13203 40371 13209
rect 41049 13243 41107 13249
rect 41049 13209 41061 13243
rect 41095 13240 41107 13243
rect 41966 13240 41972 13252
rect 41095 13212 41972 13240
rect 41095 13209 41107 13212
rect 41049 13203 41107 13209
rect 41966 13200 41972 13212
rect 42024 13200 42030 13252
rect 26191 13144 27108 13172
rect 28537 13175 28595 13181
rect 26191 13141 26203 13144
rect 26145 13135 26203 13141
rect 28537 13141 28549 13175
rect 28583 13172 28595 13175
rect 28718 13172 28724 13184
rect 28583 13144 28724 13172
rect 28583 13141 28595 13144
rect 28537 13135 28595 13141
rect 28718 13132 28724 13144
rect 28776 13132 28782 13184
rect 30377 13175 30435 13181
rect 30377 13141 30389 13175
rect 30423 13172 30435 13175
rect 30466 13172 30472 13184
rect 30423 13144 30472 13172
rect 30423 13141 30435 13144
rect 30377 13135 30435 13141
rect 30466 13132 30472 13144
rect 30524 13132 30530 13184
rect 34149 13175 34207 13181
rect 34149 13141 34161 13175
rect 34195 13172 34207 13175
rect 35618 13172 35624 13184
rect 34195 13144 35624 13172
rect 34195 13141 34207 13144
rect 34149 13135 34207 13141
rect 35618 13132 35624 13144
rect 35676 13132 35682 13184
rect 38562 13172 38568 13184
rect 38523 13144 38568 13172
rect 38562 13132 38568 13144
rect 38620 13132 38626 13184
rect 39209 13175 39267 13181
rect 39209 13141 39221 13175
rect 39255 13172 39267 13175
rect 40218 13172 40224 13184
rect 39255 13144 40224 13172
rect 39255 13141 39267 13144
rect 39209 13135 39267 13141
rect 40218 13132 40224 13144
rect 40276 13132 40282 13184
rect 40494 13172 40500 13184
rect 40455 13144 40500 13172
rect 40494 13132 40500 13144
rect 40552 13172 40558 13184
rect 41233 13175 41291 13181
rect 41233 13172 41245 13175
rect 40552 13144 41245 13172
rect 40552 13132 40558 13144
rect 41233 13141 41245 13144
rect 41279 13141 41291 13175
rect 41233 13135 41291 13141
rect 1104 13082 45056 13104
rect 1104 13030 11898 13082
rect 11950 13030 11962 13082
rect 12014 13030 12026 13082
rect 12078 13030 12090 13082
rect 12142 13030 12154 13082
rect 12206 13030 22846 13082
rect 22898 13030 22910 13082
rect 22962 13030 22974 13082
rect 23026 13030 23038 13082
rect 23090 13030 23102 13082
rect 23154 13030 33794 13082
rect 33846 13030 33858 13082
rect 33910 13030 33922 13082
rect 33974 13030 33986 13082
rect 34038 13030 34050 13082
rect 34102 13030 44742 13082
rect 44794 13030 44806 13082
rect 44858 13030 44870 13082
rect 44922 13030 44934 13082
rect 44986 13030 44998 13082
rect 45050 13030 45056 13082
rect 1104 13008 45056 13030
rect 22278 12968 22284 12980
rect 3160 12940 22094 12968
rect 22239 12940 22284 12968
rect 3160 12841 3188 12940
rect 4700 12903 4758 12909
rect 4700 12869 4712 12903
rect 4746 12900 4758 12903
rect 5350 12900 5356 12912
rect 4746 12872 5356 12900
rect 4746 12869 4758 12872
rect 4700 12863 4758 12869
rect 5350 12860 5356 12872
rect 5408 12860 5414 12912
rect 8570 12860 8576 12912
rect 8628 12900 8634 12912
rect 8665 12903 8723 12909
rect 8665 12900 8677 12903
rect 8628 12872 8677 12900
rect 8628 12860 8634 12872
rect 8665 12869 8677 12872
rect 8711 12869 8723 12903
rect 9030 12900 9036 12912
rect 8991 12872 9036 12900
rect 8665 12863 8723 12869
rect 9030 12860 9036 12872
rect 9088 12860 9094 12912
rect 9784 12872 10640 12900
rect 3145 12835 3203 12841
rect 3145 12801 3157 12835
rect 3191 12801 3203 12835
rect 4430 12832 4436 12844
rect 4391 12804 4436 12832
rect 3145 12795 3203 12801
rect 4430 12792 4436 12804
rect 4488 12792 4494 12844
rect 8754 12792 8760 12844
rect 8812 12832 8818 12844
rect 8849 12835 8907 12841
rect 8849 12832 8861 12835
rect 8812 12804 8861 12832
rect 8812 12792 8818 12804
rect 8849 12801 8861 12804
rect 8895 12832 8907 12835
rect 9784 12832 9812 12872
rect 8895 12804 9812 12832
rect 9861 12835 9919 12841
rect 8895 12801 8907 12804
rect 8849 12795 8907 12801
rect 9861 12801 9873 12835
rect 9907 12832 9919 12835
rect 10502 12832 10508 12844
rect 9907 12804 10508 12832
rect 9907 12801 9919 12804
rect 9861 12795 9919 12801
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 9769 12767 9827 12773
rect 9769 12764 9781 12767
rect 8444 12736 9781 12764
rect 8444 12724 8450 12736
rect 9769 12733 9781 12736
rect 9815 12733 9827 12767
rect 10612 12764 10640 12872
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 13633 12903 13691 12909
rect 13633 12900 13645 12903
rect 12584 12872 13645 12900
rect 12584 12860 12590 12872
rect 13633 12869 13645 12872
rect 13679 12869 13691 12903
rect 13633 12863 13691 12869
rect 13817 12903 13875 12909
rect 13817 12869 13829 12903
rect 13863 12900 13875 12903
rect 13863 12872 14780 12900
rect 13863 12869 13875 12872
rect 13817 12863 13875 12869
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 11977 12835 12035 12841
rect 11977 12832 11989 12835
rect 10744 12804 11989 12832
rect 10744 12792 10750 12804
rect 11977 12801 11989 12804
rect 12023 12801 12035 12835
rect 12986 12832 12992 12844
rect 12947 12804 12992 12832
rect 11977 12795 12035 12801
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13449 12835 13507 12841
rect 13449 12801 13461 12835
rect 13495 12832 13507 12835
rect 13906 12832 13912 12844
rect 13495 12804 13912 12832
rect 13495 12801 13507 12804
rect 13449 12795 13507 12801
rect 13464 12764 13492 12795
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 14458 12832 14464 12844
rect 14419 12804 14464 12832
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 14642 12832 14648 12844
rect 14603 12804 14648 12832
rect 14642 12792 14648 12804
rect 14700 12792 14706 12844
rect 14752 12841 14780 12872
rect 15286 12860 15292 12912
rect 15344 12900 15350 12912
rect 15930 12900 15936 12912
rect 15344 12872 15936 12900
rect 15344 12860 15350 12872
rect 15488 12841 15516 12872
rect 15930 12860 15936 12872
rect 15988 12860 15994 12912
rect 17770 12860 17776 12912
rect 17828 12860 17834 12912
rect 22066 12900 22094 12940
rect 22278 12928 22284 12940
rect 22336 12928 22342 12980
rect 22370 12928 22376 12980
rect 22428 12968 22434 12980
rect 23290 12968 23296 12980
rect 22428 12940 22473 12968
rect 23251 12940 23296 12968
rect 22428 12928 22434 12940
rect 23290 12928 23296 12940
rect 23348 12928 23354 12980
rect 23842 12968 23848 12980
rect 23803 12940 23848 12968
rect 23842 12928 23848 12940
rect 23900 12928 23906 12980
rect 24026 12968 24032 12980
rect 23987 12940 24032 12968
rect 24026 12928 24032 12940
rect 24084 12928 24090 12980
rect 33505 12971 33563 12977
rect 24136 12940 31754 12968
rect 24136 12900 24164 12940
rect 18984 12872 21588 12900
rect 22066 12872 24164 12900
rect 14737 12835 14795 12841
rect 14737 12801 14749 12835
rect 14783 12801 14795 12835
rect 15197 12835 15255 12841
rect 15197 12832 15209 12835
rect 14737 12795 14795 12801
rect 14844 12804 15209 12832
rect 10612 12736 13492 12764
rect 9769 12727 9827 12733
rect 10229 12699 10287 12705
rect 10229 12665 10241 12699
rect 10275 12696 10287 12699
rect 14844 12696 14872 12804
rect 15197 12801 15209 12804
rect 15243 12801 15255 12835
rect 15381 12835 15439 12841
rect 15381 12832 15393 12835
rect 15197 12795 15255 12801
rect 15304 12804 15393 12832
rect 15304 12776 15332 12804
rect 15381 12801 15393 12804
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 15473 12835 15531 12841
rect 15473 12801 15485 12835
rect 15519 12801 15531 12835
rect 15473 12795 15531 12801
rect 15749 12835 15807 12841
rect 15749 12801 15761 12835
rect 15795 12832 15807 12835
rect 16206 12832 16212 12844
rect 15795 12804 16212 12832
rect 15795 12801 15807 12804
rect 15749 12795 15807 12801
rect 16206 12792 16212 12804
rect 16264 12792 16270 12844
rect 16666 12832 16672 12844
rect 16627 12804 16672 12832
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 17862 12792 17868 12844
rect 17920 12832 17926 12844
rect 18463 12835 18521 12841
rect 18463 12832 18475 12835
rect 17920 12804 18475 12832
rect 17920 12792 17926 12804
rect 18463 12801 18475 12804
rect 18509 12801 18521 12835
rect 18463 12795 18521 12801
rect 15286 12724 15292 12776
rect 15344 12724 15350 12776
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12764 15623 12767
rect 16298 12764 16304 12776
rect 15611 12736 16304 12764
rect 15611 12733 15623 12736
rect 15565 12727 15623 12733
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 17034 12764 17040 12776
rect 16995 12736 17040 12764
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 10275 12668 14872 12696
rect 10275 12665 10287 12668
rect 10229 12659 10287 12665
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 2961 12631 3019 12637
rect 2961 12628 2973 12631
rect 2832 12600 2973 12628
rect 2832 12588 2838 12600
rect 2961 12597 2973 12600
rect 3007 12597 3019 12631
rect 2961 12591 3019 12597
rect 5813 12631 5871 12637
rect 5813 12597 5825 12631
rect 5859 12628 5871 12631
rect 5994 12628 6000 12640
rect 5859 12600 6000 12628
rect 5859 12597 5871 12600
rect 5813 12591 5871 12597
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 10870 12628 10876 12640
rect 10831 12600 10876 12628
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 12069 12631 12127 12637
rect 12069 12597 12081 12631
rect 12115 12628 12127 12631
rect 12158 12628 12164 12640
rect 12115 12600 12164 12628
rect 12115 12597 12127 12600
rect 12069 12591 12127 12597
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 12805 12631 12863 12637
rect 12805 12597 12817 12631
rect 12851 12628 12863 12631
rect 13354 12628 13360 12640
rect 12851 12600 13360 12628
rect 12851 12597 12863 12600
rect 12805 12591 12863 12597
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 14461 12631 14519 12637
rect 14461 12597 14473 12631
rect 14507 12628 14519 12631
rect 15838 12628 15844 12640
rect 14507 12600 15844 12628
rect 14507 12597 14519 12600
rect 14461 12591 14519 12597
rect 15838 12588 15844 12600
rect 15896 12588 15902 12640
rect 15933 12631 15991 12637
rect 15933 12597 15945 12631
rect 15979 12628 15991 12631
rect 18984 12628 19012 12872
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12832 19947 12835
rect 20901 12835 20959 12841
rect 19935 12804 20668 12832
rect 19935 12801 19947 12804
rect 19889 12795 19947 12801
rect 20254 12764 20260 12776
rect 20215 12736 20260 12764
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 19705 12699 19763 12705
rect 19705 12665 19717 12699
rect 19751 12696 19763 12699
rect 20533 12699 20591 12705
rect 19751 12668 20484 12696
rect 19751 12665 19763 12668
rect 19705 12659 19763 12665
rect 15979 12600 19012 12628
rect 20456 12628 20484 12668
rect 20533 12665 20545 12699
rect 20579 12696 20591 12699
rect 20640 12696 20668 12804
rect 20901 12801 20913 12835
rect 20947 12832 20959 12835
rect 21560 12832 21588 12872
rect 25130 12860 25136 12912
rect 25188 12900 25194 12912
rect 25225 12903 25283 12909
rect 25225 12900 25237 12903
rect 25188 12872 25237 12900
rect 25188 12860 25194 12872
rect 25225 12869 25237 12872
rect 25271 12869 25283 12903
rect 25425 12903 25483 12909
rect 25425 12900 25437 12903
rect 25225 12863 25283 12869
rect 25332 12872 25437 12900
rect 23109 12835 23167 12841
rect 20947 12804 21496 12832
rect 21560 12804 22232 12832
rect 20947 12801 20959 12804
rect 20901 12795 20959 12801
rect 20990 12764 20996 12776
rect 20951 12736 20996 12764
rect 20990 12724 20996 12736
rect 21048 12724 21054 12776
rect 21082 12724 21088 12776
rect 21140 12764 21146 12776
rect 21468 12764 21496 12804
rect 22094 12764 22100 12776
rect 21140 12736 21185 12764
rect 21468 12736 22100 12764
rect 21140 12724 21146 12736
rect 22094 12724 22100 12736
rect 22152 12724 22158 12776
rect 20579 12668 20668 12696
rect 20579 12665 20591 12668
rect 20533 12659 20591 12665
rect 21358 12656 21364 12708
rect 21416 12696 21422 12708
rect 21913 12699 21971 12705
rect 21913 12696 21925 12699
rect 21416 12668 21925 12696
rect 21416 12656 21422 12668
rect 21913 12665 21925 12668
rect 21959 12665 21971 12699
rect 22204 12696 22232 12804
rect 23109 12801 23121 12835
rect 23155 12801 23167 12835
rect 23382 12832 23388 12844
rect 23343 12804 23388 12832
rect 23109 12795 23167 12801
rect 22462 12724 22468 12776
rect 22520 12764 22526 12776
rect 23124 12764 23152 12795
rect 23382 12792 23388 12804
rect 23440 12792 23446 12844
rect 23970 12835 24028 12841
rect 23970 12832 23982 12835
rect 23676 12804 23982 12832
rect 23474 12764 23480 12776
rect 22520 12736 22565 12764
rect 23124 12736 23480 12764
rect 22520 12724 22526 12736
rect 23474 12724 23480 12736
rect 23532 12724 23538 12776
rect 23014 12696 23020 12708
rect 22204 12668 23020 12696
rect 21913 12659 21971 12665
rect 23014 12656 23020 12668
rect 23072 12656 23078 12708
rect 23382 12656 23388 12708
rect 23440 12696 23446 12708
rect 23676 12696 23704 12804
rect 23970 12801 23982 12804
rect 24016 12801 24028 12835
rect 23970 12795 24028 12801
rect 24210 12792 24216 12844
rect 24268 12832 24274 12844
rect 25332 12832 25360 12872
rect 25425 12869 25437 12872
rect 25471 12869 25483 12903
rect 25425 12863 25483 12869
rect 27982 12860 27988 12912
rect 28040 12860 28046 12912
rect 30466 12860 30472 12912
rect 30524 12860 30530 12912
rect 31726 12900 31754 12940
rect 33505 12937 33517 12971
rect 33551 12968 33563 12971
rect 34425 12971 34483 12977
rect 34425 12968 34437 12971
rect 33551 12940 34437 12968
rect 33551 12937 33563 12940
rect 33505 12931 33563 12937
rect 34425 12937 34437 12940
rect 34471 12937 34483 12971
rect 35618 12968 35624 12980
rect 35579 12940 35624 12968
rect 34425 12931 34483 12937
rect 35618 12928 35624 12940
rect 35676 12928 35682 12980
rect 38378 12928 38384 12980
rect 38436 12968 38442 12980
rect 38657 12971 38715 12977
rect 38657 12968 38669 12971
rect 38436 12940 38669 12968
rect 38436 12928 38442 12940
rect 38657 12937 38669 12940
rect 38703 12937 38715 12971
rect 38657 12931 38715 12937
rect 39114 12928 39120 12980
rect 39172 12968 39178 12980
rect 39409 12971 39467 12977
rect 39409 12968 39421 12971
rect 39172 12940 39421 12968
rect 39172 12928 39178 12940
rect 39409 12937 39421 12940
rect 39455 12937 39467 12971
rect 39409 12931 39467 12937
rect 31726 12872 34008 12900
rect 26237 12835 26295 12841
rect 26237 12832 26249 12835
rect 24268 12804 26249 12832
rect 24268 12792 24274 12804
rect 26237 12801 26249 12804
rect 26283 12801 26295 12835
rect 26237 12795 26295 12801
rect 30742 12792 30748 12844
rect 30800 12832 30806 12844
rect 31573 12835 31631 12841
rect 31573 12832 31585 12835
rect 30800 12804 31585 12832
rect 30800 12792 30806 12804
rect 31573 12801 31585 12804
rect 31619 12801 31631 12835
rect 32125 12835 32183 12841
rect 32125 12832 32137 12835
rect 31573 12795 31631 12801
rect 31726 12804 32137 12832
rect 24489 12767 24547 12773
rect 24489 12733 24501 12767
rect 24535 12764 24547 12767
rect 25314 12764 25320 12776
rect 24535 12736 25320 12764
rect 24535 12733 24547 12736
rect 24489 12727 24547 12733
rect 25314 12724 25320 12736
rect 25372 12724 25378 12776
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 25424 12736 26065 12764
rect 23440 12668 23704 12696
rect 23440 12656 23446 12668
rect 24578 12656 24584 12708
rect 24636 12696 24642 12708
rect 25424 12696 25452 12736
rect 26053 12733 26065 12736
rect 26099 12733 26111 12767
rect 26053 12727 26111 12733
rect 26973 12767 27031 12773
rect 26973 12733 26985 12767
rect 27019 12733 27031 12767
rect 27246 12764 27252 12776
rect 27207 12736 27252 12764
rect 26973 12727 27031 12733
rect 24636 12668 25452 12696
rect 24636 12656 24642 12668
rect 20898 12628 20904 12640
rect 20456 12600 20904 12628
rect 15979 12597 15991 12600
rect 15933 12591 15991 12597
rect 20898 12588 20904 12600
rect 20956 12588 20962 12640
rect 22278 12588 22284 12640
rect 22336 12628 22342 12640
rect 23109 12631 23167 12637
rect 23109 12628 23121 12631
rect 22336 12600 23121 12628
rect 22336 12588 22342 12600
rect 23109 12597 23121 12600
rect 23155 12597 23167 12631
rect 23109 12591 23167 12597
rect 24397 12631 24455 12637
rect 24397 12597 24409 12631
rect 24443 12628 24455 12631
rect 25038 12628 25044 12640
rect 24443 12600 25044 12628
rect 24443 12597 24455 12600
rect 24397 12591 24455 12597
rect 25038 12588 25044 12600
rect 25096 12588 25102 12640
rect 25424 12637 25452 12668
rect 25593 12699 25651 12705
rect 25593 12665 25605 12699
rect 25639 12696 25651 12699
rect 26694 12696 26700 12708
rect 25639 12668 26700 12696
rect 25639 12665 25651 12668
rect 25593 12659 25651 12665
rect 26694 12656 26700 12668
rect 26752 12656 26758 12708
rect 25409 12631 25467 12637
rect 25409 12597 25421 12631
rect 25455 12597 25467 12631
rect 25409 12591 25467 12597
rect 26421 12631 26479 12637
rect 26421 12597 26433 12631
rect 26467 12628 26479 12631
rect 26510 12628 26516 12640
rect 26467 12600 26516 12628
rect 26467 12597 26479 12600
rect 26421 12591 26479 12597
rect 26510 12588 26516 12600
rect 26568 12588 26574 12640
rect 26786 12588 26792 12640
rect 26844 12628 26850 12640
rect 26988 12628 27016 12727
rect 27246 12724 27252 12736
rect 27304 12724 27310 12776
rect 29181 12767 29239 12773
rect 29181 12733 29193 12767
rect 29227 12733 29239 12767
rect 29454 12764 29460 12776
rect 29415 12736 29460 12764
rect 29181 12727 29239 12733
rect 29196 12696 29224 12727
rect 29454 12724 29460 12736
rect 29512 12724 29518 12776
rect 30190 12724 30196 12776
rect 30248 12764 30254 12776
rect 31726 12764 31754 12804
rect 32125 12801 32137 12804
rect 32171 12801 32183 12835
rect 32381 12835 32439 12841
rect 32381 12832 32393 12835
rect 32125 12795 32183 12801
rect 32232 12804 32393 12832
rect 32232 12764 32260 12804
rect 32381 12801 32393 12804
rect 32427 12801 32439 12835
rect 32381 12795 32439 12801
rect 30248 12736 31754 12764
rect 32048 12736 32260 12764
rect 30248 12724 30254 12736
rect 28276 12668 29224 12696
rect 28276 12628 28304 12668
rect 26844 12600 28304 12628
rect 28721 12631 28779 12637
rect 26844 12588 26850 12600
rect 28721 12597 28733 12631
rect 28767 12628 28779 12631
rect 29086 12628 29092 12640
rect 28767 12600 29092 12628
rect 28767 12597 28779 12600
rect 28721 12591 28779 12597
rect 29086 12588 29092 12600
rect 29144 12588 29150 12640
rect 29196 12628 29224 12668
rect 31389 12699 31447 12705
rect 31389 12665 31401 12699
rect 31435 12696 31447 12699
rect 32048 12696 32076 12736
rect 33980 12705 34008 12872
rect 34514 12860 34520 12912
rect 34572 12900 34578 12912
rect 39209 12903 39267 12909
rect 34572 12872 35756 12900
rect 34572 12860 34578 12872
rect 34330 12832 34336 12844
rect 34291 12804 34336 12832
rect 34330 12792 34336 12804
rect 34388 12792 34394 12844
rect 35529 12835 35587 12841
rect 35529 12801 35541 12835
rect 35575 12801 35587 12835
rect 35529 12795 35587 12801
rect 34514 12764 34520 12776
rect 34475 12736 34520 12764
rect 34514 12724 34520 12736
rect 34572 12724 34578 12776
rect 31435 12668 32076 12696
rect 33965 12699 34023 12705
rect 31435 12665 31447 12668
rect 31389 12659 31447 12665
rect 33965 12665 33977 12699
rect 34011 12665 34023 12699
rect 35544 12696 35572 12795
rect 35728 12773 35756 12872
rect 37292 12872 38976 12900
rect 35713 12767 35771 12773
rect 35713 12733 35725 12767
rect 35759 12733 35771 12767
rect 35713 12727 35771 12733
rect 36998 12724 37004 12776
rect 37056 12764 37062 12776
rect 37292 12773 37320 12872
rect 37550 12841 37556 12844
rect 37544 12795 37556 12841
rect 37608 12832 37614 12844
rect 38948 12832 38976 12872
rect 39209 12869 39221 12903
rect 39255 12900 39267 12903
rect 39758 12900 39764 12912
rect 39255 12872 39764 12900
rect 39255 12869 39267 12872
rect 39209 12863 39267 12869
rect 39758 12860 39764 12872
rect 39816 12860 39822 12912
rect 40497 12835 40555 12841
rect 40497 12832 40509 12835
rect 37608 12804 37644 12832
rect 38948 12804 40509 12832
rect 37550 12792 37556 12795
rect 37608 12792 37614 12804
rect 40497 12801 40509 12804
rect 40543 12832 40555 12835
rect 40586 12832 40592 12844
rect 40543 12804 40592 12832
rect 40543 12801 40555 12804
rect 40497 12795 40555 12801
rect 40586 12792 40592 12804
rect 40644 12792 40650 12844
rect 40764 12835 40822 12841
rect 40764 12801 40776 12835
rect 40810 12832 40822 12835
rect 42702 12832 42708 12844
rect 40810 12804 42708 12832
rect 40810 12801 40822 12804
rect 40764 12795 40822 12801
rect 42702 12792 42708 12804
rect 42760 12792 42766 12844
rect 37277 12767 37335 12773
rect 37277 12764 37289 12767
rect 37056 12736 37289 12764
rect 37056 12724 37062 12736
rect 37277 12733 37289 12736
rect 37323 12733 37335 12767
rect 40034 12764 40040 12776
rect 37277 12727 37335 12733
rect 38304 12736 40040 12764
rect 33965 12659 34023 12665
rect 34072 12668 35572 12696
rect 30190 12628 30196 12640
rect 29196 12600 30196 12628
rect 30190 12588 30196 12600
rect 30248 12588 30254 12640
rect 30466 12588 30472 12640
rect 30524 12628 30530 12640
rect 30929 12631 30987 12637
rect 30929 12628 30941 12631
rect 30524 12600 30941 12628
rect 30524 12588 30530 12600
rect 30929 12597 30941 12600
rect 30975 12597 30987 12631
rect 30929 12591 30987 12597
rect 33594 12588 33600 12640
rect 33652 12628 33658 12640
rect 34072 12628 34100 12668
rect 33652 12600 34100 12628
rect 35161 12631 35219 12637
rect 33652 12588 33658 12600
rect 35161 12597 35173 12631
rect 35207 12628 35219 12631
rect 38304 12628 38332 12736
rect 40034 12724 40040 12736
rect 40092 12724 40098 12776
rect 38562 12656 38568 12708
rect 38620 12696 38626 12708
rect 38620 12668 39436 12696
rect 38620 12656 38626 12668
rect 39408 12637 39436 12668
rect 35207 12600 38332 12628
rect 39393 12631 39451 12637
rect 35207 12597 35219 12600
rect 35161 12591 35219 12597
rect 39393 12597 39405 12631
rect 39439 12597 39451 12631
rect 39393 12591 39451 12597
rect 39577 12631 39635 12637
rect 39577 12597 39589 12631
rect 39623 12628 39635 12631
rect 39666 12628 39672 12640
rect 39623 12600 39672 12628
rect 39623 12597 39635 12600
rect 39577 12591 39635 12597
rect 39666 12588 39672 12600
rect 39724 12588 39730 12640
rect 41877 12631 41935 12637
rect 41877 12597 41889 12631
rect 41923 12628 41935 12631
rect 41966 12628 41972 12640
rect 41923 12600 41972 12628
rect 41923 12597 41935 12600
rect 41877 12591 41935 12597
rect 41966 12588 41972 12600
rect 42024 12588 42030 12640
rect 44082 12588 44088 12640
rect 44140 12628 44146 12640
rect 44177 12631 44235 12637
rect 44177 12628 44189 12631
rect 44140 12600 44189 12628
rect 44140 12588 44146 12600
rect 44177 12597 44189 12600
rect 44223 12597 44235 12631
rect 44177 12591 44235 12597
rect 1104 12538 44896 12560
rect 1104 12486 6424 12538
rect 6476 12486 6488 12538
rect 6540 12486 6552 12538
rect 6604 12486 6616 12538
rect 6668 12486 6680 12538
rect 6732 12486 17372 12538
rect 17424 12486 17436 12538
rect 17488 12486 17500 12538
rect 17552 12486 17564 12538
rect 17616 12486 17628 12538
rect 17680 12486 28320 12538
rect 28372 12486 28384 12538
rect 28436 12486 28448 12538
rect 28500 12486 28512 12538
rect 28564 12486 28576 12538
rect 28628 12486 39268 12538
rect 39320 12486 39332 12538
rect 39384 12486 39396 12538
rect 39448 12486 39460 12538
rect 39512 12486 39524 12538
rect 39576 12486 44896 12538
rect 1104 12464 44896 12486
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 6089 12427 6147 12433
rect 6089 12424 6101 12427
rect 5500 12396 6101 12424
rect 5500 12384 5506 12396
rect 6089 12393 6101 12396
rect 6135 12424 6147 12427
rect 12066 12424 12072 12436
rect 6135 12396 12072 12424
rect 6135 12393 6147 12396
rect 6089 12387 6147 12393
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 12250 12384 12256 12436
rect 12308 12424 12314 12436
rect 14185 12427 14243 12433
rect 12308 12396 14136 12424
rect 12308 12384 12314 12396
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 8260 12328 10088 12356
rect 8260 12316 8266 12328
rect 4430 12248 4436 12300
rect 4488 12288 4494 12300
rect 4709 12291 4767 12297
rect 4709 12288 4721 12291
rect 4488 12260 4721 12288
rect 4488 12248 4494 12260
rect 4709 12257 4721 12260
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 9953 12291 10011 12297
rect 9953 12288 9965 12291
rect 9640 12260 9965 12288
rect 9640 12248 9646 12260
rect 9953 12257 9965 12260
rect 9999 12257 10011 12291
rect 10060 12288 10088 12328
rect 12342 12316 12348 12368
rect 12400 12356 12406 12368
rect 12400 12328 13676 12356
rect 12400 12316 12406 12328
rect 11057 12291 11115 12297
rect 11057 12288 11069 12291
rect 10060 12260 11069 12288
rect 9953 12251 10011 12257
rect 11057 12257 11069 12260
rect 11103 12257 11115 12291
rect 11057 12251 11115 12257
rect 12526 12248 12532 12300
rect 12584 12288 12590 12300
rect 13648 12288 13676 12328
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 14108 12356 14136 12396
rect 14185 12393 14197 12427
rect 14231 12424 14243 12427
rect 14642 12424 14648 12436
rect 14231 12396 14648 12424
rect 14231 12393 14243 12396
rect 14185 12387 14243 12393
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 14921 12427 14979 12433
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 15470 12424 15476 12436
rect 14967 12396 15476 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 15764 12396 21680 12424
rect 15764 12356 15792 12396
rect 16482 12356 16488 12368
rect 13780 12328 13952 12356
rect 14108 12328 15792 12356
rect 15856 12328 16488 12356
rect 13780 12316 13786 12328
rect 13924 12288 13952 12328
rect 15749 12291 15807 12297
rect 12584 12260 13584 12288
rect 13648 12260 13768 12288
rect 13924 12260 14320 12288
rect 12584 12248 12590 12260
rect 13556 12232 13584 12260
rect 2590 12220 2596 12232
rect 2551 12192 2596 12220
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 2682 12180 2688 12232
rect 2740 12220 2746 12232
rect 4157 12223 4215 12229
rect 4157 12220 4169 12223
rect 2740 12192 4169 12220
rect 2740 12180 2746 12192
rect 4157 12189 4169 12192
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 6822 12220 6828 12232
rect 6687 12192 6828 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12220 8447 12223
rect 8846 12220 8852 12232
rect 8435 12192 8852 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 8938 12180 8944 12232
rect 8996 12220 9002 12232
rect 10778 12220 10784 12232
rect 8996 12192 10784 12220
rect 8996 12180 9002 12192
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12220 13047 12223
rect 13078 12220 13084 12232
rect 13035 12192 13084 12220
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 13078 12180 13084 12192
rect 13136 12180 13142 12232
rect 13538 12180 13544 12232
rect 13596 12180 13602 12232
rect 4976 12155 5034 12161
rect 4976 12121 4988 12155
rect 5022 12152 5034 12155
rect 6546 12152 6552 12164
rect 5022 12124 6552 12152
rect 5022 12121 5034 12124
rect 4976 12115 5034 12121
rect 6546 12112 6552 12124
rect 6604 12112 6610 12164
rect 9769 12155 9827 12161
rect 9769 12121 9781 12155
rect 9815 12152 9827 12155
rect 10318 12152 10324 12164
rect 9815 12124 10324 12152
rect 9815 12121 9827 12124
rect 9769 12115 9827 12121
rect 10318 12112 10324 12124
rect 10376 12112 10382 12164
rect 11514 12112 11520 12164
rect 11572 12112 11578 12164
rect 13740 12152 13768 12260
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 14292 12229 14320 12260
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 15856 12288 15884 12328
rect 16482 12316 16488 12328
rect 16540 12316 16546 12368
rect 16945 12359 17003 12365
rect 16945 12325 16957 12359
rect 16991 12356 17003 12359
rect 17770 12356 17776 12368
rect 16991 12328 17776 12356
rect 16991 12325 17003 12328
rect 16945 12319 17003 12325
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 20438 12356 20444 12368
rect 18064 12328 20444 12356
rect 16022 12288 16028 12300
rect 15795 12260 15884 12288
rect 15983 12260 16028 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 16022 12248 16028 12260
rect 16080 12248 16086 12300
rect 16234 12291 16292 12297
rect 16234 12257 16246 12291
rect 16280 12288 16292 12291
rect 18064 12288 18092 12328
rect 20438 12316 20444 12328
rect 20496 12316 20502 12368
rect 21652 12356 21680 12396
rect 22094 12384 22100 12436
rect 22152 12424 22158 12436
rect 22327 12427 22385 12433
rect 22327 12424 22339 12427
rect 22152 12396 22339 12424
rect 22152 12384 22158 12396
rect 22327 12393 22339 12396
rect 22373 12424 22385 12427
rect 23198 12424 23204 12436
rect 22373 12396 23204 12424
rect 22373 12393 22385 12396
rect 22327 12387 22385 12393
rect 23198 12384 23204 12396
rect 23256 12384 23262 12436
rect 23661 12427 23719 12433
rect 23661 12393 23673 12427
rect 23707 12424 23719 12427
rect 24210 12424 24216 12436
rect 23707 12396 24216 12424
rect 23707 12393 23719 12396
rect 23661 12387 23719 12393
rect 24210 12384 24216 12396
rect 24268 12384 24274 12436
rect 24578 12424 24584 12436
rect 24539 12396 24584 12424
rect 24578 12384 24584 12396
rect 24636 12384 24642 12436
rect 25222 12424 25228 12436
rect 25183 12396 25228 12424
rect 25222 12384 25228 12396
rect 25280 12384 25286 12436
rect 25314 12384 25320 12436
rect 25372 12424 25378 12436
rect 25685 12427 25743 12433
rect 25685 12424 25697 12427
rect 25372 12396 25697 12424
rect 25372 12384 25378 12396
rect 25685 12393 25697 12396
rect 25731 12393 25743 12427
rect 25685 12387 25743 12393
rect 26326 12384 26332 12436
rect 26384 12424 26390 12436
rect 26421 12427 26479 12433
rect 26421 12424 26433 12427
rect 26384 12396 26433 12424
rect 26384 12384 26390 12396
rect 26421 12393 26433 12396
rect 26467 12393 26479 12427
rect 27798 12424 27804 12436
rect 27759 12396 27804 12424
rect 26421 12387 26479 12393
rect 27798 12384 27804 12396
rect 27856 12384 27862 12436
rect 28813 12427 28871 12433
rect 28813 12393 28825 12427
rect 28859 12424 28871 12427
rect 29086 12424 29092 12436
rect 28859 12396 29092 12424
rect 28859 12393 28871 12396
rect 28813 12387 28871 12393
rect 29086 12384 29092 12396
rect 29144 12384 29150 12436
rect 29454 12384 29460 12436
rect 29512 12424 29518 12436
rect 29549 12427 29607 12433
rect 29549 12424 29561 12427
rect 29512 12396 29561 12424
rect 29512 12384 29518 12396
rect 29549 12393 29561 12396
rect 29595 12393 29607 12427
rect 29549 12387 29607 12393
rect 29914 12384 29920 12436
rect 29972 12424 29978 12436
rect 30466 12424 30472 12436
rect 29972 12396 30472 12424
rect 29972 12384 29978 12396
rect 30466 12384 30472 12396
rect 30524 12384 30530 12436
rect 30558 12384 30564 12436
rect 30616 12424 30622 12436
rect 33134 12424 33140 12436
rect 30616 12396 33140 12424
rect 30616 12384 30622 12396
rect 33134 12384 33140 12396
rect 33192 12384 33198 12436
rect 33229 12427 33287 12433
rect 33229 12393 33241 12427
rect 33275 12424 33287 12427
rect 34330 12424 34336 12436
rect 33275 12396 34336 12424
rect 33275 12393 33287 12396
rect 33229 12387 33287 12393
rect 34330 12384 34336 12396
rect 34388 12384 34394 12436
rect 37734 12424 37740 12436
rect 36188 12396 37740 12424
rect 22554 12356 22560 12368
rect 21652 12328 22560 12356
rect 22554 12316 22560 12328
rect 22612 12316 22618 12368
rect 24670 12316 24676 12368
rect 24728 12356 24734 12368
rect 26234 12356 26240 12368
rect 24728 12328 26240 12356
rect 24728 12316 24734 12328
rect 26234 12316 26240 12328
rect 26292 12316 26298 12368
rect 28997 12359 29055 12365
rect 26344 12328 27844 12356
rect 16280 12260 18092 12288
rect 18141 12291 18199 12297
rect 16280 12257 16292 12260
rect 16234 12251 16292 12257
rect 18141 12257 18153 12291
rect 18187 12288 18199 12291
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 18187 12260 19809 12288
rect 18187 12257 18199 12260
rect 18141 12251 18199 12257
rect 19797 12257 19809 12260
rect 19843 12288 19855 12291
rect 20346 12288 20352 12300
rect 19843 12260 20352 12288
rect 19843 12257 19855 12260
rect 19797 12251 19855 12257
rect 20346 12248 20352 12260
rect 20404 12288 20410 12300
rect 20898 12288 20904 12300
rect 20404 12260 20760 12288
rect 20859 12260 20904 12288
rect 20404 12248 20410 12260
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13964 12192 14105 12220
rect 13964 12180 13970 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12189 14335 12223
rect 14826 12220 14832 12232
rect 14787 12192 14832 12220
rect 14277 12183 14335 12189
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 16117 12223 16175 12229
rect 16117 12220 16129 12223
rect 15896 12192 16129 12220
rect 15896 12180 15902 12192
rect 16117 12189 16129 12192
rect 16163 12189 16175 12223
rect 16758 12220 16764 12232
rect 16117 12183 16175 12189
rect 16224 12192 16764 12220
rect 16224 12152 16252 12192
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 16850 12180 16856 12232
rect 16908 12220 16914 12232
rect 17862 12220 17868 12232
rect 16908 12192 16953 12220
rect 17823 12192 17868 12220
rect 16908 12180 16914 12192
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 18414 12180 18420 12232
rect 18472 12220 18478 12232
rect 19150 12220 19156 12232
rect 18472 12192 19156 12220
rect 18472 12180 18478 12192
rect 19150 12180 19156 12192
rect 19208 12220 19214 12232
rect 19613 12223 19671 12229
rect 19613 12220 19625 12223
rect 19208 12192 19625 12220
rect 19208 12180 19214 12192
rect 19613 12189 19625 12192
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 20533 12223 20591 12229
rect 20533 12189 20545 12223
rect 20579 12220 20591 12223
rect 20622 12220 20628 12232
rect 20579 12192 20628 12220
rect 20579 12189 20591 12192
rect 20533 12183 20591 12189
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 20732 12220 20760 12260
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 22462 12288 22468 12300
rect 21008 12260 22468 12288
rect 21008 12220 21036 12260
rect 22462 12248 22468 12260
rect 22520 12248 22526 12300
rect 25222 12248 25228 12300
rect 25280 12288 25286 12300
rect 26344 12288 26372 12328
rect 25280 12260 26372 12288
rect 25280 12248 25286 12260
rect 26510 12248 26516 12300
rect 26568 12288 26574 12300
rect 27065 12291 27123 12297
rect 27065 12288 27077 12291
rect 26568 12260 27077 12288
rect 26568 12248 26574 12260
rect 27065 12257 27077 12260
rect 27111 12288 27123 12291
rect 27430 12288 27436 12300
rect 27111 12260 27436 12288
rect 27111 12257 27123 12260
rect 27065 12251 27123 12257
rect 27430 12248 27436 12260
rect 27488 12248 27494 12300
rect 20732 12192 21036 12220
rect 23014 12180 23020 12232
rect 23072 12220 23078 12232
rect 23201 12223 23259 12229
rect 23201 12220 23213 12223
rect 23072 12192 23213 12220
rect 23072 12180 23078 12192
rect 23201 12189 23213 12192
rect 23247 12220 23259 12223
rect 23382 12220 23388 12232
rect 23247 12192 23388 12220
rect 23247 12189 23259 12192
rect 23201 12183 23259 12189
rect 23382 12180 23388 12192
rect 23440 12180 23446 12232
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12220 23903 12223
rect 24026 12220 24032 12232
rect 23891 12192 24032 12220
rect 23891 12189 23903 12192
rect 23845 12183 23903 12189
rect 13740 12124 16252 12152
rect 16408 12124 19932 12152
rect 2958 12044 2964 12096
rect 3016 12084 3022 12096
rect 3237 12087 3295 12093
rect 3237 12084 3249 12087
rect 3016 12056 3249 12084
rect 3016 12044 3022 12056
rect 3237 12053 3249 12056
rect 3283 12053 3295 12087
rect 3237 12047 3295 12053
rect 3878 12044 3884 12096
rect 3936 12084 3942 12096
rect 3973 12087 4031 12093
rect 3973 12084 3985 12087
rect 3936 12056 3985 12084
rect 3936 12044 3942 12056
rect 3973 12053 3985 12056
rect 4019 12053 4031 12087
rect 7190 12084 7196 12096
rect 7151 12056 7196 12084
rect 3973 12047 4031 12053
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 8205 12087 8263 12093
rect 8205 12053 8217 12087
rect 8251 12084 8263 12087
rect 9214 12084 9220 12096
rect 8251 12056 9220 12084
rect 8251 12053 8263 12056
rect 8205 12047 8263 12053
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 9398 12084 9404 12096
rect 9359 12056 9404 12084
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 9858 12044 9864 12096
rect 9916 12084 9922 12096
rect 9916 12056 9961 12084
rect 9916 12044 9922 12056
rect 10226 12044 10232 12096
rect 10284 12084 10290 12096
rect 12342 12084 12348 12096
rect 10284 12056 12348 12084
rect 10284 12044 10290 12056
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12618 12044 12624 12096
rect 12676 12084 12682 12096
rect 16408 12093 16436 12124
rect 13173 12087 13231 12093
rect 13173 12084 13185 12087
rect 12676 12056 13185 12084
rect 12676 12044 12682 12056
rect 13173 12053 13185 12056
rect 13219 12053 13231 12087
rect 13173 12047 13231 12053
rect 16393 12087 16451 12093
rect 16393 12053 16405 12087
rect 16439 12053 16451 12087
rect 16393 12047 16451 12053
rect 17218 12044 17224 12096
rect 17276 12084 17282 12096
rect 17497 12087 17555 12093
rect 17497 12084 17509 12087
rect 17276 12056 17509 12084
rect 17276 12044 17282 12056
rect 17497 12053 17509 12056
rect 17543 12053 17555 12087
rect 17497 12047 17555 12053
rect 17586 12044 17592 12096
rect 17644 12084 17650 12096
rect 17954 12084 17960 12096
rect 17644 12056 17960 12084
rect 17644 12044 17650 12056
rect 17954 12044 17960 12056
rect 18012 12044 18018 12096
rect 18046 12044 18052 12096
rect 18104 12084 18110 12096
rect 19245 12087 19303 12093
rect 19245 12084 19257 12087
rect 18104 12056 19257 12084
rect 18104 12044 18110 12056
rect 19245 12053 19257 12056
rect 19291 12053 19303 12087
rect 19245 12047 19303 12053
rect 19705 12087 19763 12093
rect 19705 12053 19717 12087
rect 19751 12084 19763 12087
rect 19794 12084 19800 12096
rect 19751 12056 19800 12084
rect 19751 12053 19763 12056
rect 19705 12047 19763 12053
rect 19794 12044 19800 12056
rect 19852 12044 19858 12096
rect 19904 12084 19932 12124
rect 21266 12112 21272 12164
rect 21324 12112 21330 12164
rect 23860 12152 23888 12183
rect 24026 12180 24032 12192
rect 24084 12180 24090 12232
rect 25409 12223 25467 12229
rect 25409 12220 25421 12223
rect 24412 12192 25421 12220
rect 24412 12161 24440 12192
rect 25409 12189 25421 12192
rect 25455 12189 25467 12223
rect 25409 12183 25467 12189
rect 25501 12223 25559 12229
rect 25501 12189 25513 12223
rect 25547 12220 25559 12223
rect 26881 12223 26939 12229
rect 26881 12220 26893 12223
rect 25547 12192 26893 12220
rect 25547 12189 25559 12192
rect 25501 12183 25559 12189
rect 26881 12189 26893 12192
rect 26927 12189 26939 12223
rect 26881 12183 26939 12189
rect 22066 12124 23888 12152
rect 24397 12155 24455 12161
rect 22066 12084 22094 12124
rect 24397 12121 24409 12155
rect 24443 12121 24455 12155
rect 24397 12115 24455 12121
rect 24486 12112 24492 12164
rect 24544 12152 24550 12164
rect 25225 12155 25283 12161
rect 25225 12152 25237 12155
rect 24544 12124 25237 12152
rect 24544 12112 24550 12124
rect 25225 12121 25237 12124
rect 25271 12121 25283 12155
rect 25424 12152 25452 12183
rect 26418 12152 26424 12164
rect 25424 12124 26424 12152
rect 25225 12115 25283 12121
rect 26418 12112 26424 12124
rect 26476 12112 26482 12164
rect 26896 12152 26924 12183
rect 27614 12180 27620 12232
rect 27672 12220 27678 12232
rect 27709 12223 27767 12229
rect 27709 12220 27721 12223
rect 27672 12192 27721 12220
rect 27672 12180 27678 12192
rect 27709 12189 27721 12192
rect 27755 12189 27767 12223
rect 27816 12220 27844 12328
rect 28997 12325 29009 12359
rect 29043 12356 29055 12359
rect 30742 12356 30748 12368
rect 29043 12328 30748 12356
rect 29043 12325 29055 12328
rect 28997 12319 29055 12325
rect 30742 12316 30748 12328
rect 30800 12316 30806 12368
rect 31294 12288 31300 12300
rect 30024 12260 31300 12288
rect 30024 12232 30052 12260
rect 31294 12248 31300 12260
rect 31352 12248 31358 12300
rect 33873 12291 33931 12297
rect 33873 12257 33885 12291
rect 33919 12288 33931 12291
rect 34238 12288 34244 12300
rect 33919 12260 34244 12288
rect 33919 12257 33931 12260
rect 33873 12251 33931 12257
rect 34238 12248 34244 12260
rect 34296 12248 34302 12300
rect 36188 12297 36216 12396
rect 37734 12384 37740 12396
rect 37792 12384 37798 12436
rect 40494 12424 40500 12436
rect 40328 12396 40500 12424
rect 38010 12316 38016 12368
rect 38068 12356 38074 12368
rect 39850 12356 39856 12368
rect 38068 12328 39856 12356
rect 38068 12316 38074 12328
rect 39850 12316 39856 12328
rect 39908 12316 39914 12368
rect 36173 12291 36231 12297
rect 36173 12257 36185 12291
rect 36219 12257 36231 12291
rect 36538 12288 36544 12300
rect 36451 12260 36544 12288
rect 36173 12251 36231 12257
rect 36538 12248 36544 12260
rect 36596 12288 36602 12300
rect 40328 12297 40356 12396
rect 40494 12384 40500 12396
rect 40552 12384 40558 12436
rect 42702 12384 42708 12436
rect 42760 12424 42766 12436
rect 42889 12427 42947 12433
rect 42889 12424 42901 12427
rect 42760 12396 42901 12424
rect 42760 12384 42766 12396
rect 42889 12393 42901 12396
rect 42935 12393 42947 12427
rect 42889 12387 42947 12393
rect 40402 12316 40408 12368
rect 40460 12356 40466 12368
rect 40460 12328 40540 12356
rect 40460 12316 40466 12328
rect 40512 12297 40540 12328
rect 40314 12291 40372 12297
rect 36596 12260 37136 12288
rect 36596 12248 36602 12260
rect 28629 12223 28687 12229
rect 28629 12220 28641 12223
rect 27816 12192 28641 12220
rect 27709 12183 27767 12189
rect 28629 12189 28641 12192
rect 28675 12189 28687 12223
rect 28629 12183 28687 12189
rect 28721 12223 28779 12229
rect 28721 12189 28733 12223
rect 28767 12189 28779 12223
rect 28721 12183 28779 12189
rect 28736 12152 28764 12183
rect 29086 12180 29092 12232
rect 29144 12220 29150 12232
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 29144 12192 29745 12220
rect 29144 12180 29150 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 30006 12220 30012 12232
rect 29967 12192 30012 12220
rect 29733 12183 29791 12189
rect 26896 12124 28764 12152
rect 29748 12152 29776 12183
rect 30006 12180 30012 12192
rect 30064 12180 30070 12232
rect 30282 12180 30288 12232
rect 30340 12220 30346 12232
rect 31021 12223 31079 12229
rect 31021 12220 31033 12223
rect 30340 12192 31033 12220
rect 30340 12180 30346 12192
rect 31021 12189 31033 12192
rect 31067 12189 31079 12223
rect 31021 12183 31079 12189
rect 33318 12180 33324 12232
rect 33376 12220 33382 12232
rect 33597 12223 33655 12229
rect 33597 12220 33609 12223
rect 33376 12192 33609 12220
rect 33376 12180 33382 12192
rect 33597 12189 33609 12192
rect 33643 12189 33655 12223
rect 33597 12183 33655 12189
rect 33689 12223 33747 12229
rect 33689 12189 33701 12223
rect 33735 12220 33747 12223
rect 34146 12220 34152 12232
rect 33735 12192 34152 12220
rect 33735 12189 33747 12192
rect 33689 12183 33747 12189
rect 34146 12180 34152 12192
rect 34204 12180 34210 12232
rect 36357 12223 36415 12229
rect 36357 12189 36369 12223
rect 36403 12189 36415 12223
rect 36998 12220 37004 12232
rect 36959 12192 37004 12220
rect 36357 12183 36415 12189
rect 29748 12124 30052 12152
rect 19904 12056 22094 12084
rect 23017 12087 23075 12093
rect 23017 12053 23029 12087
rect 23063 12084 23075 12087
rect 23474 12084 23480 12096
rect 23063 12056 23480 12084
rect 23063 12053 23075 12056
rect 23017 12047 23075 12053
rect 23474 12044 23480 12056
rect 23532 12044 23538 12096
rect 24210 12044 24216 12096
rect 24268 12084 24274 12096
rect 24597 12087 24655 12093
rect 24597 12084 24609 12087
rect 24268 12056 24609 12084
rect 24268 12044 24274 12056
rect 24597 12053 24609 12056
rect 24643 12053 24655 12087
rect 24762 12084 24768 12096
rect 24723 12056 24768 12084
rect 24597 12047 24655 12053
rect 24762 12044 24768 12056
rect 24820 12044 24826 12096
rect 25038 12044 25044 12096
rect 25096 12084 25102 12096
rect 26789 12087 26847 12093
rect 26789 12084 26801 12087
rect 25096 12056 26801 12084
rect 25096 12044 25102 12056
rect 26789 12053 26801 12056
rect 26835 12084 26847 12087
rect 28626 12084 28632 12096
rect 26835 12056 28632 12084
rect 26835 12053 26847 12056
rect 26789 12047 26847 12053
rect 28626 12044 28632 12056
rect 28684 12044 28690 12096
rect 28736 12084 28764 12124
rect 29914 12084 29920 12096
rect 28736 12056 29920 12084
rect 29914 12044 29920 12056
rect 29972 12044 29978 12096
rect 30024 12084 30052 12124
rect 30190 12112 30196 12164
rect 30248 12152 30254 12164
rect 30374 12152 30380 12164
rect 30248 12124 30380 12152
rect 30248 12112 30254 12124
rect 30374 12112 30380 12124
rect 30432 12112 30438 12164
rect 30650 12112 30656 12164
rect 30708 12152 30714 12164
rect 31297 12155 31355 12161
rect 31297 12152 31309 12155
rect 30708 12124 31309 12152
rect 30708 12112 30714 12124
rect 31297 12121 31309 12124
rect 31343 12121 31355 12155
rect 33502 12152 33508 12164
rect 32522 12124 33508 12152
rect 31297 12115 31355 12121
rect 33502 12112 33508 12124
rect 33560 12112 33566 12164
rect 30742 12084 30748 12096
rect 30024 12056 30748 12084
rect 30742 12044 30748 12056
rect 30800 12044 30806 12096
rect 31202 12044 31208 12096
rect 31260 12084 31266 12096
rect 32769 12087 32827 12093
rect 32769 12084 32781 12087
rect 31260 12056 32781 12084
rect 31260 12044 31266 12056
rect 32769 12053 32781 12056
rect 32815 12053 32827 12087
rect 36372 12084 36400 12183
rect 36998 12180 37004 12192
rect 37056 12180 37062 12232
rect 37108 12220 37136 12260
rect 38028 12260 39252 12288
rect 38028 12220 38056 12260
rect 39022 12220 39028 12232
rect 37108 12192 38056 12220
rect 38983 12192 39028 12220
rect 39022 12180 39028 12192
rect 39080 12180 39086 12232
rect 39224 12229 39252 12260
rect 40314 12257 40326 12291
rect 40360 12257 40372 12291
rect 40314 12251 40372 12257
rect 40497 12291 40555 12297
rect 40497 12257 40509 12291
rect 40543 12257 40555 12291
rect 40497 12251 40555 12257
rect 40586 12248 40592 12300
rect 40644 12288 40650 12300
rect 41049 12291 41107 12297
rect 41049 12288 41061 12291
rect 40644 12260 41061 12288
rect 40644 12248 40650 12260
rect 41049 12257 41061 12260
rect 41095 12257 41107 12291
rect 41049 12251 41107 12257
rect 42610 12248 42616 12300
rect 42668 12288 42674 12300
rect 42668 12260 43116 12288
rect 42668 12248 42674 12260
rect 39209 12223 39267 12229
rect 39209 12189 39221 12223
rect 39255 12189 39267 12223
rect 39209 12183 39267 12189
rect 39298 12180 39304 12232
rect 39356 12220 39362 12232
rect 39356 12192 39401 12220
rect 39356 12180 39362 12192
rect 39666 12180 39672 12232
rect 39724 12220 39730 12232
rect 43088 12229 43116 12260
rect 40222 12223 40280 12229
rect 39724 12214 40172 12220
rect 40222 12214 40234 12223
rect 39724 12192 40234 12214
rect 39724 12180 39730 12192
rect 40144 12189 40234 12192
rect 40268 12189 40280 12223
rect 40144 12186 40280 12189
rect 40222 12183 40280 12186
rect 40405 12223 40463 12229
rect 40405 12189 40417 12223
rect 40451 12189 40463 12223
rect 42889 12223 42947 12229
rect 42889 12220 42901 12223
rect 40405 12183 40463 12189
rect 41386 12192 42901 12220
rect 37268 12155 37326 12161
rect 37268 12121 37280 12155
rect 37314 12121 37326 12155
rect 38841 12155 38899 12161
rect 38841 12152 38853 12155
rect 37268 12115 37326 12121
rect 37476 12124 38853 12152
rect 37182 12084 37188 12096
rect 36372 12056 37188 12084
rect 32769 12047 32827 12053
rect 37182 12044 37188 12056
rect 37240 12044 37246 12096
rect 37292 12084 37320 12115
rect 37476 12084 37504 12124
rect 38841 12121 38853 12124
rect 38887 12121 38899 12155
rect 38841 12115 38899 12121
rect 39850 12112 39856 12164
rect 39908 12152 39914 12164
rect 40310 12152 40316 12164
rect 39908 12124 40316 12152
rect 39908 12112 39914 12124
rect 40310 12112 40316 12124
rect 40368 12112 40374 12164
rect 40420 12152 40448 12183
rect 40770 12152 40776 12164
rect 40420 12124 40776 12152
rect 40770 12112 40776 12124
rect 40828 12112 40834 12164
rect 41046 12112 41052 12164
rect 41104 12152 41110 12164
rect 41294 12155 41352 12161
rect 41294 12152 41306 12155
rect 41104 12124 41306 12152
rect 41104 12112 41110 12124
rect 41294 12121 41306 12124
rect 41340 12121 41352 12155
rect 41294 12115 41352 12121
rect 37292 12056 37504 12084
rect 38286 12044 38292 12096
rect 38344 12084 38350 12096
rect 38381 12087 38439 12093
rect 38381 12084 38393 12087
rect 38344 12056 38393 12084
rect 38344 12044 38350 12056
rect 38381 12053 38393 12056
rect 38427 12084 38439 12087
rect 39298 12084 39304 12096
rect 38427 12056 39304 12084
rect 38427 12053 38439 12056
rect 38381 12047 38439 12053
rect 39298 12044 39304 12056
rect 39356 12044 39362 12096
rect 40037 12087 40095 12093
rect 40037 12053 40049 12087
rect 40083 12084 40095 12087
rect 41386 12084 41414 12192
rect 42889 12189 42901 12192
rect 42935 12189 42947 12223
rect 42889 12183 42947 12189
rect 43073 12223 43131 12229
rect 43073 12189 43085 12223
rect 43119 12189 43131 12223
rect 43073 12183 43131 12189
rect 42426 12084 42432 12096
rect 40083 12056 41414 12084
rect 42387 12056 42432 12084
rect 40083 12053 40095 12056
rect 40037 12047 40095 12053
rect 42426 12044 42432 12056
rect 42484 12044 42490 12096
rect 1104 11994 45056 12016
rect 1104 11942 11898 11994
rect 11950 11942 11962 11994
rect 12014 11942 12026 11994
rect 12078 11942 12090 11994
rect 12142 11942 12154 11994
rect 12206 11942 22846 11994
rect 22898 11942 22910 11994
rect 22962 11942 22974 11994
rect 23026 11942 23038 11994
rect 23090 11942 23102 11994
rect 23154 11942 33794 11994
rect 33846 11942 33858 11994
rect 33910 11942 33922 11994
rect 33974 11942 33986 11994
rect 34038 11942 34050 11994
rect 34102 11942 44742 11994
rect 44794 11942 44806 11994
rect 44858 11942 44870 11994
rect 44922 11942 44934 11994
rect 44986 11942 44998 11994
rect 45050 11942 45056 11994
rect 1104 11920 45056 11942
rect 2590 11840 2596 11892
rect 2648 11880 2654 11892
rect 4433 11883 4491 11889
rect 4433 11880 4445 11883
rect 2648 11852 4445 11880
rect 2648 11840 2654 11852
rect 4433 11849 4445 11852
rect 4479 11880 4491 11883
rect 4614 11880 4620 11892
rect 4479 11852 4620 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 5077 11883 5135 11889
rect 5077 11849 5089 11883
rect 5123 11849 5135 11883
rect 5442 11880 5448 11892
rect 5403 11852 5448 11880
rect 5077 11843 5135 11849
rect 3694 11812 3700 11824
rect 3068 11784 3700 11812
rect 3068 11753 3096 11784
rect 3694 11772 3700 11784
rect 3752 11772 3758 11824
rect 5092 11812 5120 11843
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 5537 11883 5595 11889
rect 5537 11849 5549 11883
rect 5583 11880 5595 11883
rect 7190 11880 7196 11892
rect 5583 11852 7196 11880
rect 5583 11849 5595 11852
rect 5537 11843 5595 11849
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 9916 11852 13461 11880
rect 9916 11840 9922 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 17034 11880 17040 11892
rect 16995 11852 17040 11880
rect 13449 11843 13507 11849
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 19150 11840 19156 11892
rect 19208 11880 19214 11892
rect 19613 11883 19671 11889
rect 19613 11880 19625 11883
rect 19208 11852 19625 11880
rect 19208 11840 19214 11852
rect 19613 11849 19625 11852
rect 19659 11849 19671 11883
rect 19613 11843 19671 11849
rect 19702 11840 19708 11892
rect 19760 11880 19766 11892
rect 20441 11883 20499 11889
rect 20441 11880 20453 11883
rect 19760 11852 20453 11880
rect 19760 11840 19766 11852
rect 20441 11849 20453 11852
rect 20487 11880 20499 11883
rect 21082 11880 21088 11892
rect 20487 11852 21088 11880
rect 20487 11849 20499 11852
rect 20441 11843 20499 11849
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 21177 11883 21235 11889
rect 21177 11849 21189 11883
rect 21223 11880 21235 11883
rect 21266 11880 21272 11892
rect 21223 11852 21272 11880
rect 21223 11849 21235 11852
rect 21177 11843 21235 11849
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 22649 11883 22707 11889
rect 22649 11849 22661 11883
rect 22695 11880 22707 11883
rect 22738 11880 22744 11892
rect 22695 11852 22744 11880
rect 22695 11849 22707 11852
rect 22649 11843 22707 11849
rect 22738 11840 22744 11852
rect 22796 11840 22802 11892
rect 23768 11852 26280 11880
rect 9214 11812 9220 11824
rect 5092 11784 6776 11812
rect 9175 11784 9220 11812
rect 6748 11753 6776 11784
rect 9214 11772 9220 11784
rect 9272 11772 9278 11824
rect 10594 11812 10600 11824
rect 10442 11784 10600 11812
rect 10594 11772 10600 11784
rect 10652 11772 10658 11824
rect 11977 11815 12035 11821
rect 11977 11781 11989 11815
rect 12023 11812 12035 11815
rect 12526 11812 12532 11824
rect 12023 11784 12532 11812
rect 12023 11781 12035 11784
rect 11977 11775 12035 11781
rect 12526 11772 12532 11784
rect 12584 11772 12590 11824
rect 18230 11812 18236 11824
rect 14292 11784 18236 11812
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 3320 11747 3378 11753
rect 3320 11713 3332 11747
rect 3366 11744 3378 11747
rect 6733 11747 6791 11753
rect 3366 11716 6684 11744
rect 3366 11713 3378 11716
rect 3320 11707 3378 11713
rect 4246 11636 4252 11688
rect 4304 11676 4310 11688
rect 5721 11679 5779 11685
rect 5721 11676 5733 11679
rect 4304 11648 5733 11676
rect 4304 11636 4310 11648
rect 5721 11645 5733 11648
rect 5767 11676 5779 11679
rect 5767 11648 6408 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 6086 11608 6092 11620
rect 4120 11580 6092 11608
rect 4120 11568 4126 11580
rect 6086 11568 6092 11580
rect 6144 11568 6150 11620
rect 6380 11540 6408 11648
rect 6546 11608 6552 11620
rect 6507 11580 6552 11608
rect 6546 11568 6552 11580
rect 6604 11568 6610 11620
rect 6656 11608 6684 11716
rect 6733 11713 6745 11747
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 11698 11704 11704 11756
rect 11756 11744 11762 11756
rect 12066 11744 12072 11756
rect 11756 11716 12072 11744
rect 11756 11704 11762 11716
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 12158 11704 12164 11756
rect 12216 11744 12222 11756
rect 14292 11744 14320 11784
rect 18230 11772 18236 11784
rect 18288 11772 18294 11824
rect 18598 11772 18604 11824
rect 18656 11772 18662 11824
rect 23768 11812 23796 11852
rect 19444 11784 23796 11812
rect 23845 11815 23903 11821
rect 12216 11716 14320 11744
rect 14369 11747 14427 11753
rect 12216 11704 12222 11716
rect 14369 11713 14381 11747
rect 14415 11744 14427 11747
rect 15197 11747 15255 11753
rect 14415 11716 14872 11744
rect 14415 11713 14427 11716
rect 14369 11707 14427 11713
rect 7469 11679 7527 11685
rect 7469 11645 7481 11679
rect 7515 11676 7527 11679
rect 8478 11676 8484 11688
rect 7515 11648 8484 11676
rect 7515 11645 7527 11648
rect 7469 11639 7527 11645
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 8938 11676 8944 11688
rect 8899 11648 8944 11676
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 10226 11676 10232 11688
rect 9048 11648 10232 11676
rect 9048 11608 9076 11648
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 10502 11636 10508 11688
rect 10560 11676 10566 11688
rect 10689 11679 10747 11685
rect 10689 11676 10701 11679
rect 10560 11648 10701 11676
rect 10560 11636 10566 11648
rect 10689 11645 10701 11648
rect 10735 11645 10747 11679
rect 10689 11639 10747 11645
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 11609 11611 11667 11617
rect 11609 11608 11621 11611
rect 6656 11580 9076 11608
rect 10244 11580 11621 11608
rect 7282 11540 7288 11552
rect 6380 11512 7288 11540
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 8018 11540 8024 11552
rect 7979 11512 8024 11540
rect 8018 11500 8024 11512
rect 8076 11500 8082 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 10244 11540 10272 11580
rect 11609 11577 11621 11580
rect 11655 11577 11667 11611
rect 11609 11571 11667 11577
rect 11698 11568 11704 11620
rect 11756 11608 11762 11620
rect 12268 11608 12296 11639
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 12400 11648 12817 11676
rect 12400 11636 12406 11648
rect 12805 11645 12817 11648
rect 12851 11645 12863 11679
rect 12805 11639 12863 11645
rect 13446 11608 13452 11620
rect 11756 11580 13452 11608
rect 11756 11568 11762 11580
rect 13446 11568 13452 11580
rect 13504 11568 13510 11620
rect 14844 11617 14872 11716
rect 15197 11713 15209 11747
rect 15243 11744 15255 11747
rect 15930 11744 15936 11756
rect 15243 11716 15936 11744
rect 15243 11713 15255 11716
rect 15197 11707 15255 11713
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 17218 11744 17224 11756
rect 17179 11716 17224 11744
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 15289 11679 15347 11685
rect 15289 11645 15301 11679
rect 15335 11645 15347 11679
rect 15470 11676 15476 11688
rect 15431 11648 15476 11676
rect 15289 11639 15347 11645
rect 14829 11611 14887 11617
rect 14829 11577 14841 11611
rect 14875 11577 14887 11611
rect 14829 11571 14887 11577
rect 15194 11568 15200 11620
rect 15252 11608 15258 11620
rect 15304 11608 15332 11639
rect 15470 11636 15476 11648
rect 15528 11636 15534 11688
rect 15746 11636 15752 11688
rect 15804 11676 15810 11688
rect 16666 11676 16672 11688
rect 15804 11648 16672 11676
rect 15804 11636 15810 11648
rect 16666 11636 16672 11648
rect 16724 11676 16730 11688
rect 17862 11676 17868 11688
rect 16724 11648 17868 11676
rect 16724 11636 16730 11648
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 18138 11676 18144 11688
rect 18099 11648 18144 11676
rect 18138 11636 18144 11648
rect 18196 11636 18202 11688
rect 18230 11636 18236 11688
rect 18288 11676 18294 11688
rect 19444 11676 19472 11784
rect 23845 11781 23857 11815
rect 23891 11781 23903 11815
rect 23845 11775 23903 11781
rect 20346 11744 20352 11756
rect 20307 11716 20352 11744
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 21085 11747 21143 11753
rect 21085 11744 21097 11747
rect 20456 11716 21097 11744
rect 18288 11648 19472 11676
rect 18288 11636 18294 11648
rect 20070 11636 20076 11688
rect 20128 11676 20134 11688
rect 20456 11676 20484 11716
rect 21085 11713 21097 11716
rect 21131 11713 21143 11747
rect 21821 11747 21879 11753
rect 21821 11744 21833 11747
rect 21085 11707 21143 11713
rect 21192 11716 21833 11744
rect 20128 11648 20484 11676
rect 20128 11636 20134 11648
rect 20990 11636 20996 11688
rect 21048 11676 21054 11688
rect 21192 11676 21220 11716
rect 21821 11713 21833 11716
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 22002 11704 22008 11756
rect 22060 11744 22066 11756
rect 22557 11747 22615 11753
rect 22557 11744 22569 11747
rect 22060 11716 22569 11744
rect 22060 11704 22066 11716
rect 22557 11713 22569 11716
rect 22603 11713 22615 11747
rect 22557 11707 22615 11713
rect 23201 11747 23259 11753
rect 23201 11713 23213 11747
rect 23247 11713 23259 11747
rect 23201 11707 23259 11713
rect 23385 11747 23443 11753
rect 23385 11713 23397 11747
rect 23431 11744 23443 11747
rect 23474 11744 23480 11756
rect 23431 11716 23480 11744
rect 23431 11713 23443 11716
rect 23385 11707 23443 11713
rect 21048 11648 21220 11676
rect 23216 11676 23244 11707
rect 23474 11704 23480 11716
rect 23532 11704 23538 11756
rect 23860 11744 23888 11775
rect 23934 11772 23940 11824
rect 23992 11812 23998 11824
rect 24061 11815 24119 11821
rect 24061 11812 24073 11815
rect 23992 11784 24073 11812
rect 23992 11772 23998 11784
rect 24061 11781 24073 11784
rect 24107 11812 24119 11815
rect 24210 11812 24216 11824
rect 24107 11784 24216 11812
rect 24107 11781 24119 11784
rect 24061 11775 24119 11781
rect 24210 11772 24216 11784
rect 24268 11772 24274 11824
rect 26252 11812 26280 11852
rect 26326 11840 26332 11892
rect 26384 11880 26390 11892
rect 26786 11880 26792 11892
rect 26384 11852 26792 11880
rect 26384 11840 26390 11852
rect 26786 11840 26792 11852
rect 26844 11840 26850 11892
rect 26973 11883 27031 11889
rect 26973 11849 26985 11883
rect 27019 11880 27031 11883
rect 27246 11880 27252 11892
rect 27019 11852 27252 11880
rect 27019 11849 27031 11852
rect 26973 11843 27031 11849
rect 27246 11840 27252 11852
rect 27304 11840 27310 11892
rect 27982 11840 27988 11892
rect 28040 11880 28046 11892
rect 28353 11883 28411 11889
rect 28353 11880 28365 11883
rect 28040 11852 28365 11880
rect 28040 11840 28046 11852
rect 28353 11849 28365 11852
rect 28399 11849 28411 11883
rect 28353 11843 28411 11849
rect 28626 11840 28632 11892
rect 28684 11880 28690 11892
rect 29914 11880 29920 11892
rect 28684 11852 29684 11880
rect 29875 11852 29920 11880
rect 28684 11840 28690 11852
rect 29454 11812 29460 11824
rect 26252 11784 29460 11812
rect 29454 11772 29460 11784
rect 29512 11772 29518 11824
rect 29656 11821 29684 11852
rect 29914 11840 29920 11852
rect 29972 11840 29978 11892
rect 30650 11880 30656 11892
rect 30611 11852 30656 11880
rect 30650 11840 30656 11852
rect 30708 11840 30714 11892
rect 33226 11880 33232 11892
rect 33187 11852 33232 11880
rect 33226 11840 33232 11852
rect 33284 11840 33290 11892
rect 33502 11840 33508 11892
rect 33560 11880 33566 11892
rect 33965 11883 34023 11889
rect 33965 11880 33977 11883
rect 33560 11852 33977 11880
rect 33560 11840 33566 11852
rect 33965 11849 33977 11852
rect 34011 11849 34023 11883
rect 34698 11880 34704 11892
rect 34611 11852 34704 11880
rect 33965 11843 34023 11849
rect 34698 11840 34704 11852
rect 34756 11880 34762 11892
rect 37277 11883 37335 11889
rect 34756 11852 36768 11880
rect 34756 11840 34762 11852
rect 29641 11815 29699 11821
rect 29641 11781 29653 11815
rect 29687 11781 29699 11815
rect 29641 11775 29699 11781
rect 36740 11812 36768 11852
rect 37277 11849 37289 11883
rect 37323 11880 37335 11883
rect 37550 11880 37556 11892
rect 37323 11852 37556 11880
rect 37323 11849 37335 11852
rect 37277 11843 37335 11849
rect 37550 11840 37556 11852
rect 37608 11840 37614 11892
rect 38295 11883 38353 11889
rect 38295 11849 38307 11883
rect 38341 11880 38353 11883
rect 39022 11880 39028 11892
rect 38341 11852 39028 11880
rect 38341 11849 38353 11852
rect 38295 11843 38353 11849
rect 39022 11840 39028 11852
rect 39080 11840 39086 11892
rect 39942 11840 39948 11892
rect 40000 11880 40006 11892
rect 41598 11880 41604 11892
rect 40000 11852 41604 11880
rect 40000 11840 40006 11852
rect 41598 11840 41604 11852
rect 41656 11840 41662 11892
rect 36740 11784 37587 11812
rect 24486 11744 24492 11756
rect 23860 11716 24492 11744
rect 24486 11704 24492 11716
rect 24544 11704 24550 11756
rect 24670 11744 24676 11756
rect 24631 11716 24676 11744
rect 24670 11704 24676 11716
rect 24728 11704 24734 11756
rect 26082 11716 26648 11744
rect 23934 11676 23940 11688
rect 23216 11648 23940 11676
rect 21048 11636 21054 11648
rect 23934 11636 23940 11648
rect 23992 11636 23998 11688
rect 24213 11611 24271 11617
rect 24213 11608 24225 11611
rect 15252 11580 15332 11608
rect 19352 11580 24225 11608
rect 15252 11568 15258 11580
rect 8444 11512 10272 11540
rect 8444 11500 8450 11512
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 12710 11540 12716 11552
rect 12124 11512 12716 11540
rect 12124 11500 12130 11512
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 14090 11500 14096 11552
rect 14148 11540 14154 11552
rect 14185 11543 14243 11549
rect 14185 11540 14197 11543
rect 14148 11512 14197 11540
rect 14148 11500 14154 11512
rect 14185 11509 14197 11512
rect 14231 11509 14243 11543
rect 14185 11503 14243 11509
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 19352 11540 19380 11580
rect 24213 11577 24225 11580
rect 24259 11577 24271 11611
rect 24504 11608 24532 11704
rect 24949 11679 25007 11685
rect 24949 11645 24961 11679
rect 24995 11676 25007 11679
rect 26142 11676 26148 11688
rect 24995 11648 26148 11676
rect 24995 11645 25007 11648
rect 24949 11639 25007 11645
rect 26142 11636 26148 11648
rect 26200 11636 26206 11688
rect 26418 11676 26424 11688
rect 26379 11648 26424 11676
rect 26418 11636 26424 11648
rect 26476 11636 26482 11688
rect 26620 11676 26648 11716
rect 26694 11704 26700 11756
rect 26752 11744 26758 11756
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 26752 11716 27169 11744
rect 26752 11704 26758 11716
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 27246 11704 27252 11756
rect 27304 11744 27310 11756
rect 27614 11744 27620 11756
rect 27304 11716 27620 11744
rect 27304 11704 27310 11716
rect 27614 11704 27620 11716
rect 27672 11704 27678 11756
rect 28261 11747 28319 11753
rect 28261 11713 28273 11747
rect 28307 11744 28319 11747
rect 28810 11744 28816 11756
rect 28307 11716 28816 11744
rect 28307 11713 28319 11716
rect 28261 11707 28319 11713
rect 28810 11704 28816 11716
rect 28868 11704 28874 11756
rect 29365 11747 29423 11753
rect 29365 11713 29377 11747
rect 29411 11713 29423 11747
rect 29549 11747 29607 11753
rect 29549 11744 29561 11747
rect 29365 11707 29423 11713
rect 29472 11716 29561 11744
rect 27709 11679 27767 11685
rect 27709 11676 27721 11679
rect 26620 11648 27721 11676
rect 27709 11645 27721 11648
rect 27755 11645 27767 11679
rect 27709 11639 27767 11645
rect 24504 11580 24808 11608
rect 24213 11571 24271 11577
rect 16724 11512 19380 11540
rect 16724 11500 16730 11512
rect 20070 11500 20076 11552
rect 20128 11540 20134 11552
rect 22002 11540 22008 11552
rect 20128 11512 22008 11540
rect 20128 11500 20134 11512
rect 22002 11500 22008 11512
rect 22060 11500 22066 11552
rect 23290 11540 23296 11552
rect 23251 11512 23296 11540
rect 23290 11500 23296 11512
rect 23348 11500 23354 11552
rect 23474 11500 23480 11552
rect 23532 11540 23538 11552
rect 24029 11543 24087 11549
rect 24029 11540 24041 11543
rect 23532 11512 24041 11540
rect 23532 11500 23538 11512
rect 24029 11509 24041 11512
rect 24075 11540 24087 11543
rect 24578 11540 24584 11552
rect 24075 11512 24584 11540
rect 24075 11509 24087 11512
rect 24029 11503 24087 11509
rect 24578 11500 24584 11512
rect 24636 11500 24642 11552
rect 24780 11540 24808 11580
rect 25958 11568 25964 11620
rect 26016 11608 26022 11620
rect 27338 11608 27344 11620
rect 26016 11580 27344 11608
rect 26016 11568 26022 11580
rect 27338 11568 27344 11580
rect 27396 11568 27402 11620
rect 29380 11608 29408 11707
rect 29472 11676 29500 11716
rect 29549 11713 29561 11716
rect 29595 11713 29607 11747
rect 29549 11707 29607 11713
rect 29730 11704 29736 11756
rect 29788 11744 29794 11756
rect 30929 11747 30987 11753
rect 30929 11744 30941 11747
rect 29788 11716 29833 11744
rect 29923 11716 30941 11744
rect 29788 11704 29794 11716
rect 29923 11676 29951 11716
rect 30929 11713 30941 11716
rect 30975 11744 30987 11747
rect 32585 11747 32643 11753
rect 30975 11716 32536 11744
rect 30975 11713 30987 11716
rect 30929 11707 30987 11713
rect 30834 11676 30840 11688
rect 29472 11648 29951 11676
rect 30795 11648 30840 11676
rect 30834 11636 30840 11648
rect 30892 11636 30898 11688
rect 31202 11676 31208 11688
rect 30944 11648 31208 11676
rect 30650 11608 30656 11620
rect 29380 11580 30656 11608
rect 30650 11568 30656 11580
rect 30708 11568 30714 11620
rect 30944 11540 30972 11648
rect 31202 11636 31208 11648
rect 31260 11636 31266 11688
rect 31294 11636 31300 11688
rect 31352 11676 31358 11688
rect 32508 11676 32536 11716
rect 32585 11713 32597 11747
rect 32631 11744 32643 11747
rect 33226 11744 33232 11756
rect 32631 11716 33232 11744
rect 32631 11713 32643 11716
rect 32585 11707 32643 11713
rect 33226 11704 33232 11716
rect 33284 11704 33290 11756
rect 33410 11744 33416 11756
rect 33371 11716 33416 11744
rect 33410 11704 33416 11716
rect 33468 11704 33474 11756
rect 33873 11747 33931 11753
rect 33873 11713 33885 11747
rect 33919 11744 33931 11747
rect 34146 11744 34152 11756
rect 33919 11716 34152 11744
rect 33919 11713 33931 11716
rect 33873 11707 33931 11713
rect 32766 11676 32772 11688
rect 31352 11648 31397 11676
rect 32508 11648 32772 11676
rect 31352 11636 31358 11648
rect 32766 11636 32772 11648
rect 32824 11636 32830 11688
rect 33134 11636 33140 11688
rect 33192 11676 33198 11688
rect 33888 11676 33916 11707
rect 34146 11704 34152 11716
rect 34204 11704 34210 11756
rect 34606 11744 34612 11756
rect 34567 11716 34612 11744
rect 34606 11704 34612 11716
rect 34664 11704 34670 11756
rect 36538 11744 36544 11756
rect 36499 11716 36544 11744
rect 36538 11704 36544 11716
rect 36596 11704 36602 11756
rect 36740 11753 36768 11784
rect 36725 11747 36783 11753
rect 36725 11713 36737 11747
rect 36771 11713 36783 11747
rect 36725 11707 36783 11713
rect 37461 11747 37519 11753
rect 37461 11713 37473 11747
rect 37507 11713 37519 11747
rect 37461 11707 37519 11713
rect 33192 11648 33916 11676
rect 36633 11679 36691 11685
rect 33192 11636 33198 11648
rect 36633 11645 36645 11679
rect 36679 11676 36691 11679
rect 37476 11676 37504 11707
rect 36679 11648 37504 11676
rect 37559 11676 37587 11784
rect 37642 11772 37648 11824
rect 37700 11812 37706 11824
rect 38562 11812 38568 11824
rect 37700 11784 38240 11812
rect 37700 11772 37706 11784
rect 37734 11744 37740 11756
rect 37695 11716 37740 11744
rect 37734 11704 37740 11716
rect 37792 11704 37798 11756
rect 38212 11753 38240 11784
rect 38396 11784 38568 11812
rect 38197 11747 38255 11753
rect 38197 11713 38209 11747
rect 38243 11744 38255 11747
rect 38286 11744 38292 11756
rect 38243 11716 38292 11744
rect 38243 11713 38255 11716
rect 38197 11707 38255 11713
rect 38286 11704 38292 11716
rect 38344 11704 38350 11756
rect 38396 11753 38424 11784
rect 38562 11772 38568 11784
rect 38620 11772 38626 11824
rect 39298 11772 39304 11824
rect 39356 11812 39362 11824
rect 40126 11812 40132 11824
rect 39356 11784 40132 11812
rect 39356 11772 39362 11784
rect 40126 11772 40132 11784
rect 40184 11772 40190 11824
rect 40221 11815 40279 11821
rect 40221 11781 40233 11815
rect 40267 11812 40279 11815
rect 40494 11812 40500 11824
rect 40267 11784 40500 11812
rect 40267 11781 40279 11784
rect 40221 11775 40279 11781
rect 40494 11772 40500 11784
rect 40552 11812 40558 11824
rect 41506 11812 41512 11824
rect 40552 11784 41512 11812
rect 40552 11772 40558 11784
rect 41506 11772 41512 11784
rect 41564 11772 41570 11824
rect 38381 11747 38439 11753
rect 38381 11713 38393 11747
rect 38427 11713 38439 11747
rect 38381 11707 38439 11713
rect 38470 11704 38476 11756
rect 38528 11744 38534 11756
rect 38930 11744 38936 11756
rect 38528 11716 38573 11744
rect 38891 11716 38936 11744
rect 38528 11704 38534 11716
rect 38930 11704 38936 11716
rect 38988 11704 38994 11756
rect 39022 11704 39028 11756
rect 39080 11744 39086 11756
rect 39209 11747 39267 11753
rect 39080 11716 39125 11744
rect 39080 11704 39086 11716
rect 39209 11713 39221 11747
rect 39255 11713 39267 11747
rect 39209 11707 39267 11713
rect 39398 11747 39456 11753
rect 39398 11713 39410 11747
rect 39444 11744 39456 11747
rect 39758 11744 39764 11756
rect 39444 11716 39764 11744
rect 39444 11713 39456 11716
rect 39398 11707 39456 11713
rect 38010 11676 38016 11688
rect 37559 11648 38016 11676
rect 36679 11645 36691 11648
rect 36633 11639 36691 11645
rect 38010 11636 38016 11648
rect 38068 11636 38074 11688
rect 38102 11636 38108 11688
rect 38160 11676 38166 11688
rect 39224 11676 39252 11707
rect 39758 11704 39764 11716
rect 39816 11704 39822 11756
rect 39942 11704 39948 11756
rect 40000 11744 40006 11756
rect 40313 11747 40371 11753
rect 40313 11744 40325 11747
rect 40000 11716 40325 11744
rect 40000 11704 40006 11716
rect 40313 11713 40325 11716
rect 40359 11713 40371 11747
rect 40313 11707 40371 11713
rect 40402 11704 40408 11756
rect 40460 11744 40466 11756
rect 40460 11716 40505 11744
rect 40460 11704 40466 11716
rect 40586 11704 40592 11756
rect 40644 11744 40650 11756
rect 40644 11716 40689 11744
rect 40644 11704 40650 11716
rect 40770 11704 40776 11756
rect 40828 11744 40834 11756
rect 41049 11747 41107 11753
rect 41049 11744 41061 11747
rect 40828 11716 41061 11744
rect 40828 11704 40834 11716
rect 41049 11713 41061 11716
rect 41095 11744 41107 11747
rect 41966 11744 41972 11756
rect 41095 11716 41972 11744
rect 41095 11713 41107 11716
rect 41049 11707 41107 11713
rect 41966 11704 41972 11716
rect 42024 11704 42030 11756
rect 42426 11676 42432 11688
rect 38160 11648 41184 11676
rect 42387 11648 42432 11676
rect 38160 11636 38166 11648
rect 40037 11611 40095 11617
rect 40037 11608 40049 11611
rect 39224 11580 40049 11608
rect 24780 11512 30972 11540
rect 31938 11500 31944 11552
rect 31996 11540 32002 11552
rect 32677 11543 32735 11549
rect 32677 11540 32689 11543
rect 31996 11512 32689 11540
rect 31996 11500 32002 11512
rect 32677 11509 32689 11512
rect 32723 11509 32735 11543
rect 32677 11503 32735 11509
rect 37274 11500 37280 11552
rect 37332 11540 37338 11552
rect 37550 11540 37556 11552
rect 37332 11512 37556 11540
rect 37332 11500 37338 11512
rect 37550 11500 37556 11512
rect 37608 11540 37614 11552
rect 37645 11543 37703 11549
rect 37645 11540 37657 11543
rect 37608 11512 37657 11540
rect 37608 11500 37614 11512
rect 37645 11509 37657 11512
rect 37691 11540 37703 11543
rect 38470 11540 38476 11552
rect 37691 11512 38476 11540
rect 37691 11509 37703 11512
rect 37645 11503 37703 11509
rect 38470 11500 38476 11512
rect 38528 11500 38534 11552
rect 39022 11500 39028 11552
rect 39080 11540 39086 11552
rect 39224 11540 39252 11580
rect 40037 11577 40049 11580
rect 40083 11608 40095 11611
rect 40310 11608 40316 11620
rect 40083 11580 40316 11608
rect 40083 11577 40095 11580
rect 40037 11571 40095 11577
rect 40310 11568 40316 11580
rect 40368 11568 40374 11620
rect 39080 11512 39252 11540
rect 39577 11543 39635 11549
rect 39080 11500 39086 11512
rect 39577 11509 39589 11543
rect 39623 11540 39635 11543
rect 40494 11540 40500 11552
rect 39623 11512 40500 11540
rect 39623 11509 39635 11512
rect 39577 11503 39635 11509
rect 40494 11500 40500 11512
rect 40552 11500 40558 11552
rect 41156 11549 41184 11648
rect 42426 11636 42432 11648
rect 42484 11636 42490 11688
rect 42702 11676 42708 11688
rect 42663 11648 42708 11676
rect 42702 11636 42708 11648
rect 42760 11636 42766 11688
rect 41141 11543 41199 11549
rect 41141 11509 41153 11543
rect 41187 11509 41199 11543
rect 41141 11503 41199 11509
rect 41322 11500 41328 11552
rect 41380 11540 41386 11552
rect 41509 11543 41567 11549
rect 41509 11540 41521 11543
rect 41380 11512 41521 11540
rect 41380 11500 41386 11512
rect 41509 11509 41521 11512
rect 41555 11509 41567 11543
rect 41509 11503 41567 11509
rect 1104 11450 44896 11472
rect 1104 11398 6424 11450
rect 6476 11398 6488 11450
rect 6540 11398 6552 11450
rect 6604 11398 6616 11450
rect 6668 11398 6680 11450
rect 6732 11398 17372 11450
rect 17424 11398 17436 11450
rect 17488 11398 17500 11450
rect 17552 11398 17564 11450
rect 17616 11398 17628 11450
rect 17680 11398 28320 11450
rect 28372 11398 28384 11450
rect 28436 11398 28448 11450
rect 28500 11398 28512 11450
rect 28564 11398 28576 11450
rect 28628 11398 39268 11450
rect 39320 11398 39332 11450
rect 39384 11398 39396 11450
rect 39448 11398 39460 11450
rect 39512 11398 39524 11450
rect 39576 11398 44896 11450
rect 1104 11376 44896 11398
rect 2501 11339 2559 11345
rect 2501 11305 2513 11339
rect 2547 11336 2559 11339
rect 2682 11336 2688 11348
rect 2547 11308 2688 11336
rect 2547 11305 2559 11308
rect 2501 11299 2559 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 8202 11336 8208 11348
rect 4212 11308 7420 11336
rect 8163 11308 8208 11336
rect 4212 11296 4218 11308
rect 2958 11200 2964 11212
rect 2919 11172 2964 11200
rect 2958 11160 2964 11172
rect 3016 11160 3022 11212
rect 3145 11203 3203 11209
rect 3145 11169 3157 11203
rect 3191 11200 3203 11203
rect 4246 11200 4252 11212
rect 3191 11172 4252 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 7392 11200 7420 11308
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 10318 11336 10324 11348
rect 8904 11308 9904 11336
rect 10279 11308 10324 11336
rect 8904 11296 8910 11308
rect 7745 11271 7803 11277
rect 7745 11237 7757 11271
rect 7791 11268 7803 11271
rect 8478 11268 8484 11280
rect 7791 11240 8484 11268
rect 7791 11237 7803 11240
rect 7745 11231 7803 11237
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 9876 11268 9904 11308
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 12618 11336 12624 11348
rect 10468 11308 12624 11336
rect 10468 11296 10474 11308
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 12805 11339 12863 11345
rect 12805 11305 12817 11339
rect 12851 11336 12863 11339
rect 12986 11336 12992 11348
rect 12851 11308 12992 11336
rect 12851 11305 12863 11308
rect 12805 11299 12863 11305
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 15930 11336 15936 11348
rect 13740 11308 15516 11336
rect 15891 11308 15936 11336
rect 10781 11271 10839 11277
rect 10781 11268 10793 11271
rect 9876 11240 10793 11268
rect 10781 11237 10793 11240
rect 10827 11237 10839 11271
rect 12158 11268 12164 11280
rect 10781 11231 10839 11237
rect 10888 11240 12164 11268
rect 10888 11200 10916 11240
rect 12158 11228 12164 11240
rect 12216 11228 12222 11280
rect 12345 11271 12403 11277
rect 12345 11237 12357 11271
rect 12391 11268 12403 11271
rect 12434 11268 12440 11280
rect 12391 11240 12440 11268
rect 12391 11237 12403 11240
rect 12345 11231 12403 11237
rect 12434 11228 12440 11240
rect 12492 11268 12498 11280
rect 13740 11268 13768 11308
rect 12492 11240 13768 11268
rect 15488 11268 15516 11308
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 17865 11339 17923 11345
rect 17865 11305 17877 11339
rect 17911 11336 17923 11339
rect 18138 11336 18144 11348
rect 17911 11308 18144 11336
rect 17911 11305 17923 11308
rect 17865 11299 17923 11305
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 18598 11336 18604 11348
rect 18559 11308 18604 11336
rect 18598 11296 18604 11308
rect 18656 11296 18662 11348
rect 20070 11336 20076 11348
rect 19352 11308 20076 11336
rect 16574 11268 16580 11280
rect 15488 11240 16580 11268
rect 12492 11228 12498 11240
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 16850 11228 16856 11280
rect 16908 11268 16914 11280
rect 19352 11268 19380 11308
rect 20070 11296 20076 11308
rect 20128 11296 20134 11348
rect 20346 11296 20352 11348
rect 20404 11336 20410 11348
rect 20717 11339 20775 11345
rect 20717 11336 20729 11339
rect 20404 11308 20729 11336
rect 20404 11296 20410 11308
rect 20717 11305 20729 11308
rect 20763 11305 20775 11339
rect 20717 11299 20775 11305
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 25958 11336 25964 11348
rect 23256 11308 25964 11336
rect 23256 11296 23262 11308
rect 25958 11296 25964 11308
rect 26016 11296 26022 11348
rect 26142 11336 26148 11348
rect 26103 11308 26148 11336
rect 26142 11296 26148 11308
rect 26200 11296 26206 11348
rect 30650 11336 30656 11348
rect 26252 11308 30512 11336
rect 30611 11308 30656 11336
rect 26252 11268 26280 11308
rect 27249 11271 27307 11277
rect 27249 11268 27261 11271
rect 16908 11240 19380 11268
rect 20364 11240 26280 11268
rect 26344 11240 27261 11268
rect 16908 11228 16914 11240
rect 7392 11172 9076 11200
rect 3694 11092 3700 11144
rect 3752 11132 3758 11144
rect 4614 11141 4620 11144
rect 4341 11135 4399 11141
rect 4341 11132 4353 11135
rect 3752 11104 4353 11132
rect 3752 11092 3758 11104
rect 4341 11101 4353 11104
rect 4387 11101 4399 11135
rect 4608 11132 4620 11141
rect 4575 11104 4620 11132
rect 4341 11095 4399 11101
rect 4608 11095 4620 11104
rect 4614 11092 4620 11095
rect 4672 11092 4678 11144
rect 6365 11135 6423 11141
rect 6365 11101 6377 11135
rect 6411 11132 6423 11135
rect 8294 11132 8300 11144
rect 6411 11104 8300 11132
rect 6411 11101 6423 11104
rect 6365 11095 6423 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 8938 11132 8944 11144
rect 8444 11104 8489 11132
rect 8899 11104 8944 11132
rect 8444 11092 8450 11104
rect 8938 11092 8944 11104
rect 8996 11092 9002 11144
rect 9048 11132 9076 11172
rect 9968 11172 10916 11200
rect 11425 11203 11483 11209
rect 9968 11132 9996 11172
rect 11425 11169 11437 11203
rect 11471 11200 11483 11203
rect 11698 11200 11704 11212
rect 11471 11172 11704 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 13446 11200 13452 11212
rect 13407 11172 13452 11200
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 14182 11200 14188 11212
rect 14095 11172 14188 11200
rect 14182 11160 14188 11172
rect 14240 11200 14246 11212
rect 15746 11200 15752 11212
rect 14240 11172 15752 11200
rect 14240 11160 14246 11172
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 17862 11160 17868 11212
rect 17920 11200 17926 11212
rect 17920 11172 19380 11200
rect 17920 11160 17926 11172
rect 9048 11104 9996 11132
rect 10502 11092 10508 11144
rect 10560 11132 10566 11144
rect 11149 11135 11207 11141
rect 11149 11132 11161 11135
rect 10560 11104 11161 11132
rect 10560 11092 10566 11104
rect 11149 11101 11161 11104
rect 11195 11101 11207 11135
rect 11149 11095 11207 11101
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12250 11132 12256 11144
rect 12207 11104 12256 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 12526 11092 12532 11144
rect 12584 11132 12590 11144
rect 13265 11135 13323 11141
rect 13265 11132 13277 11135
rect 12584 11104 13277 11132
rect 12584 11092 12590 11104
rect 13265 11101 13277 11104
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 14090 11092 14096 11144
rect 14148 11132 14154 11144
rect 16666 11132 16672 11144
rect 14148 11104 14228 11132
rect 16627 11104 16672 11132
rect 14148 11092 14154 11104
rect 2869 11067 2927 11073
rect 2869 11033 2881 11067
rect 2915 11064 2927 11067
rect 5166 11064 5172 11076
rect 2915 11036 5172 11064
rect 2915 11033 2927 11036
rect 2869 11027 2927 11033
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 6632 11067 6690 11073
rect 6632 11064 6644 11067
rect 5736 11036 6644 11064
rect 5736 11005 5764 11036
rect 6632 11033 6644 11036
rect 6678 11064 6690 11067
rect 6822 11064 6828 11076
rect 6678 11036 6828 11064
rect 6678 11033 6690 11036
rect 6632 11027 6690 11033
rect 6822 11024 6828 11036
rect 6880 11024 6886 11076
rect 9030 11024 9036 11076
rect 9088 11064 9094 11076
rect 9186 11067 9244 11073
rect 9186 11064 9198 11067
rect 9088 11036 9198 11064
rect 9088 11024 9094 11036
rect 9186 11033 9198 11036
rect 9232 11033 9244 11067
rect 9186 11027 9244 11033
rect 9582 11024 9588 11076
rect 9640 11064 9646 11076
rect 10410 11064 10416 11076
rect 9640 11036 10416 11064
rect 9640 11024 9646 11036
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 11238 11064 11244 11076
rect 11199 11036 11244 11064
rect 11238 11024 11244 11036
rect 11296 11024 11302 11076
rect 13173 11067 13231 11073
rect 13173 11033 13185 11067
rect 13219 11064 13231 11067
rect 13998 11064 14004 11076
rect 13219 11036 14004 11064
rect 13219 11033 13231 11036
rect 13173 11027 13231 11033
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 14200 11064 14228 11104
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 18046 11132 18052 11144
rect 18007 11104 18052 11132
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18506 11132 18512 11144
rect 18467 11104 18512 11132
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 19352 11141 19380 11172
rect 19337 11135 19395 11141
rect 19337 11101 19349 11135
rect 19383 11132 19395 11135
rect 19886 11132 19892 11144
rect 19383 11104 19892 11132
rect 19383 11101 19395 11104
rect 19337 11095 19395 11101
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 14461 11067 14519 11073
rect 14461 11064 14473 11067
rect 14200 11036 14473 11064
rect 14461 11033 14473 11036
rect 14507 11033 14519 11067
rect 14461 11027 14519 11033
rect 15470 11024 15476 11076
rect 15528 11024 15534 11076
rect 18322 11024 18328 11076
rect 18380 11064 18386 11076
rect 19604 11067 19662 11073
rect 18380 11036 19564 11064
rect 18380 11024 18386 11036
rect 5721 10999 5779 11005
rect 5721 10965 5733 10999
rect 5767 10965 5779 10999
rect 5721 10959 5779 10965
rect 10226 10956 10232 11008
rect 10284 10996 10290 11008
rect 12434 10996 12440 11008
rect 10284 10968 12440 10996
rect 10284 10956 10290 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 15838 10996 15844 11008
rect 12676 10968 15844 10996
rect 12676 10956 12682 10968
rect 15838 10956 15844 10968
rect 15896 10956 15902 11008
rect 16022 10956 16028 11008
rect 16080 10996 16086 11008
rect 16485 10999 16543 11005
rect 16485 10996 16497 10999
rect 16080 10968 16497 10996
rect 16080 10956 16086 10968
rect 16485 10965 16497 10968
rect 16531 10965 16543 10999
rect 16485 10959 16543 10965
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 19334 10996 19340 11008
rect 16632 10968 19340 10996
rect 16632 10956 16638 10968
rect 19334 10956 19340 10968
rect 19392 10956 19398 11008
rect 19536 10996 19564 11036
rect 19604 11033 19616 11067
rect 19650 11064 19662 11067
rect 19702 11064 19708 11076
rect 19650 11036 19708 11064
rect 19650 11033 19662 11036
rect 19604 11027 19662 11033
rect 19702 11024 19708 11036
rect 19760 11024 19766 11076
rect 20364 11064 20392 11240
rect 20438 11160 20444 11212
rect 20496 11200 20502 11212
rect 20496 11172 20944 11200
rect 20496 11160 20502 11172
rect 19812 11036 20392 11064
rect 20916 11064 20944 11172
rect 22094 11160 22100 11212
rect 22152 11200 22158 11212
rect 22649 11203 22707 11209
rect 22649 11200 22661 11203
rect 22152 11172 22661 11200
rect 22152 11160 22158 11172
rect 22649 11169 22661 11172
rect 22695 11200 22707 11203
rect 23198 11200 23204 11212
rect 22695 11172 23204 11200
rect 22695 11169 22707 11172
rect 22649 11163 22707 11169
rect 23198 11160 23204 11172
rect 23256 11160 23262 11212
rect 23290 11160 23296 11212
rect 23348 11200 23354 11212
rect 26344 11209 26372 11240
rect 27249 11237 27261 11240
rect 27295 11237 27307 11271
rect 27249 11231 27307 11237
rect 27430 11228 27436 11280
rect 27488 11268 27494 11280
rect 29730 11268 29736 11280
rect 27488 11240 29736 11268
rect 27488 11228 27494 11240
rect 29730 11228 29736 11240
rect 29788 11228 29794 11280
rect 30006 11268 30012 11280
rect 29840 11240 30012 11268
rect 26329 11203 26387 11209
rect 23348 11172 25268 11200
rect 23348 11160 23354 11172
rect 22370 11092 22376 11144
rect 22428 11132 22434 11144
rect 22465 11135 22523 11141
rect 22465 11132 22477 11135
rect 22428 11104 22477 11132
rect 22428 11092 22434 11104
rect 22465 11101 22477 11104
rect 22511 11101 22523 11135
rect 22465 11095 22523 11101
rect 22557 11135 22615 11141
rect 22557 11101 22569 11135
rect 22603 11132 22615 11135
rect 23566 11132 23572 11144
rect 22603 11104 23572 11132
rect 22603 11101 22615 11104
rect 22557 11095 22615 11101
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 23845 11135 23903 11141
rect 23845 11101 23857 11135
rect 23891 11132 23903 11135
rect 24762 11132 24768 11144
rect 23891 11104 24768 11132
rect 23891 11101 23903 11104
rect 23845 11095 23903 11101
rect 24762 11092 24768 11104
rect 24820 11092 24826 11144
rect 24949 11135 25007 11141
rect 24949 11101 24961 11135
rect 24995 11132 25007 11135
rect 25130 11132 25136 11144
rect 24995 11104 25136 11132
rect 24995 11101 25007 11104
rect 24949 11095 25007 11101
rect 25130 11092 25136 11104
rect 25188 11092 25194 11144
rect 25240 11141 25268 11172
rect 26329 11169 26341 11203
rect 26375 11169 26387 11203
rect 26329 11163 26387 11169
rect 26510 11160 26516 11212
rect 26568 11200 26574 11212
rect 26697 11203 26755 11209
rect 26697 11200 26709 11203
rect 26568 11172 26709 11200
rect 26568 11160 26574 11172
rect 26697 11169 26709 11172
rect 26743 11169 26755 11203
rect 26697 11163 26755 11169
rect 25225 11135 25283 11141
rect 25225 11101 25237 11135
rect 25271 11132 25283 11135
rect 26421 11135 26479 11141
rect 25271 11104 26372 11132
rect 25271 11101 25283 11104
rect 25225 11095 25283 11101
rect 22278 11064 22284 11076
rect 20916 11036 22284 11064
rect 19812 10996 19840 11036
rect 22278 11024 22284 11036
rect 22336 11024 22342 11076
rect 26234 11064 26240 11076
rect 25240 11036 26240 11064
rect 25240 11008 25268 11036
rect 26234 11024 26240 11036
rect 26292 11024 26298 11076
rect 26344 11064 26372 11104
rect 26421 11101 26433 11135
rect 26467 11132 26479 11135
rect 26970 11132 26976 11144
rect 26467 11104 26976 11132
rect 26467 11101 26479 11104
rect 26421 11095 26479 11101
rect 26970 11092 26976 11104
rect 27028 11092 27034 11144
rect 27433 11135 27491 11141
rect 27433 11101 27445 11135
rect 27479 11132 27491 11135
rect 27614 11132 27620 11144
rect 27479 11104 27620 11132
rect 27479 11101 27491 11104
rect 27433 11095 27491 11101
rect 27614 11092 27620 11104
rect 27672 11092 27678 11144
rect 26789 11067 26847 11073
rect 26789 11064 26801 11067
rect 26344 11036 26801 11064
rect 26789 11033 26801 11036
rect 26835 11064 26847 11067
rect 29840 11064 29868 11240
rect 30006 11228 30012 11240
rect 30064 11228 30070 11280
rect 30006 11132 30012 11144
rect 29967 11104 30012 11132
rect 30006 11092 30012 11104
rect 30064 11092 30070 11144
rect 26835 11036 29868 11064
rect 30101 11067 30159 11073
rect 26835 11033 26847 11036
rect 26789 11027 26847 11033
rect 30101 11033 30113 11067
rect 30147 11064 30159 11067
rect 30374 11064 30380 11076
rect 30147 11036 30380 11064
rect 30147 11033 30159 11036
rect 30101 11027 30159 11033
rect 30374 11024 30380 11036
rect 30432 11024 30438 11076
rect 30484 11064 30512 11308
rect 30650 11296 30656 11308
rect 30708 11296 30714 11348
rect 31021 11339 31079 11345
rect 31021 11305 31033 11339
rect 31067 11336 31079 11339
rect 33410 11336 33416 11348
rect 31067 11308 33416 11336
rect 31067 11305 31079 11308
rect 31021 11299 31079 11305
rect 33410 11296 33416 11308
rect 33468 11296 33474 11348
rect 40586 11336 40592 11348
rect 36556 11308 40592 11336
rect 30668 11200 30696 11296
rect 30834 11228 30840 11280
rect 30892 11268 30898 11280
rect 31481 11271 31539 11277
rect 31481 11268 31493 11271
rect 30892 11240 31493 11268
rect 30892 11228 30898 11240
rect 31481 11237 31493 11240
rect 31527 11237 31539 11271
rect 31481 11231 31539 11237
rect 33686 11200 33692 11212
rect 30668 11172 31524 11200
rect 30650 11132 30656 11144
rect 30611 11104 30656 11132
rect 30650 11092 30656 11104
rect 30708 11092 30714 11144
rect 30742 11092 30748 11144
rect 30800 11132 30806 11144
rect 31496 11141 31524 11172
rect 32416 11172 33692 11200
rect 31481 11135 31539 11141
rect 30800 11104 30845 11132
rect 30800 11092 30806 11104
rect 31481 11101 31493 11135
rect 31527 11132 31539 11135
rect 31938 11132 31944 11144
rect 31527 11104 31944 11132
rect 31527 11101 31539 11104
rect 31481 11095 31539 11101
rect 31938 11092 31944 11104
rect 31996 11092 32002 11144
rect 32306 11132 32312 11144
rect 32267 11104 32312 11132
rect 32306 11092 32312 11104
rect 32364 11092 32370 11144
rect 32416 11064 32444 11172
rect 33686 11160 33692 11172
rect 33744 11160 33750 11212
rect 34103 11203 34161 11209
rect 34103 11169 34115 11203
rect 34149 11200 34161 11203
rect 34606 11200 34612 11212
rect 34149 11172 34612 11200
rect 34149 11169 34161 11172
rect 34103 11163 34161 11169
rect 34606 11160 34612 11172
rect 34664 11200 34670 11212
rect 34701 11203 34759 11209
rect 34701 11200 34713 11203
rect 34664 11172 34713 11200
rect 34664 11160 34670 11172
rect 34701 11169 34713 11172
rect 34747 11169 34759 11203
rect 34701 11163 34759 11169
rect 32582 11092 32588 11144
rect 32640 11132 32646 11144
rect 32677 11135 32735 11141
rect 32677 11132 32689 11135
rect 32640 11104 32689 11132
rect 32640 11092 32646 11104
rect 32677 11101 32689 11104
rect 32723 11101 32735 11135
rect 34974 11132 34980 11144
rect 34935 11104 34980 11132
rect 32677 11095 32735 11101
rect 34974 11092 34980 11104
rect 35032 11092 35038 11144
rect 36556 11141 36584 11308
rect 40586 11296 40592 11308
rect 40644 11296 40650 11348
rect 41046 11336 41052 11348
rect 41007 11308 41052 11336
rect 41046 11296 41052 11308
rect 41104 11296 41110 11348
rect 42058 11336 42064 11348
rect 42019 11308 42064 11336
rect 42058 11296 42064 11308
rect 42116 11296 42122 11348
rect 37185 11271 37243 11277
rect 37185 11237 37197 11271
rect 37231 11268 37243 11271
rect 37458 11268 37464 11280
rect 37231 11240 37464 11268
rect 37231 11237 37243 11240
rect 37185 11231 37243 11237
rect 37458 11228 37464 11240
rect 37516 11228 37522 11280
rect 39301 11271 39359 11277
rect 39301 11268 39313 11271
rect 39224 11240 39313 11268
rect 36998 11160 37004 11212
rect 37056 11200 37062 11212
rect 37918 11200 37924 11212
rect 37056 11172 37924 11200
rect 37056 11160 37062 11172
rect 37918 11160 37924 11172
rect 37976 11160 37982 11212
rect 36541 11135 36599 11141
rect 36541 11101 36553 11135
rect 36587 11101 36599 11135
rect 36541 11095 36599 11101
rect 36725 11135 36783 11141
rect 36725 11101 36737 11135
rect 36771 11132 36783 11135
rect 37461 11135 37519 11141
rect 36771 11104 37412 11132
rect 36771 11101 36783 11104
rect 36725 11095 36783 11101
rect 35618 11064 35624 11076
rect 30484 11036 32444 11064
rect 33718 11036 35624 11064
rect 35618 11024 35624 11036
rect 35676 11024 35682 11076
rect 37182 11064 37188 11076
rect 37143 11036 37188 11064
rect 37182 11024 37188 11036
rect 37240 11024 37246 11076
rect 37384 11073 37412 11104
rect 37461 11101 37473 11135
rect 37507 11134 37519 11135
rect 37550 11134 37556 11144
rect 37507 11106 37556 11134
rect 37507 11101 37519 11106
rect 37461 11095 37519 11101
rect 37550 11092 37556 11106
rect 37608 11092 37614 11144
rect 38562 11132 38568 11144
rect 37660 11104 38568 11132
rect 37369 11067 37427 11073
rect 37369 11033 37381 11067
rect 37415 11033 37427 11067
rect 37369 11027 37427 11033
rect 19536 10968 19840 10996
rect 19886 10956 19892 11008
rect 19944 10996 19950 11008
rect 20622 10996 20628 11008
rect 19944 10968 20628 10996
rect 19944 10956 19950 10968
rect 20622 10956 20628 10968
rect 20680 10956 20686 11008
rect 22097 10999 22155 11005
rect 22097 10965 22109 10999
rect 22143 10996 22155 10999
rect 22370 10996 22376 11008
rect 22143 10968 22376 10996
rect 22143 10965 22155 10968
rect 22097 10959 22155 10965
rect 22370 10956 22376 10968
rect 22428 10956 22434 11008
rect 23658 10996 23664 11008
rect 23619 10968 23664 10996
rect 23658 10956 23664 10968
rect 23716 10956 23722 11008
rect 24762 10996 24768 11008
rect 24723 10968 24768 10996
rect 24762 10956 24768 10968
rect 24820 10956 24826 11008
rect 25133 10999 25191 11005
rect 25133 10965 25145 10999
rect 25179 10996 25191 10999
rect 25222 10996 25228 11008
rect 25179 10968 25228 10996
rect 25179 10965 25191 10968
rect 25133 10959 25191 10965
rect 25222 10956 25228 10968
rect 25280 10956 25286 11008
rect 27246 10956 27252 11008
rect 27304 10996 27310 11008
rect 30190 10996 30196 11008
rect 27304 10968 30196 10996
rect 27304 10956 27310 10968
rect 30190 10956 30196 10968
rect 30248 10956 30254 11008
rect 36722 10996 36728 11008
rect 36683 10968 36728 10996
rect 36722 10956 36728 10968
rect 36780 10956 36786 11008
rect 37384 10996 37412 11027
rect 37660 10996 37688 11104
rect 38562 11092 38568 11104
rect 38620 11092 38626 11144
rect 38654 11092 38660 11144
rect 38712 11132 38718 11144
rect 39224 11132 39252 11240
rect 39301 11237 39313 11240
rect 39347 11268 39359 11271
rect 39942 11268 39948 11280
rect 39347 11240 39948 11268
rect 39347 11237 39359 11240
rect 39301 11231 39359 11237
rect 39942 11228 39948 11240
rect 40000 11228 40006 11280
rect 41322 11200 41328 11212
rect 39868 11172 41328 11200
rect 39868 11141 39896 11172
rect 41322 11160 41328 11172
rect 41380 11160 41386 11212
rect 41506 11160 41512 11212
rect 41564 11200 41570 11212
rect 42702 11200 42708 11212
rect 41564 11172 42708 11200
rect 41564 11160 41570 11172
rect 42702 11160 42708 11172
rect 42760 11160 42766 11212
rect 42812 11172 43668 11200
rect 38712 11104 39252 11132
rect 39853 11135 39911 11141
rect 38712 11092 38718 11104
rect 39853 11101 39865 11135
rect 39899 11101 39911 11135
rect 39853 11095 39911 11101
rect 40037 11135 40095 11141
rect 40037 11101 40049 11135
rect 40083 11101 40095 11135
rect 40037 11095 40095 11101
rect 40129 11135 40187 11141
rect 40129 11101 40141 11135
rect 40175 11101 40187 11135
rect 40129 11095 40187 11101
rect 37734 11024 37740 11076
rect 37792 11064 37798 11076
rect 38166 11067 38224 11073
rect 38166 11064 38178 11067
rect 37792 11036 38178 11064
rect 37792 11024 37798 11036
rect 38166 11033 38178 11036
rect 38212 11033 38224 11067
rect 39758 11064 39764 11076
rect 38166 11027 38224 11033
rect 38580 11036 39764 11064
rect 37384 10968 37688 10996
rect 37826 10956 37832 11008
rect 37884 10996 37890 11008
rect 38580 10996 38608 11036
rect 39758 11024 39764 11036
rect 39816 11064 39822 11076
rect 40052 11064 40080 11095
rect 39816 11036 40080 11064
rect 39816 11024 39822 11036
rect 40144 11008 40172 11095
rect 40218 11092 40224 11144
rect 40276 11132 40282 11144
rect 40276 11104 40321 11132
rect 40276 11092 40282 11104
rect 40402 11092 40408 11144
rect 40460 11132 40466 11144
rect 40460 11104 40505 11132
rect 40460 11092 40466 11104
rect 40954 11092 40960 11144
rect 41012 11132 41018 11144
rect 41233 11135 41291 11141
rect 41233 11132 41245 11135
rect 41012 11104 41245 11132
rect 41012 11092 41018 11104
rect 41233 11101 41245 11104
rect 41279 11101 41291 11135
rect 41414 11132 41420 11144
rect 41375 11104 41420 11132
rect 41233 11095 41291 11101
rect 41414 11092 41420 11104
rect 41472 11092 41478 11144
rect 41966 11132 41972 11144
rect 41927 11104 41972 11132
rect 41966 11092 41972 11104
rect 42024 11092 42030 11144
rect 42426 11092 42432 11144
rect 42484 11132 42490 11144
rect 42812 11141 42840 11172
rect 43640 11141 43668 11172
rect 42797 11135 42855 11141
rect 42797 11132 42809 11135
rect 42484 11104 42809 11132
rect 42484 11092 42490 11104
rect 42797 11101 42809 11104
rect 42843 11101 42855 11135
rect 42797 11095 42855 11101
rect 43441 11135 43499 11141
rect 43441 11101 43453 11135
rect 43487 11101 43499 11135
rect 43441 11095 43499 11101
rect 43625 11135 43683 11141
rect 43625 11101 43637 11135
rect 43671 11101 43683 11135
rect 43625 11095 43683 11101
rect 40236 11064 40264 11092
rect 41506 11064 41512 11076
rect 40236 11036 41512 11064
rect 41506 11024 41512 11036
rect 41564 11024 41570 11076
rect 42518 11024 42524 11076
rect 42576 11064 42582 11076
rect 42613 11067 42671 11073
rect 42613 11064 42625 11067
rect 42576 11036 42625 11064
rect 42576 11024 42582 11036
rect 42613 11033 42625 11036
rect 42659 11064 42671 11067
rect 43456 11064 43484 11095
rect 42659 11036 43484 11064
rect 42659 11033 42671 11036
rect 42613 11027 42671 11033
rect 37884 10968 38608 10996
rect 37884 10956 37890 10968
rect 40126 10956 40132 11008
rect 40184 10956 40190 11008
rect 40589 10999 40647 11005
rect 40589 10965 40601 10999
rect 40635 10996 40647 10999
rect 41046 10996 41052 11008
rect 40635 10968 41052 10996
rect 40635 10965 40647 10968
rect 40589 10959 40647 10965
rect 41046 10956 41052 10968
rect 41104 10956 41110 11008
rect 42886 10956 42892 11008
rect 42944 10996 42950 11008
rect 42981 10999 43039 11005
rect 42981 10996 42993 10999
rect 42944 10968 42993 10996
rect 42944 10956 42950 10968
rect 42981 10965 42993 10968
rect 43027 10965 43039 10999
rect 43530 10996 43536 11008
rect 43491 10968 43536 10996
rect 42981 10959 43039 10965
rect 43530 10956 43536 10968
rect 43588 10956 43594 11008
rect 1104 10906 45056 10928
rect 1104 10854 11898 10906
rect 11950 10854 11962 10906
rect 12014 10854 12026 10906
rect 12078 10854 12090 10906
rect 12142 10854 12154 10906
rect 12206 10854 22846 10906
rect 22898 10854 22910 10906
rect 22962 10854 22974 10906
rect 23026 10854 23038 10906
rect 23090 10854 23102 10906
rect 23154 10854 33794 10906
rect 33846 10854 33858 10906
rect 33910 10854 33922 10906
rect 33974 10854 33986 10906
rect 34038 10854 34050 10906
rect 34102 10854 44742 10906
rect 44794 10854 44806 10906
rect 44858 10854 44870 10906
rect 44922 10854 44934 10906
rect 44986 10854 44998 10906
rect 45050 10854 45056 10906
rect 1104 10832 45056 10854
rect 3237 10795 3295 10801
rect 3237 10761 3249 10795
rect 3283 10792 3295 10795
rect 3326 10792 3332 10804
rect 3283 10764 3332 10792
rect 3283 10761 3295 10764
rect 3237 10755 3295 10761
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 6270 10792 6276 10804
rect 3712 10764 6276 10792
rect 2774 10724 2780 10736
rect 1412 10696 2780 10724
rect 1412 10665 1440 10696
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 3712 10724 3740 10764
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 7101 10795 7159 10801
rect 7101 10761 7113 10795
rect 7147 10792 7159 10795
rect 8018 10792 8024 10804
rect 7147 10764 8024 10792
rect 7147 10761 7159 10764
rect 7101 10755 7159 10761
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 10594 10792 10600 10804
rect 10152 10764 10600 10792
rect 4430 10724 4436 10736
rect 2976 10696 3740 10724
rect 3804 10696 4436 10724
rect 1397 10659 1455 10665
rect 1397 10625 1409 10659
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 2409 10659 2467 10665
rect 2409 10625 2421 10659
rect 2455 10656 2467 10659
rect 2976 10656 3004 10696
rect 3804 10665 3832 10696
rect 4430 10684 4436 10696
rect 4488 10684 4494 10736
rect 7009 10727 7067 10733
rect 7009 10693 7021 10727
rect 7055 10724 7067 10727
rect 10152 10724 10180 10764
rect 10594 10752 10600 10764
rect 10652 10792 10658 10804
rect 14182 10792 14188 10804
rect 10652 10764 12020 10792
rect 10652 10752 10658 10764
rect 7055 10696 10180 10724
rect 7055 10693 7067 10696
rect 7009 10687 7067 10693
rect 10318 10684 10324 10736
rect 10376 10724 10382 10736
rect 10376 10696 10824 10724
rect 10376 10684 10382 10696
rect 2455 10628 3004 10656
rect 3053 10659 3111 10665
rect 2455 10625 2467 10628
rect 2409 10619 2467 10625
rect 3053 10625 3065 10659
rect 3099 10625 3111 10659
rect 3053 10619 3111 10625
rect 3789 10659 3847 10665
rect 3789 10625 3801 10659
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 2866 10588 2872 10600
rect 2827 10560 2872 10588
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 2222 10452 2228 10464
rect 2183 10424 2228 10452
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 3068 10452 3096 10619
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 4045 10659 4103 10665
rect 4045 10656 4057 10659
rect 3936 10628 4057 10656
rect 3936 10616 3942 10628
rect 4045 10625 4057 10628
rect 4091 10625 4103 10659
rect 4045 10619 4103 10625
rect 7837 10659 7895 10665
rect 7837 10625 7849 10659
rect 7883 10656 7895 10659
rect 10686 10656 10692 10668
rect 7883 10628 10692 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 10686 10616 10692 10628
rect 10744 10616 10750 10668
rect 10796 10665 10824 10696
rect 11992 10665 12020 10764
rect 13188 10764 14188 10792
rect 13188 10724 13216 10764
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 14274 10752 14280 10804
rect 14332 10792 14338 10804
rect 14826 10792 14832 10804
rect 14332 10764 14832 10792
rect 14332 10752 14338 10764
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 15381 10795 15439 10801
rect 15381 10761 15393 10795
rect 15427 10792 15439 10795
rect 15470 10792 15476 10804
rect 15427 10764 15476 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 22002 10792 22008 10804
rect 15896 10764 22008 10792
rect 15896 10752 15902 10764
rect 22002 10752 22008 10764
rect 22060 10752 22066 10804
rect 22189 10795 22247 10801
rect 22189 10761 22201 10795
rect 22235 10792 22247 10795
rect 22370 10792 22376 10804
rect 22235 10764 22376 10792
rect 22235 10761 22247 10764
rect 22189 10755 22247 10761
rect 22370 10752 22376 10764
rect 22428 10752 22434 10804
rect 26234 10792 26240 10804
rect 26195 10764 26240 10792
rect 26234 10752 26240 10764
rect 26292 10752 26298 10804
rect 32306 10752 32312 10804
rect 32364 10792 32370 10804
rect 35069 10795 35127 10801
rect 35069 10792 35081 10795
rect 32364 10764 35081 10792
rect 32364 10752 32370 10764
rect 35069 10761 35081 10764
rect 35115 10792 35127 10795
rect 36998 10792 37004 10804
rect 35115 10764 37004 10792
rect 35115 10761 35127 10764
rect 35069 10755 35127 10761
rect 36998 10752 37004 10764
rect 37056 10752 37062 10804
rect 39666 10792 39672 10804
rect 37568 10764 39672 10792
rect 13354 10724 13360 10736
rect 13096 10696 13216 10724
rect 13315 10696 13360 10724
rect 13096 10665 13124 10696
rect 13354 10684 13360 10696
rect 13412 10684 13418 10736
rect 15010 10724 15016 10736
rect 14582 10696 15016 10724
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 21910 10724 21916 10736
rect 16224 10696 21916 10724
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10625 13139 10659
rect 15286 10656 15292 10668
rect 15247 10628 15292 10656
rect 13081 10619 13139 10625
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 16117 10659 16175 10665
rect 16117 10625 16129 10659
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 7282 10588 7288 10600
rect 7195 10560 7288 10588
rect 7282 10548 7288 10560
rect 7340 10588 7346 10600
rect 9582 10588 9588 10600
rect 7340 10560 9588 10588
rect 7340 10548 7346 10560
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 10410 10548 10416 10600
rect 10468 10588 10474 10600
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 10468 10560 10609 10588
rect 10468 10548 10474 10560
rect 10597 10557 10609 10560
rect 10643 10588 10655 10591
rect 11793 10591 11851 10597
rect 11793 10588 11805 10591
rect 10643 10560 11805 10588
rect 10643 10557 10655 10560
rect 10597 10551 10655 10557
rect 11793 10557 11805 10560
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 12207 10560 14504 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 4982 10480 4988 10532
rect 5040 10520 5046 10532
rect 10226 10520 10232 10532
rect 5040 10492 10232 10520
rect 5040 10480 5046 10492
rect 10226 10480 10232 10492
rect 10284 10480 10290 10532
rect 10965 10523 11023 10529
rect 10965 10489 10977 10523
rect 11011 10520 11023 10523
rect 14476 10520 14504 10560
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 16132 10588 16160 10619
rect 14608 10560 16160 10588
rect 14608 10548 14614 10560
rect 16224 10520 16252 10696
rect 21910 10684 21916 10696
rect 21968 10684 21974 10736
rect 24670 10724 24676 10736
rect 24504 10696 24676 10724
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10625 17739 10659
rect 20990 10656 20996 10668
rect 20951 10628 20996 10656
rect 17681 10619 17739 10625
rect 17696 10588 17724 10619
rect 20990 10616 20996 10628
rect 21048 10616 21054 10668
rect 23014 10656 23020 10668
rect 22975 10628 23020 10656
rect 23014 10616 23020 10628
rect 23072 10616 23078 10668
rect 24504 10665 24532 10696
rect 24670 10684 24676 10696
rect 24728 10684 24734 10736
rect 24762 10684 24768 10736
rect 24820 10724 24826 10736
rect 24820 10696 24865 10724
rect 24820 10684 24826 10696
rect 25222 10684 25228 10736
rect 25280 10684 25286 10736
rect 33781 10727 33839 10733
rect 33781 10724 33793 10727
rect 28736 10696 33793 10724
rect 28736 10668 28764 10696
rect 33781 10693 33793 10696
rect 33827 10693 33839 10727
rect 33781 10687 33839 10693
rect 37369 10681 37427 10687
rect 24489 10659 24547 10665
rect 24489 10625 24501 10659
rect 24535 10625 24547 10659
rect 24489 10619 24547 10625
rect 28629 10659 28687 10665
rect 28629 10625 28641 10659
rect 28675 10656 28687 10659
rect 28718 10656 28724 10668
rect 28675 10628 28724 10656
rect 28675 10625 28687 10628
rect 28629 10619 28687 10625
rect 28718 10616 28724 10628
rect 28776 10616 28782 10668
rect 28810 10616 28816 10668
rect 28868 10656 28874 10668
rect 30837 10659 30895 10665
rect 30837 10656 30849 10659
rect 28868 10628 30849 10656
rect 28868 10616 28874 10628
rect 30837 10625 30849 10628
rect 30883 10625 30895 10659
rect 32582 10656 32588 10668
rect 32543 10628 32588 10656
rect 30837 10619 30895 10625
rect 32582 10616 32588 10628
rect 32640 10616 32646 10668
rect 32769 10659 32827 10665
rect 32769 10625 32781 10659
rect 32815 10625 32827 10659
rect 32769 10619 32827 10625
rect 32953 10659 33011 10665
rect 32953 10625 32965 10659
rect 32999 10625 33011 10659
rect 32953 10619 33011 10625
rect 33045 10659 33103 10665
rect 33045 10625 33057 10659
rect 33091 10656 33103 10659
rect 35802 10656 35808 10668
rect 33091 10628 35808 10656
rect 33091 10625 33103 10628
rect 33045 10619 33103 10625
rect 18506 10588 18512 10600
rect 17696 10560 18512 10588
rect 18506 10548 18512 10560
rect 18564 10588 18570 10600
rect 22278 10588 22284 10600
rect 18564 10560 21220 10588
rect 22239 10560 22284 10588
rect 18564 10548 18570 10560
rect 21192 10529 21220 10560
rect 22278 10548 22284 10560
rect 22336 10548 22342 10600
rect 22462 10588 22468 10600
rect 22423 10560 22468 10588
rect 22462 10548 22468 10560
rect 22520 10548 22526 10600
rect 30282 10588 30288 10600
rect 30243 10560 30288 10588
rect 30282 10548 30288 10560
rect 30340 10548 30346 10600
rect 32784 10588 32812 10619
rect 30392 10560 32812 10588
rect 32968 10588 32996 10619
rect 35802 10616 35808 10628
rect 35860 10616 35866 10668
rect 35986 10656 35992 10668
rect 35947 10628 35992 10656
rect 35986 10616 35992 10628
rect 36044 10616 36050 10668
rect 37369 10647 37381 10681
rect 37415 10678 37427 10681
rect 37415 10662 37504 10678
rect 37568 10662 37596 10764
rect 39666 10752 39672 10764
rect 39724 10792 39730 10804
rect 41414 10792 41420 10804
rect 39724 10764 41420 10792
rect 39724 10752 39730 10764
rect 41414 10752 41420 10764
rect 41472 10752 41478 10804
rect 38286 10724 38292 10736
rect 38247 10696 38292 10724
rect 38286 10684 38292 10696
rect 38344 10684 38350 10736
rect 42886 10724 42892 10736
rect 42847 10696 42892 10724
rect 42886 10684 42892 10696
rect 42944 10684 42950 10736
rect 37415 10650 37596 10662
rect 37415 10647 37427 10650
rect 37369 10641 37427 10647
rect 37476 10634 37596 10650
rect 38105 10659 38163 10665
rect 38105 10625 38117 10659
rect 38151 10625 38163 10659
rect 38105 10619 38163 10625
rect 38933 10659 38991 10665
rect 38933 10625 38945 10659
rect 38979 10656 38991 10659
rect 39114 10656 39120 10668
rect 38979 10628 39120 10656
rect 38979 10625 38991 10628
rect 38933 10619 38991 10625
rect 34974 10588 34980 10600
rect 32968 10560 34980 10588
rect 11011 10492 12434 10520
rect 14476 10492 16252 10520
rect 21177 10523 21235 10529
rect 11011 10489 11023 10492
rect 10965 10483 11023 10489
rect 5074 10452 5080 10464
rect 3068 10424 5080 10452
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 6641 10455 6699 10461
rect 5224 10424 5269 10452
rect 5224 10412 5230 10424
rect 6641 10421 6653 10455
rect 6687 10452 6699 10455
rect 8202 10452 8208 10464
rect 6687 10424 8208 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8938 10412 8944 10464
rect 8996 10452 9002 10464
rect 9214 10452 9220 10464
rect 8996 10424 9220 10452
rect 8996 10412 9002 10424
rect 9214 10412 9220 10424
rect 9272 10452 9278 10464
rect 9309 10455 9367 10461
rect 9309 10452 9321 10455
rect 9272 10424 9321 10452
rect 9272 10412 9278 10424
rect 9309 10421 9321 10424
rect 9355 10421 9367 10455
rect 12406 10452 12434 10492
rect 21177 10489 21189 10523
rect 21223 10520 21235 10523
rect 21726 10520 21732 10532
rect 21223 10492 21732 10520
rect 21223 10489 21235 10492
rect 21177 10483 21235 10489
rect 21726 10480 21732 10492
rect 21784 10480 21790 10532
rect 21910 10480 21916 10532
rect 21968 10520 21974 10532
rect 21968 10492 23336 10520
rect 21968 10480 21974 10492
rect 15470 10452 15476 10464
rect 12406 10424 15476 10452
rect 9309 10415 9367 10421
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 15562 10412 15568 10464
rect 15620 10452 15626 10464
rect 15933 10455 15991 10461
rect 15933 10452 15945 10455
rect 15620 10424 15945 10452
rect 15620 10412 15626 10424
rect 15933 10421 15945 10424
rect 15979 10421 15991 10455
rect 17770 10452 17776 10464
rect 17731 10424 17776 10452
rect 15933 10415 15991 10421
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 21821 10455 21879 10461
rect 21821 10421 21833 10455
rect 21867 10452 21879 10455
rect 22462 10452 22468 10464
rect 21867 10424 22468 10452
rect 21867 10421 21879 10424
rect 21821 10415 21879 10421
rect 22462 10412 22468 10424
rect 22520 10412 22526 10464
rect 23109 10455 23167 10461
rect 23109 10421 23121 10455
rect 23155 10452 23167 10455
rect 23198 10452 23204 10464
rect 23155 10424 23204 10452
rect 23155 10421 23167 10424
rect 23109 10415 23167 10421
rect 23198 10412 23204 10424
rect 23256 10412 23262 10464
rect 23308 10452 23336 10492
rect 25774 10480 25780 10532
rect 25832 10520 25838 10532
rect 30392 10520 30420 10560
rect 34974 10548 34980 10560
rect 35032 10588 35038 10600
rect 36538 10588 36544 10600
rect 35032 10560 36544 10588
rect 35032 10548 35038 10560
rect 36538 10548 36544 10560
rect 36596 10548 36602 10600
rect 37458 10548 37464 10600
rect 37516 10588 37522 10600
rect 37516 10560 37561 10588
rect 37516 10548 37522 10560
rect 37642 10548 37648 10600
rect 37700 10588 37706 10600
rect 37700 10560 37745 10588
rect 37700 10548 37706 10560
rect 34054 10520 34060 10532
rect 25832 10492 30420 10520
rect 30484 10492 34060 10520
rect 25832 10480 25838 10492
rect 30484 10452 30512 10492
rect 34054 10480 34060 10492
rect 34112 10480 34118 10532
rect 36081 10523 36139 10529
rect 36081 10489 36093 10523
rect 36127 10520 36139 10523
rect 37274 10520 37280 10532
rect 36127 10492 37280 10520
rect 36127 10489 36139 10492
rect 36081 10483 36139 10489
rect 37274 10480 37280 10492
rect 37332 10480 37338 10532
rect 37366 10480 37372 10532
rect 37424 10520 37430 10532
rect 38120 10520 38148 10619
rect 39114 10616 39120 10628
rect 39172 10616 39178 10668
rect 40494 10616 40500 10668
rect 40552 10656 40558 10668
rect 40773 10659 40831 10665
rect 40773 10656 40785 10659
rect 40552 10628 40785 10656
rect 40552 10616 40558 10628
rect 40773 10625 40785 10628
rect 40819 10625 40831 10659
rect 40773 10619 40831 10625
rect 40957 10659 41015 10665
rect 40957 10625 40969 10659
rect 41003 10656 41015 10659
rect 41598 10656 41604 10668
rect 41003 10628 41414 10656
rect 41559 10628 41604 10656
rect 41003 10625 41015 10628
rect 40957 10619 41015 10625
rect 38470 10548 38476 10600
rect 38528 10588 38534 10600
rect 39209 10591 39267 10597
rect 39209 10588 39221 10591
rect 38528 10560 39221 10588
rect 38528 10548 38534 10560
rect 39209 10557 39221 10560
rect 39255 10557 39267 10591
rect 39209 10551 39267 10557
rect 40865 10591 40923 10597
rect 40865 10557 40877 10591
rect 40911 10557 40923 10591
rect 41046 10588 41052 10600
rect 41007 10560 41052 10588
rect 40865 10551 40923 10557
rect 40494 10520 40500 10532
rect 37424 10492 37469 10520
rect 38120 10492 40500 10520
rect 37424 10480 37430 10492
rect 40494 10480 40500 10492
rect 40552 10480 40558 10532
rect 40880 10520 40908 10551
rect 41046 10548 41052 10560
rect 41104 10548 41110 10600
rect 41230 10520 41236 10532
rect 40880 10492 41236 10520
rect 41230 10480 41236 10492
rect 41288 10480 41294 10532
rect 41386 10520 41414 10628
rect 41598 10616 41604 10628
rect 41656 10616 41662 10668
rect 42613 10659 42671 10665
rect 42613 10625 42625 10659
rect 42659 10625 42671 10659
rect 42794 10656 42800 10668
rect 42755 10628 42800 10656
rect 42613 10619 42671 10625
rect 42628 10588 42656 10619
rect 42794 10616 42800 10628
rect 42852 10616 42858 10668
rect 42981 10659 43039 10665
rect 42981 10625 42993 10659
rect 43027 10656 43039 10659
rect 43530 10656 43536 10668
rect 43027 10628 43536 10656
rect 43027 10625 43039 10628
rect 42981 10619 43039 10625
rect 43530 10616 43536 10628
rect 43588 10616 43594 10668
rect 44174 10656 44180 10668
rect 44135 10628 44180 10656
rect 44174 10616 44180 10628
rect 44232 10616 44238 10668
rect 43346 10588 43352 10600
rect 42628 10560 43352 10588
rect 43346 10548 43352 10560
rect 43404 10548 43410 10600
rect 43165 10523 43223 10529
rect 43165 10520 43177 10523
rect 41386 10492 43177 10520
rect 43165 10489 43177 10492
rect 43211 10489 43223 10523
rect 43165 10483 43223 10489
rect 23308 10424 30512 10452
rect 30929 10455 30987 10461
rect 30929 10421 30941 10455
rect 30975 10452 30987 10455
rect 32490 10452 32496 10464
rect 30975 10424 32496 10452
rect 30975 10421 30987 10424
rect 30929 10415 30987 10421
rect 32490 10412 32496 10424
rect 32548 10412 32554 10464
rect 32766 10412 32772 10464
rect 32824 10452 32830 10464
rect 38473 10455 38531 10461
rect 38473 10452 38485 10455
rect 32824 10424 38485 10452
rect 32824 10412 32830 10424
rect 38473 10421 38485 10424
rect 38519 10421 38531 10455
rect 40586 10452 40592 10464
rect 40547 10424 40592 10452
rect 38473 10415 38531 10421
rect 40586 10412 40592 10424
rect 40644 10412 40650 10464
rect 40770 10412 40776 10464
rect 40828 10452 40834 10464
rect 41693 10455 41751 10461
rect 41693 10452 41705 10455
rect 40828 10424 41705 10452
rect 40828 10412 40834 10424
rect 41693 10421 41705 10424
rect 41739 10452 41751 10455
rect 42702 10452 42708 10464
rect 41739 10424 42708 10452
rect 41739 10421 41751 10424
rect 41693 10415 41751 10421
rect 42702 10412 42708 10424
rect 42760 10412 42766 10464
rect 1104 10362 44896 10384
rect 1104 10310 6424 10362
rect 6476 10310 6488 10362
rect 6540 10310 6552 10362
rect 6604 10310 6616 10362
rect 6668 10310 6680 10362
rect 6732 10310 17372 10362
rect 17424 10310 17436 10362
rect 17488 10310 17500 10362
rect 17552 10310 17564 10362
rect 17616 10310 17628 10362
rect 17680 10310 28320 10362
rect 28372 10310 28384 10362
rect 28436 10310 28448 10362
rect 28500 10310 28512 10362
rect 28564 10310 28576 10362
rect 28628 10310 39268 10362
rect 39320 10310 39332 10362
rect 39384 10310 39396 10362
rect 39448 10310 39460 10362
rect 39512 10310 39524 10362
rect 39576 10310 44896 10362
rect 1104 10288 44896 10310
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 4982 10248 4988 10260
rect 2924 10220 4988 10248
rect 2924 10208 2930 10220
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 5074 10208 5080 10260
rect 5132 10248 5138 10260
rect 5169 10251 5227 10257
rect 5169 10248 5181 10251
rect 5132 10220 5181 10248
rect 5132 10208 5138 10220
rect 5169 10217 5181 10220
rect 5215 10217 5227 10251
rect 5169 10211 5227 10217
rect 8941 10251 8999 10257
rect 8941 10217 8953 10251
rect 8987 10248 8999 10251
rect 9030 10248 9036 10260
rect 8987 10220 9036 10248
rect 8987 10217 8999 10220
rect 8941 10211 8999 10217
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 11054 10248 11060 10260
rect 10967 10220 11060 10248
rect 11054 10208 11060 10220
rect 11112 10248 11118 10260
rect 12342 10248 12348 10260
rect 11112 10220 12348 10248
rect 11112 10208 11118 10220
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 13078 10248 13084 10260
rect 12544 10220 13084 10248
rect 10686 10140 10692 10192
rect 10744 10180 10750 10192
rect 12434 10180 12440 10192
rect 10744 10152 12440 10180
rect 10744 10140 10750 10152
rect 12434 10140 12440 10152
rect 12492 10140 12498 10192
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 9490 10112 9496 10124
rect 8352 10084 9496 10112
rect 8352 10072 8358 10084
rect 9490 10072 9496 10084
rect 9548 10112 9554 10124
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9548 10084 9689 10112
rect 9548 10072 9554 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 12544 10112 12572 10220
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 14461 10251 14519 10257
rect 14461 10217 14473 10251
rect 14507 10248 14519 10251
rect 14550 10248 14556 10260
rect 14507 10220 14556 10248
rect 14507 10217 14519 10220
rect 14461 10211 14519 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 15010 10248 15016 10260
rect 14971 10220 15016 10248
rect 15010 10208 15016 10220
rect 15068 10208 15074 10260
rect 19702 10248 19708 10260
rect 19663 10220 19708 10248
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 22005 10251 22063 10257
rect 19812 10220 21588 10248
rect 13096 10180 13124 10208
rect 13096 10152 15884 10180
rect 12400 10084 12572 10112
rect 12713 10115 12771 10121
rect 12400 10072 12406 10084
rect 12713 10081 12725 10115
rect 12759 10112 12771 10115
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 12759 10084 14105 10112
rect 12759 10081 12771 10084
rect 12713 10075 12771 10081
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 15746 10112 15752 10124
rect 15707 10084 15752 10112
rect 14093 10075 14151 10081
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10044 2743 10047
rect 3234 10044 3240 10056
rect 2731 10016 3240 10044
rect 2731 10013 2743 10016
rect 2685 10007 2743 10013
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10044 3847 10047
rect 4430 10044 4436 10056
rect 3835 10016 4436 10044
rect 3835 10013 3847 10016
rect 3789 10007 3847 10013
rect 4430 10004 4436 10016
rect 4488 10004 4494 10056
rect 6086 10044 6092 10056
rect 6047 10016 6092 10044
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9398 10044 9404 10056
rect 9171 10016 9404 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 11517 10047 11575 10053
rect 11517 10044 11529 10047
rect 11388 10016 11529 10044
rect 11388 10004 11394 10016
rect 11517 10013 11529 10016
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 2222 9936 2228 9988
rect 2280 9976 2286 9988
rect 4034 9979 4092 9985
rect 4034 9976 4046 9979
rect 2280 9948 4046 9976
rect 2280 9936 2286 9948
rect 4034 9945 4046 9948
rect 4080 9945 4092 9979
rect 6822 9976 6828 9988
rect 4034 9939 4092 9945
rect 5092 9948 6828 9976
rect 3237 9911 3295 9917
rect 3237 9877 3249 9911
rect 3283 9908 3295 9911
rect 5092 9908 5120 9948
rect 6822 9936 6828 9948
rect 6880 9936 6886 9988
rect 8478 9936 8484 9988
rect 8536 9976 8542 9988
rect 9922 9979 9980 9985
rect 9922 9976 9934 9979
rect 8536 9948 9934 9976
rect 8536 9936 8542 9948
rect 9922 9945 9934 9948
rect 9968 9945 9980 9979
rect 9922 9939 9980 9945
rect 10410 9936 10416 9988
rect 10468 9976 10474 9988
rect 12728 9976 12756 10075
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 15856 10112 15884 10152
rect 17497 10115 17555 10121
rect 17497 10112 17509 10115
rect 15856 10084 17509 10112
rect 17497 10081 17509 10084
rect 17543 10081 17555 10115
rect 19812 10112 19840 10220
rect 21560 10180 21588 10220
rect 22005 10217 22017 10251
rect 22051 10248 22063 10251
rect 22278 10248 22284 10260
rect 22051 10220 22284 10248
rect 22051 10217 22063 10220
rect 22005 10211 22063 10217
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 22649 10251 22707 10257
rect 22649 10217 22661 10251
rect 22695 10248 22707 10251
rect 23014 10248 23020 10260
rect 22695 10220 23020 10248
rect 22695 10217 22707 10220
rect 22649 10211 22707 10217
rect 22664 10180 22692 10211
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 23753 10251 23811 10257
rect 23753 10217 23765 10251
rect 23799 10248 23811 10251
rect 25222 10248 25228 10260
rect 23799 10220 25228 10248
rect 23799 10217 23811 10220
rect 23753 10211 23811 10217
rect 25222 10208 25228 10220
rect 25280 10208 25286 10260
rect 25593 10251 25651 10257
rect 25593 10217 25605 10251
rect 25639 10248 25651 10251
rect 27246 10248 27252 10260
rect 25639 10220 27252 10248
rect 25639 10217 25651 10220
rect 25593 10211 25651 10217
rect 27246 10208 27252 10220
rect 27304 10208 27310 10260
rect 28966 10220 33180 10248
rect 21560 10152 22692 10180
rect 26970 10140 26976 10192
rect 27028 10180 27034 10192
rect 28966 10180 28994 10220
rect 27028 10152 28994 10180
rect 33152 10180 33180 10220
rect 33226 10208 33232 10260
rect 33284 10248 33290 10260
rect 33505 10251 33563 10257
rect 33505 10248 33517 10251
rect 33284 10220 33517 10248
rect 33284 10208 33290 10220
rect 33505 10217 33517 10220
rect 33551 10217 33563 10251
rect 35618 10248 35624 10260
rect 35579 10220 35624 10248
rect 33505 10211 33563 10217
rect 35618 10208 35624 10220
rect 35676 10208 35682 10260
rect 35802 10208 35808 10260
rect 35860 10248 35866 10260
rect 36265 10251 36323 10257
rect 36265 10248 36277 10251
rect 35860 10220 36277 10248
rect 35860 10208 35866 10220
rect 36265 10217 36277 10220
rect 36311 10217 36323 10251
rect 39301 10251 39359 10257
rect 36265 10211 36323 10217
rect 36372 10220 39252 10248
rect 36372 10180 36400 10220
rect 37550 10180 37556 10192
rect 33152 10152 36400 10180
rect 37292 10152 37556 10180
rect 27028 10140 27034 10152
rect 20622 10112 20628 10124
rect 17497 10075 17555 10081
rect 19306 10084 19840 10112
rect 20583 10084 20628 10112
rect 12894 10044 12900 10056
rect 12855 10016 12900 10044
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 14274 10044 14280 10056
rect 14235 10016 14280 10044
rect 14274 10004 14280 10016
rect 14332 10004 14338 10056
rect 14921 10047 14979 10053
rect 14921 10013 14933 10047
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 10468 9948 12756 9976
rect 10468 9936 10474 9948
rect 7374 9908 7380 9920
rect 3283 9880 5120 9908
rect 7335 9880 7380 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 12161 9911 12219 9917
rect 12161 9877 12173 9911
rect 12207 9908 12219 9911
rect 12250 9908 12256 9920
rect 12207 9880 12256 9908
rect 12207 9877 12219 9880
rect 12161 9871 12219 9877
rect 12250 9868 12256 9880
rect 12308 9868 12314 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12986 9908 12992 9920
rect 12492 9880 12992 9908
rect 12492 9868 12498 9880
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 13081 9911 13139 9917
rect 13081 9877 13093 9911
rect 13127 9908 13139 9911
rect 13630 9908 13636 9920
rect 13127 9880 13636 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 14936 9908 14964 10007
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18509 10047 18567 10053
rect 18509 10044 18521 10047
rect 18380 10016 18521 10044
rect 18380 10004 18386 10016
rect 18509 10013 18521 10016
rect 18555 10044 18567 10047
rect 19306 10044 19334 10084
rect 20622 10072 20628 10084
rect 20680 10072 20686 10124
rect 21726 10072 21732 10124
rect 21784 10112 21790 10124
rect 28810 10112 28816 10124
rect 21784 10084 28816 10112
rect 21784 10072 21790 10084
rect 19886 10044 19892 10056
rect 18555 10016 19334 10044
rect 19847 10016 19892 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 21174 10004 21180 10056
rect 21232 10044 21238 10056
rect 22002 10044 22008 10056
rect 21232 10016 22008 10044
rect 21232 10004 21238 10016
rect 22002 10004 22008 10016
rect 22060 10044 22066 10056
rect 22465 10047 22523 10053
rect 22465 10044 22477 10047
rect 22060 10016 22477 10044
rect 22060 10004 22066 10016
rect 22465 10013 22477 10016
rect 22511 10013 22523 10047
rect 22465 10007 22523 10013
rect 23661 10047 23719 10053
rect 23661 10013 23673 10047
rect 23707 10044 23719 10047
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 23707 10016 24777 10044
rect 23707 10013 23719 10016
rect 23661 10007 23719 10013
rect 24765 10013 24777 10016
rect 24811 10044 24823 10047
rect 25222 10044 25228 10056
rect 24811 10016 25228 10044
rect 24811 10013 24823 10016
rect 24765 10007 24823 10013
rect 25222 10004 25228 10016
rect 25280 10004 25286 10056
rect 25406 10044 25412 10056
rect 25367 10016 25412 10044
rect 25406 10004 25412 10016
rect 25464 10004 25470 10056
rect 26694 10044 26700 10056
rect 26655 10016 26700 10044
rect 26694 10004 26700 10016
rect 26752 10004 26758 10056
rect 26970 10044 26976 10056
rect 26931 10016 26976 10044
rect 26970 10004 26976 10016
rect 27028 10004 27034 10056
rect 27433 10047 27491 10053
rect 27433 10013 27445 10047
rect 27479 10044 27491 10047
rect 27522 10044 27528 10056
rect 27479 10016 27528 10044
rect 27479 10013 27491 10016
rect 27433 10007 27491 10013
rect 27522 10004 27528 10016
rect 27580 10044 27586 10056
rect 28460 10053 28488 10084
rect 28810 10072 28816 10084
rect 28868 10072 28874 10124
rect 29549 10115 29607 10121
rect 29549 10081 29561 10115
rect 29595 10112 29607 10115
rect 30282 10112 30288 10124
rect 29595 10084 30288 10112
rect 29595 10081 29607 10084
rect 29549 10075 29607 10081
rect 30282 10072 30288 10084
rect 30340 10112 30346 10124
rect 31757 10115 31815 10121
rect 31757 10112 31769 10115
rect 30340 10084 31769 10112
rect 30340 10072 30346 10084
rect 31757 10081 31769 10084
rect 31803 10081 31815 10115
rect 31757 10075 31815 10081
rect 34146 10072 34152 10124
rect 34204 10112 34210 10124
rect 34204 10084 35572 10112
rect 34204 10072 34210 10084
rect 28445 10047 28503 10053
rect 27580 10016 27752 10044
rect 27580 10004 27586 10016
rect 16022 9976 16028 9988
rect 15983 9948 16028 9976
rect 16022 9936 16028 9948
rect 16080 9936 16086 9988
rect 17770 9976 17776 9988
rect 17250 9948 17776 9976
rect 17770 9936 17776 9948
rect 17828 9936 17834 9988
rect 20892 9979 20950 9985
rect 20892 9945 20904 9979
rect 20938 9976 20950 9979
rect 25130 9976 25136 9988
rect 20938 9948 25136 9976
rect 20938 9945 20950 9948
rect 20892 9939 20950 9945
rect 25130 9936 25136 9948
rect 25188 9936 25194 9988
rect 26881 9979 26939 9985
rect 26881 9945 26893 9979
rect 26927 9976 26939 9979
rect 27614 9976 27620 9988
rect 26927 9948 27620 9976
rect 26927 9945 26939 9948
rect 26881 9939 26939 9945
rect 27614 9936 27620 9948
rect 27672 9936 27678 9988
rect 27724 9976 27752 10016
rect 28445 10013 28457 10047
rect 28491 10013 28503 10047
rect 28445 10007 28503 10013
rect 34514 10004 34520 10056
rect 34572 10044 34578 10056
rect 34701 10047 34759 10053
rect 34701 10044 34713 10047
rect 34572 10016 34713 10044
rect 34572 10004 34578 10016
rect 34701 10013 34713 10016
rect 34747 10013 34759 10047
rect 34701 10007 34759 10013
rect 34790 10004 34796 10056
rect 34848 10044 34854 10056
rect 35544 10053 35572 10084
rect 34885 10047 34943 10053
rect 34885 10044 34897 10047
rect 34848 10016 34897 10044
rect 34848 10004 34854 10016
rect 34885 10013 34897 10016
rect 34931 10013 34943 10047
rect 34885 10007 34943 10013
rect 35529 10047 35587 10053
rect 35529 10013 35541 10047
rect 35575 10013 35587 10047
rect 36170 10044 36176 10056
rect 36131 10016 36176 10044
rect 35529 10007 35587 10013
rect 36170 10004 36176 10016
rect 36228 10004 36234 10056
rect 37292 10053 37320 10152
rect 37550 10140 37556 10152
rect 37608 10140 37614 10192
rect 39224 10180 39252 10220
rect 39301 10217 39313 10251
rect 39347 10248 39359 10251
rect 39666 10248 39672 10260
rect 39347 10220 39672 10248
rect 39347 10217 39359 10220
rect 39301 10211 39359 10217
rect 39666 10208 39672 10220
rect 39724 10248 39730 10260
rect 40126 10248 40132 10260
rect 39724 10220 40132 10248
rect 39724 10208 39730 10220
rect 40126 10208 40132 10220
rect 40184 10208 40190 10260
rect 40310 10248 40316 10260
rect 40271 10220 40316 10248
rect 40310 10208 40316 10220
rect 40368 10208 40374 10260
rect 40494 10248 40500 10260
rect 40455 10220 40500 10248
rect 40494 10208 40500 10220
rect 40552 10208 40558 10260
rect 40586 10208 40592 10260
rect 40644 10248 40650 10260
rect 40644 10220 42288 10248
rect 40644 10208 40650 10220
rect 41601 10183 41659 10189
rect 39224 10152 41414 10180
rect 37918 10112 37924 10124
rect 37879 10084 37924 10112
rect 37918 10072 37924 10084
rect 37976 10072 37982 10124
rect 41386 10112 41414 10152
rect 41601 10149 41613 10183
rect 41647 10180 41659 10183
rect 41647 10152 42196 10180
rect 41647 10149 41659 10152
rect 41601 10143 41659 10149
rect 41966 10112 41972 10124
rect 41386 10084 41972 10112
rect 41966 10072 41972 10084
rect 42024 10072 42030 10124
rect 37277 10047 37335 10053
rect 37277 10013 37289 10047
rect 37323 10013 37335 10047
rect 37277 10007 37335 10013
rect 37461 10047 37519 10053
rect 37461 10013 37473 10047
rect 37507 10044 37519 10047
rect 38470 10044 38476 10056
rect 37507 10016 38476 10044
rect 37507 10013 37519 10016
rect 37461 10007 37519 10013
rect 38470 10004 38476 10016
rect 38528 10004 38534 10056
rect 40126 10044 40132 10056
rect 40087 10016 40132 10044
rect 40126 10004 40132 10016
rect 40184 10004 40190 10056
rect 40310 10044 40316 10056
rect 40271 10016 40316 10044
rect 40310 10004 40316 10016
rect 40368 10004 40374 10056
rect 40678 10004 40684 10056
rect 40736 10044 40742 10056
rect 41138 10053 41144 10056
rect 40946 10047 41004 10053
rect 40946 10044 40958 10047
rect 40736 10016 40958 10044
rect 40736 10004 40742 10016
rect 40946 10013 40958 10016
rect 40992 10013 41004 10047
rect 40946 10007 41004 10013
rect 41105 10047 41144 10053
rect 41105 10013 41117 10047
rect 41105 10007 41144 10013
rect 41138 10004 41144 10007
rect 41196 10004 41202 10056
rect 41233 10047 41291 10053
rect 41233 10013 41245 10047
rect 41279 10013 41291 10047
rect 41233 10007 41291 10013
rect 29825 9979 29883 9985
rect 27724 9948 28672 9976
rect 15286 9908 15292 9920
rect 14936 9880 15292 9908
rect 15286 9868 15292 9880
rect 15344 9908 15350 9920
rect 16666 9908 16672 9920
rect 15344 9880 16672 9908
rect 15344 9868 15350 9880
rect 16666 9868 16672 9880
rect 16724 9908 16730 9920
rect 18322 9908 18328 9920
rect 16724 9880 18328 9908
rect 16724 9868 16730 9880
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 18506 9868 18512 9920
rect 18564 9908 18570 9920
rect 18601 9911 18659 9917
rect 18601 9908 18613 9911
rect 18564 9880 18613 9908
rect 18564 9868 18570 9880
rect 18601 9877 18613 9880
rect 18647 9877 18659 9911
rect 18601 9871 18659 9877
rect 18690 9868 18696 9920
rect 18748 9908 18754 9920
rect 22094 9908 22100 9920
rect 18748 9880 22100 9908
rect 18748 9868 18754 9880
rect 22094 9868 22100 9880
rect 22152 9868 22158 9920
rect 24857 9911 24915 9917
rect 24857 9877 24869 9911
rect 24903 9908 24915 9911
rect 24946 9908 24952 9920
rect 24903 9880 24952 9908
rect 24903 9877 24915 9880
rect 24857 9871 24915 9877
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 26326 9868 26332 9920
rect 26384 9908 26390 9920
rect 26513 9911 26571 9917
rect 26513 9908 26525 9911
rect 26384 9880 26525 9908
rect 26384 9868 26390 9880
rect 26513 9877 26525 9880
rect 26559 9877 26571 9911
rect 26513 9871 26571 9877
rect 27430 9868 27436 9920
rect 27488 9908 27494 9920
rect 27525 9911 27583 9917
rect 27525 9908 27537 9911
rect 27488 9880 27537 9908
rect 27488 9868 27494 9880
rect 27525 9877 27537 9880
rect 27571 9877 27583 9911
rect 27525 9871 27583 9877
rect 28442 9868 28448 9920
rect 28500 9908 28506 9920
rect 28537 9911 28595 9917
rect 28537 9908 28549 9911
rect 28500 9880 28549 9908
rect 28500 9868 28506 9880
rect 28537 9877 28549 9880
rect 28583 9877 28595 9911
rect 28644 9908 28672 9948
rect 29825 9945 29837 9979
rect 29871 9976 29883 9979
rect 29914 9976 29920 9988
rect 29871 9948 29920 9976
rect 29871 9945 29883 9948
rect 29825 9939 29883 9945
rect 29914 9936 29920 9948
rect 29972 9936 29978 9988
rect 30374 9936 30380 9988
rect 30432 9936 30438 9988
rect 32033 9979 32091 9985
rect 32033 9976 32045 9979
rect 31726 9948 32045 9976
rect 30006 9908 30012 9920
rect 28644 9880 30012 9908
rect 28537 9871 28595 9877
rect 30006 9868 30012 9880
rect 30064 9868 30070 9920
rect 31297 9911 31355 9917
rect 31297 9877 31309 9911
rect 31343 9908 31355 9911
rect 31726 9908 31754 9948
rect 32033 9945 32045 9948
rect 32079 9945 32091 9979
rect 32033 9939 32091 9945
rect 32490 9936 32496 9988
rect 32548 9936 32554 9988
rect 36538 9936 36544 9988
rect 36596 9976 36602 9988
rect 37642 9976 37648 9988
rect 36596 9948 37648 9976
rect 36596 9936 36602 9948
rect 37642 9936 37648 9948
rect 37700 9936 37706 9988
rect 38188 9979 38246 9985
rect 38188 9945 38200 9979
rect 38234 9976 38246 9979
rect 38838 9976 38844 9988
rect 38234 9948 38844 9976
rect 38234 9945 38246 9948
rect 38188 9939 38246 9945
rect 38838 9936 38844 9948
rect 38896 9936 38902 9988
rect 39853 9979 39911 9985
rect 39853 9945 39865 9979
rect 39899 9976 39911 9979
rect 41248 9976 41276 10007
rect 41322 10004 41328 10056
rect 41380 10044 41386 10056
rect 41506 10053 41512 10056
rect 41463 10047 41512 10053
rect 41380 10016 41425 10044
rect 41380 10004 41386 10016
rect 41463 10013 41475 10047
rect 41509 10013 41512 10047
rect 41463 10007 41512 10013
rect 41506 10004 41512 10007
rect 41564 10004 41570 10056
rect 42058 10044 42064 10056
rect 41616 10016 42064 10044
rect 41616 9976 41644 10016
rect 42058 10004 42064 10016
rect 42116 10004 42122 10056
rect 42168 10053 42196 10152
rect 42260 10053 42288 10220
rect 42794 10208 42800 10260
rect 42852 10248 42858 10260
rect 43349 10251 43407 10257
rect 43349 10248 43361 10251
rect 42852 10220 43361 10248
rect 42852 10208 42858 10220
rect 43349 10217 43361 10220
rect 43395 10217 43407 10251
rect 43349 10211 43407 10217
rect 42153 10047 42211 10053
rect 42153 10013 42165 10047
rect 42199 10013 42211 10047
rect 42153 10007 42211 10013
rect 42245 10047 42303 10053
rect 42245 10013 42257 10047
rect 42291 10013 42303 10047
rect 42245 10007 42303 10013
rect 42334 10004 42340 10056
rect 42392 10044 42398 10056
rect 42981 10047 43039 10053
rect 42392 10016 42437 10044
rect 42392 10004 42398 10016
rect 42981 10013 42993 10047
rect 43027 10044 43039 10047
rect 43438 10044 43444 10056
rect 43027 10016 43444 10044
rect 43027 10013 43039 10016
rect 42981 10007 43039 10013
rect 43438 10004 43444 10016
rect 43496 10004 43502 10056
rect 39899 9948 40908 9976
rect 41248 9948 41644 9976
rect 39899 9945 39911 9948
rect 39853 9939 39911 9945
rect 40880 9920 40908 9948
rect 41966 9936 41972 9988
rect 42024 9976 42030 9988
rect 42521 9979 42579 9985
rect 42521 9976 42533 9979
rect 42024 9948 42533 9976
rect 42024 9936 42030 9948
rect 42521 9945 42533 9948
rect 42567 9945 42579 9979
rect 42521 9939 42579 9945
rect 43165 9979 43223 9985
rect 43165 9945 43177 9979
rect 43211 9976 43223 9979
rect 43211 9948 43245 9976
rect 43211 9945 43223 9948
rect 43165 9939 43223 9945
rect 35066 9908 35072 9920
rect 31343 9880 31754 9908
rect 35027 9880 35072 9908
rect 31343 9877 31355 9880
rect 31297 9871 31355 9877
rect 35066 9868 35072 9880
rect 35124 9868 35130 9920
rect 37369 9911 37427 9917
rect 37369 9877 37381 9911
rect 37415 9908 37427 9911
rect 39022 9908 39028 9920
rect 37415 9880 39028 9908
rect 37415 9877 37427 9880
rect 37369 9871 37427 9877
rect 39022 9868 39028 9880
rect 39080 9868 39086 9920
rect 40862 9868 40868 9920
rect 40920 9868 40926 9920
rect 42150 9868 42156 9920
rect 42208 9908 42214 9920
rect 43180 9908 43208 9939
rect 43622 9908 43628 9920
rect 42208 9880 43628 9908
rect 42208 9868 42214 9880
rect 43622 9868 43628 9880
rect 43680 9868 43686 9920
rect 1104 9818 45056 9840
rect 1104 9766 11898 9818
rect 11950 9766 11962 9818
rect 12014 9766 12026 9818
rect 12078 9766 12090 9818
rect 12142 9766 12154 9818
rect 12206 9766 22846 9818
rect 22898 9766 22910 9818
rect 22962 9766 22974 9818
rect 23026 9766 23038 9818
rect 23090 9766 23102 9818
rect 23154 9766 33794 9818
rect 33846 9766 33858 9818
rect 33910 9766 33922 9818
rect 33974 9766 33986 9818
rect 34038 9766 34050 9818
rect 34102 9766 44742 9818
rect 44794 9766 44806 9818
rect 44858 9766 44870 9818
rect 44922 9766 44934 9818
rect 44986 9766 44998 9818
rect 45050 9766 45056 9818
rect 1104 9744 45056 9766
rect 5077 9707 5135 9713
rect 5077 9673 5089 9707
rect 5123 9673 5135 9707
rect 5077 9667 5135 9673
rect 11977 9707 12035 9713
rect 11977 9673 11989 9707
rect 12023 9704 12035 9707
rect 12250 9704 12256 9716
rect 12023 9676 12256 9704
rect 12023 9673 12035 9676
rect 11977 9667 12035 9673
rect 3510 9636 3516 9648
rect 1872 9608 3516 9636
rect 1872 9577 1900 9608
rect 3510 9596 3516 9608
rect 3568 9596 3574 9648
rect 3964 9639 4022 9645
rect 3964 9605 3976 9639
rect 4010 9636 4022 9639
rect 4890 9636 4896 9648
rect 4010 9608 4896 9636
rect 4010 9605 4022 9608
rect 3964 9599 4022 9605
rect 4890 9596 4896 9608
rect 4948 9596 4954 9648
rect 5092 9636 5120 9667
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 15746 9704 15752 9716
rect 14752 9676 15752 9704
rect 9760 9639 9818 9645
rect 5092 9608 7604 9636
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9537 1915 9571
rect 1857 9531 1915 9537
rect 2124 9571 2182 9577
rect 2124 9537 2136 9571
rect 2170 9568 2182 9571
rect 3418 9568 3424 9580
rect 2170 9540 3424 9568
rect 2170 9537 2182 9540
rect 2124 9531 2182 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 3620 9540 5733 9568
rect 3234 9432 3240 9444
rect 3195 9404 3240 9432
rect 3234 9392 3240 9404
rect 3292 9392 3298 9444
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 3620 9364 3648 9540
rect 5721 9537 5733 9540
rect 5767 9537 5779 9571
rect 6730 9568 6736 9580
rect 6691 9540 6736 9568
rect 5721 9531 5779 9537
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 6822 9528 6828 9580
rect 6880 9568 6886 9580
rect 7576 9577 7604 9608
rect 9760 9605 9772 9639
rect 9806 9636 9818 9639
rect 11054 9636 11060 9648
rect 9806 9608 11060 9636
rect 9806 9605 9818 9608
rect 9760 9599 9818 9605
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 11885 9639 11943 9645
rect 11885 9605 11897 9639
rect 11931 9636 11943 9639
rect 12434 9636 12440 9648
rect 11931 9608 12440 9636
rect 11931 9605 11943 9608
rect 11885 9599 11943 9605
rect 12434 9596 12440 9608
rect 12492 9636 12498 9648
rect 12894 9636 12900 9648
rect 12492 9608 12900 9636
rect 12492 9596 12498 9608
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 14752 9645 14780 9676
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 19886 9664 19892 9716
rect 19944 9704 19950 9716
rect 20165 9707 20223 9713
rect 20165 9704 20177 9707
rect 19944 9676 20177 9704
rect 19944 9664 19950 9676
rect 20165 9673 20177 9676
rect 20211 9673 20223 9707
rect 25130 9704 25136 9716
rect 25091 9676 25136 9704
rect 20165 9667 20223 9673
rect 25130 9664 25136 9676
rect 25188 9664 25194 9716
rect 25222 9664 25228 9716
rect 25280 9704 25286 9716
rect 25777 9707 25835 9713
rect 25777 9704 25789 9707
rect 25280 9676 25789 9704
rect 25280 9664 25286 9676
rect 25777 9673 25789 9676
rect 25823 9704 25835 9707
rect 27522 9704 27528 9716
rect 25823 9676 27528 9704
rect 25823 9673 25835 9676
rect 25777 9667 25835 9673
rect 27522 9664 27528 9676
rect 27580 9664 27586 9716
rect 30006 9664 30012 9716
rect 30064 9664 30070 9716
rect 31021 9707 31079 9713
rect 31021 9673 31033 9707
rect 31067 9673 31079 9707
rect 31021 9667 31079 9673
rect 32591 9707 32649 9713
rect 32591 9673 32603 9707
rect 32637 9673 32649 9707
rect 32591 9667 32649 9673
rect 33965 9707 34023 9713
rect 33965 9673 33977 9707
rect 34011 9704 34023 9707
rect 34882 9704 34888 9716
rect 34011 9676 34888 9704
rect 34011 9673 34023 9676
rect 33965 9667 34023 9673
rect 14737 9639 14795 9645
rect 14737 9605 14749 9639
rect 14783 9605 14795 9639
rect 18046 9636 18052 9648
rect 14737 9599 14795 9605
rect 17512 9608 18052 9636
rect 7561 9571 7619 9577
rect 6880 9540 6925 9568
rect 6880 9528 6886 9540
rect 7561 9537 7573 9571
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8260 9540 8861 9568
rect 8260 9528 8266 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 9490 9568 9496 9580
rect 9451 9540 9496 9568
rect 8849 9531 8907 9537
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 12342 9568 12348 9580
rect 9600 9540 12348 9568
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 6914 9500 6920 9512
rect 3752 9472 3797 9500
rect 6875 9472 6920 9500
rect 3752 9460 3758 9472
rect 6914 9460 6920 9472
rect 6972 9500 6978 9512
rect 9600 9500 9628 9540
rect 12084 9509 12112 9540
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 12986 9568 12992 9580
rect 12947 9540 12992 9568
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13538 9528 13544 9580
rect 13596 9568 13602 9580
rect 15749 9571 15807 9577
rect 15749 9568 15761 9571
rect 13596 9540 15761 9568
rect 13596 9528 13602 9540
rect 15749 9537 15761 9540
rect 15795 9537 15807 9571
rect 16666 9568 16672 9580
rect 16627 9540 16672 9568
rect 15749 9531 15807 9537
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 17512 9577 17540 9608
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 18506 9596 18512 9648
rect 18564 9596 18570 9648
rect 19334 9596 19340 9648
rect 19392 9636 19398 9648
rect 20622 9636 20628 9648
rect 19392 9608 20628 9636
rect 19392 9596 19398 9608
rect 20622 9596 20628 9608
rect 20680 9596 20686 9648
rect 23658 9636 23664 9648
rect 23619 9608 23664 9636
rect 23658 9596 23664 9608
rect 23716 9596 23722 9648
rect 24946 9636 24952 9648
rect 24886 9608 24952 9636
rect 24946 9596 24952 9608
rect 25004 9596 25010 9648
rect 28442 9596 28448 9648
rect 28500 9596 28506 9648
rect 30024 9636 30052 9664
rect 31036 9636 31064 9667
rect 31570 9636 31576 9648
rect 30024 9608 30512 9636
rect 31036 9608 31576 9636
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9537 17555 9571
rect 17497 9531 17555 9537
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 20809 9571 20867 9577
rect 20809 9568 20821 9571
rect 19484 9540 20821 9568
rect 19484 9528 19490 9540
rect 20809 9537 20821 9540
rect 20855 9537 20867 9571
rect 20809 9531 20867 9537
rect 25406 9528 25412 9580
rect 25464 9568 25470 9580
rect 25593 9571 25651 9577
rect 25593 9568 25605 9571
rect 25464 9540 25605 9568
rect 25464 9528 25470 9540
rect 25593 9537 25605 9540
rect 25639 9537 25651 9571
rect 25593 9531 25651 9537
rect 29908 9571 29966 9577
rect 29908 9537 29920 9571
rect 29954 9568 29966 9571
rect 30374 9568 30380 9580
rect 29954 9540 30380 9568
rect 29954 9537 29966 9540
rect 29908 9531 29966 9537
rect 30374 9528 30380 9540
rect 30432 9528 30438 9580
rect 30484 9568 30512 9608
rect 31570 9596 31576 9608
rect 31628 9636 31634 9648
rect 32600 9636 32628 9667
rect 34882 9664 34888 9676
rect 34940 9664 34946 9716
rect 35066 9664 35072 9716
rect 35124 9704 35130 9716
rect 38841 9707 38899 9713
rect 35124 9676 35848 9704
rect 35124 9664 35130 9676
rect 35621 9639 35679 9645
rect 35621 9636 35633 9639
rect 31628 9608 35633 9636
rect 31628 9596 31634 9608
rect 35621 9605 35633 9608
rect 35667 9605 35679 9639
rect 35820 9636 35848 9676
rect 38488 9676 38792 9704
rect 38289 9639 38347 9645
rect 35820 9608 36400 9636
rect 35621 9599 35679 9605
rect 31110 9568 31116 9580
rect 30484 9540 31116 9568
rect 31110 9528 31116 9540
rect 31168 9528 31174 9580
rect 32674 9568 32680 9580
rect 32635 9540 32680 9568
rect 32674 9528 32680 9540
rect 32732 9528 32738 9580
rect 32766 9528 32772 9580
rect 32824 9568 32830 9580
rect 33045 9571 33103 9577
rect 32824 9540 32869 9568
rect 32824 9528 32830 9540
rect 33045 9537 33057 9571
rect 33091 9568 33103 9571
rect 33226 9568 33232 9580
rect 33091 9540 33232 9568
rect 33091 9537 33103 9540
rect 33045 9531 33103 9537
rect 33226 9528 33232 9540
rect 33284 9528 33290 9580
rect 33410 9528 33416 9580
rect 33468 9568 33474 9580
rect 33873 9571 33931 9577
rect 33873 9568 33885 9571
rect 33468 9540 33885 9568
rect 33468 9528 33474 9540
rect 33873 9537 33885 9540
rect 33919 9537 33931 9571
rect 33873 9531 33931 9537
rect 34885 9571 34943 9577
rect 34885 9537 34897 9571
rect 34931 9568 34943 9571
rect 35802 9568 35808 9580
rect 34931 9540 35664 9568
rect 35763 9540 35808 9568
rect 34931 9537 34943 9540
rect 34885 9531 34943 9537
rect 6972 9472 9628 9500
rect 12069 9503 12127 9509
rect 6972 9460 6978 9472
rect 12069 9469 12081 9503
rect 12115 9469 12127 9503
rect 15838 9500 15844 9512
rect 15799 9472 15844 9500
rect 12069 9463 12127 9469
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 15930 9460 15936 9512
rect 15988 9500 15994 9512
rect 16390 9500 16396 9512
rect 15988 9472 16396 9500
rect 15988 9460 15994 9472
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 17034 9460 17040 9512
rect 17092 9500 17098 9512
rect 17773 9503 17831 9509
rect 17773 9500 17785 9503
rect 17092 9472 17785 9500
rect 17092 9460 17098 9472
rect 17773 9469 17785 9472
rect 17819 9469 17831 9503
rect 17773 9463 17831 9469
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 19751 9472 20576 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 6365 9435 6423 9441
rect 6365 9432 6377 9435
rect 4632 9404 6377 9432
rect 2832 9336 3648 9364
rect 2832 9324 2838 9336
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 4632 9364 4660 9404
rect 6365 9401 6377 9404
rect 6411 9401 6423 9435
rect 15381 9435 15439 9441
rect 6365 9395 6423 9401
rect 6656 9404 9444 9432
rect 5534 9364 5540 9376
rect 4028 9336 4660 9364
rect 5495 9336 5540 9364
rect 4028 9324 4034 9336
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 5718 9324 5724 9376
rect 5776 9364 5782 9376
rect 6656 9364 6684 9404
rect 8202 9364 8208 9376
rect 5776 9336 6684 9364
rect 8163 9336 8208 9364
rect 5776 9324 5782 9336
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 8665 9367 8723 9373
rect 8665 9333 8677 9367
rect 8711 9364 8723 9367
rect 9306 9364 9312 9376
rect 8711 9336 9312 9364
rect 8711 9333 8723 9336
rect 8665 9327 8723 9333
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 9416 9364 9444 9404
rect 15381 9401 15393 9435
rect 15427 9432 15439 9435
rect 17126 9432 17132 9444
rect 15427 9404 17132 9432
rect 15427 9401 15439 9404
rect 15381 9395 15439 9401
rect 17126 9392 17132 9404
rect 17184 9392 17190 9444
rect 19245 9435 19303 9441
rect 19245 9401 19257 9435
rect 19291 9432 19303 9435
rect 19981 9435 20039 9441
rect 19981 9432 19993 9435
rect 19291 9404 19993 9432
rect 19291 9401 19303 9404
rect 19245 9395 19303 9401
rect 19720 9376 19748 9404
rect 19981 9401 19993 9404
rect 20027 9401 20039 9435
rect 20548 9432 20576 9472
rect 20622 9460 20628 9512
rect 20680 9500 20686 9512
rect 20680 9472 20725 9500
rect 20680 9460 20686 9472
rect 21726 9460 21732 9512
rect 21784 9500 21790 9512
rect 21821 9503 21879 9509
rect 21821 9500 21833 9503
rect 21784 9472 21833 9500
rect 21784 9460 21790 9472
rect 21821 9469 21833 9472
rect 21867 9469 21879 9503
rect 21821 9463 21879 9469
rect 22002 9460 22008 9512
rect 22060 9500 22066 9512
rect 22097 9503 22155 9509
rect 22097 9500 22109 9503
rect 22060 9472 22109 9500
rect 22060 9460 22066 9472
rect 22097 9469 22109 9472
rect 22143 9469 22155 9503
rect 23382 9500 23388 9512
rect 23343 9472 23388 9500
rect 22097 9463 22155 9469
rect 21174 9432 21180 9444
rect 20548 9404 21180 9432
rect 19981 9395 20039 9401
rect 21174 9392 21180 9404
rect 21232 9392 21238 9444
rect 22112 9432 22140 9463
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 25424 9500 25452 9528
rect 23492 9472 25452 9500
rect 23492 9432 23520 9472
rect 26234 9460 26240 9512
rect 26292 9500 26298 9512
rect 27433 9503 27491 9509
rect 27433 9500 27445 9503
rect 26292 9472 27445 9500
rect 26292 9460 26298 9472
rect 27433 9469 27445 9472
rect 27479 9469 27491 9503
rect 27433 9463 27491 9469
rect 27709 9503 27767 9509
rect 27709 9469 27721 9503
rect 27755 9500 27767 9503
rect 27798 9500 27804 9512
rect 27755 9472 27804 9500
rect 27755 9469 27767 9472
rect 27709 9463 27767 9469
rect 22112 9404 23520 9432
rect 10873 9367 10931 9373
rect 10873 9364 10885 9367
rect 9416 9336 10885 9364
rect 10873 9333 10885 9336
rect 10919 9364 10931 9367
rect 11330 9364 11336 9376
rect 10919 9336 11336 9364
rect 10919 9333 10931 9336
rect 10873 9327 10931 9333
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 11514 9364 11520 9376
rect 11475 9336 11520 9364
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 14642 9324 14648 9376
rect 14700 9364 14706 9376
rect 16482 9364 16488 9376
rect 14700 9336 16488 9364
rect 14700 9324 14706 9336
rect 16482 9324 16488 9336
rect 16540 9324 16546 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 16761 9367 16819 9373
rect 16761 9364 16773 9367
rect 16724 9336 16773 9364
rect 16724 9324 16730 9336
rect 16761 9333 16773 9336
rect 16807 9333 16819 9367
rect 16761 9327 16819 9333
rect 19702 9324 19708 9376
rect 19760 9324 19766 9376
rect 20993 9367 21051 9373
rect 20993 9333 21005 9367
rect 21039 9364 21051 9367
rect 21266 9364 21272 9376
rect 21039 9336 21272 9364
rect 21039 9333 21051 9336
rect 20993 9327 21051 9333
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 27448 9364 27476 9463
rect 27798 9460 27804 9472
rect 27856 9460 27862 9512
rect 29638 9500 29644 9512
rect 29012 9472 29644 9500
rect 29012 9364 29040 9472
rect 29638 9460 29644 9472
rect 29696 9460 29702 9512
rect 32953 9503 33011 9509
rect 32953 9500 32965 9503
rect 31726 9472 32965 9500
rect 27448 9336 29040 9364
rect 29181 9367 29239 9373
rect 29181 9333 29193 9367
rect 29227 9364 29239 9367
rect 29822 9364 29828 9376
rect 29227 9336 29828 9364
rect 29227 9333 29239 9336
rect 29181 9327 29239 9333
rect 29822 9324 29828 9336
rect 29880 9364 29886 9376
rect 31726 9364 31754 9472
rect 32953 9469 32965 9472
rect 32999 9469 33011 9503
rect 32953 9463 33011 9469
rect 33134 9460 33140 9512
rect 33192 9500 33198 9512
rect 34057 9503 34115 9509
rect 34057 9500 34069 9503
rect 33192 9472 34069 9500
rect 33192 9460 33198 9472
rect 34057 9469 34069 9472
rect 34103 9500 34115 9503
rect 34238 9500 34244 9512
rect 34103 9472 34244 9500
rect 34103 9469 34115 9472
rect 34057 9463 34115 9469
rect 34238 9460 34244 9472
rect 34296 9460 34302 9512
rect 34514 9460 34520 9512
rect 34572 9500 34578 9512
rect 35161 9503 35219 9509
rect 35161 9500 35173 9503
rect 34572 9472 35173 9500
rect 34572 9460 34578 9472
rect 35161 9469 35173 9472
rect 35207 9469 35219 9503
rect 35636 9500 35664 9540
rect 35802 9528 35808 9540
rect 35860 9528 35866 9580
rect 35894 9528 35900 9580
rect 35952 9568 35958 9580
rect 36372 9577 36400 9608
rect 38289 9605 38301 9639
rect 38335 9636 38347 9639
rect 38488 9636 38516 9676
rect 38654 9636 38660 9648
rect 38335 9608 38516 9636
rect 38615 9608 38660 9636
rect 38335 9605 38347 9608
rect 38289 9599 38347 9605
rect 38654 9596 38660 9608
rect 38712 9596 38718 9648
rect 38764 9636 38792 9676
rect 38841 9673 38853 9707
rect 38887 9704 38899 9707
rect 39114 9704 39120 9716
rect 38887 9676 39120 9704
rect 38887 9673 38899 9676
rect 38841 9667 38899 9673
rect 39114 9664 39120 9676
rect 39172 9664 39178 9716
rect 40770 9674 40776 9716
rect 40696 9664 40776 9674
rect 40828 9664 40834 9716
rect 41230 9704 41236 9716
rect 41191 9676 41236 9704
rect 41230 9664 41236 9676
rect 41288 9664 41294 9716
rect 41432 9676 42012 9704
rect 39666 9636 39672 9648
rect 38764 9608 39672 9636
rect 39666 9596 39672 9608
rect 39724 9596 39730 9648
rect 40696 9646 40807 9664
rect 36357 9571 36415 9577
rect 35952 9540 35997 9568
rect 35952 9528 35958 9540
rect 36357 9537 36369 9571
rect 36403 9537 36415 9571
rect 36538 9568 36544 9580
rect 36499 9540 36544 9568
rect 36357 9531 36415 9537
rect 36538 9528 36544 9540
rect 36596 9528 36602 9580
rect 38473 9571 38531 9577
rect 38473 9537 38485 9571
rect 38519 9537 38531 9571
rect 38473 9531 38531 9537
rect 36449 9503 36507 9509
rect 36449 9500 36461 9503
rect 35636 9472 36461 9500
rect 35161 9463 35219 9469
rect 36449 9469 36461 9472
rect 36495 9469 36507 9503
rect 38488 9500 38516 9531
rect 38562 9528 38568 9580
rect 38620 9568 38626 9580
rect 38620 9540 38665 9568
rect 38620 9528 38626 9540
rect 38746 9528 38752 9580
rect 38804 9568 38810 9580
rect 38804 9540 40080 9568
rect 38804 9528 38810 9540
rect 38930 9500 38936 9512
rect 38488 9472 38936 9500
rect 36449 9463 36507 9469
rect 33505 9435 33563 9441
rect 33505 9401 33517 9435
rect 33551 9432 33563 9435
rect 33594 9432 33600 9444
rect 33551 9404 33600 9432
rect 33551 9401 33563 9404
rect 33505 9395 33563 9401
rect 33594 9392 33600 9404
rect 33652 9392 33658 9444
rect 35176 9432 35204 9463
rect 38930 9460 38936 9472
rect 38988 9460 38994 9512
rect 39301 9503 39359 9509
rect 39301 9469 39313 9503
rect 39347 9500 39359 9503
rect 39850 9500 39856 9512
rect 39347 9472 39856 9500
rect 39347 9469 39359 9472
rect 39301 9463 39359 9469
rect 39850 9460 39856 9472
rect 39908 9460 39914 9512
rect 40052 9500 40080 9540
rect 40126 9528 40132 9580
rect 40184 9568 40190 9580
rect 40696 9577 40724 9646
rect 40865 9639 40923 9645
rect 40865 9605 40877 9639
rect 40911 9636 40923 9639
rect 41432 9636 41460 9676
rect 41984 9636 42012 9676
rect 42334 9664 42340 9716
rect 42392 9704 42398 9716
rect 42429 9707 42487 9713
rect 42429 9704 42441 9707
rect 42392 9676 42441 9704
rect 42392 9664 42398 9676
rect 42429 9673 42441 9676
rect 42475 9673 42487 9707
rect 42429 9667 42487 9673
rect 40911 9608 41460 9636
rect 41524 9608 41920 9636
rect 41984 9608 42656 9636
rect 40911 9605 40923 9608
rect 40865 9599 40923 9605
rect 40589 9571 40647 9577
rect 40589 9568 40601 9571
rect 40184 9540 40601 9568
rect 40184 9528 40190 9540
rect 40589 9537 40601 9540
rect 40635 9537 40647 9571
rect 40589 9531 40647 9537
rect 40682 9571 40740 9577
rect 40682 9537 40694 9571
rect 40728 9537 40740 9571
rect 40954 9568 40960 9580
rect 40915 9540 40960 9568
rect 40682 9531 40740 9537
rect 40954 9528 40960 9540
rect 41012 9528 41018 9580
rect 41095 9571 41153 9577
rect 41095 9537 41107 9571
rect 41141 9568 41153 9571
rect 41141 9540 41276 9568
rect 41141 9537 41153 9540
rect 41095 9531 41153 9537
rect 41248 9500 41276 9540
rect 41322 9528 41328 9580
rect 41380 9568 41386 9580
rect 41524 9568 41552 9608
rect 41892 9577 41920 9608
rect 42628 9580 42656 9608
rect 43346 9596 43352 9648
rect 43404 9636 43410 9648
rect 43533 9639 43591 9645
rect 43533 9636 43545 9639
rect 43404 9608 43545 9636
rect 43404 9596 43410 9608
rect 43533 9605 43545 9608
rect 43579 9605 43591 9639
rect 43533 9599 43591 9605
rect 41380 9540 41552 9568
rect 41693 9571 41751 9577
rect 41380 9528 41386 9540
rect 41693 9537 41705 9571
rect 41739 9537 41751 9571
rect 41693 9531 41751 9537
rect 41877 9571 41935 9577
rect 41877 9537 41889 9571
rect 41923 9537 41935 9571
rect 42610 9568 42616 9580
rect 42571 9540 42616 9568
rect 41877 9531 41935 9537
rect 41708 9500 41736 9531
rect 42610 9528 42616 9540
rect 42668 9528 42674 9580
rect 42702 9528 42708 9580
rect 42760 9568 42766 9580
rect 42981 9571 43039 9577
rect 42760 9540 42805 9568
rect 42760 9528 42766 9540
rect 42981 9537 42993 9571
rect 43027 9537 43039 9571
rect 43438 9568 43444 9580
rect 43399 9540 43444 9568
rect 42981 9531 43039 9537
rect 40052 9472 41736 9500
rect 42058 9460 42064 9512
rect 42116 9500 42122 9512
rect 42518 9500 42524 9512
rect 42116 9472 42524 9500
rect 42116 9460 42122 9472
rect 42518 9460 42524 9472
rect 42576 9500 42582 9512
rect 42889 9503 42947 9509
rect 42889 9500 42901 9503
rect 42576 9472 42901 9500
rect 42576 9460 42582 9472
rect 42889 9469 42901 9472
rect 42935 9469 42947 9503
rect 42889 9463 42947 9469
rect 35802 9432 35808 9444
rect 35176 9404 35808 9432
rect 35802 9392 35808 9404
rect 35860 9392 35866 9444
rect 38470 9392 38476 9444
rect 38528 9432 38534 9444
rect 39531 9435 39589 9441
rect 39531 9432 39543 9435
rect 38528 9404 39543 9432
rect 38528 9392 38534 9404
rect 39531 9401 39543 9404
rect 39577 9401 39589 9435
rect 39531 9395 39589 9401
rect 40218 9392 40224 9444
rect 40276 9432 40282 9444
rect 42996 9432 43024 9531
rect 43438 9528 43444 9540
rect 43496 9528 43502 9580
rect 43622 9568 43628 9580
rect 43583 9540 43628 9568
rect 43622 9528 43628 9540
rect 43680 9528 43686 9580
rect 43346 9432 43352 9444
rect 40276 9404 43352 9432
rect 40276 9392 40282 9404
rect 43346 9392 43352 9404
rect 43404 9392 43410 9444
rect 29880 9336 31754 9364
rect 32309 9367 32367 9373
rect 29880 9324 29886 9336
rect 32309 9333 32321 9367
rect 32355 9364 32367 9367
rect 34422 9364 34428 9376
rect 32355 9336 34428 9364
rect 32355 9333 32367 9336
rect 32309 9327 32367 9333
rect 34422 9324 34428 9336
rect 34480 9324 34486 9376
rect 34698 9364 34704 9376
rect 34659 9336 34704 9364
rect 34698 9324 34704 9336
rect 34756 9324 34762 9376
rect 34790 9324 34796 9376
rect 34848 9364 34854 9376
rect 35069 9367 35127 9373
rect 35069 9364 35081 9367
rect 34848 9336 35081 9364
rect 34848 9324 34854 9336
rect 35069 9333 35081 9336
rect 35115 9333 35127 9367
rect 35069 9327 35127 9333
rect 35897 9367 35955 9373
rect 35897 9333 35909 9367
rect 35943 9364 35955 9367
rect 40126 9364 40132 9376
rect 35943 9336 40132 9364
rect 35943 9333 35955 9336
rect 35897 9327 35955 9333
rect 40126 9324 40132 9336
rect 40184 9324 40190 9376
rect 40862 9324 40868 9376
rect 40920 9364 40926 9376
rect 41506 9364 41512 9376
rect 40920 9336 41512 9364
rect 40920 9324 40926 9336
rect 41506 9324 41512 9336
rect 41564 9324 41570 9376
rect 41690 9364 41696 9376
rect 41651 9336 41696 9364
rect 41690 9324 41696 9336
rect 41748 9324 41754 9376
rect 1104 9274 44896 9296
rect 1104 9222 6424 9274
rect 6476 9222 6488 9274
rect 6540 9222 6552 9274
rect 6604 9222 6616 9274
rect 6668 9222 6680 9274
rect 6732 9222 17372 9274
rect 17424 9222 17436 9274
rect 17488 9222 17500 9274
rect 17552 9222 17564 9274
rect 17616 9222 17628 9274
rect 17680 9222 28320 9274
rect 28372 9222 28384 9274
rect 28436 9222 28448 9274
rect 28500 9222 28512 9274
rect 28564 9222 28576 9274
rect 28628 9222 39268 9274
rect 39320 9222 39332 9274
rect 39384 9222 39396 9274
rect 39448 9222 39460 9274
rect 39512 9222 39524 9274
rect 39576 9222 44896 9274
rect 1104 9200 44896 9222
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 5718 9160 5724 9172
rect 3476 9132 5724 9160
rect 3476 9120 3482 9132
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 5813 9163 5871 9169
rect 5813 9129 5825 9163
rect 5859 9160 5871 9163
rect 6822 9160 6828 9172
rect 5859 9132 6828 9160
rect 5859 9129 5871 9132
rect 5813 9123 5871 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 11977 9163 12035 9169
rect 11977 9129 11989 9163
rect 12023 9160 12035 9163
rect 12434 9160 12440 9172
rect 12023 9132 12440 9160
rect 12023 9129 12035 9132
rect 11977 9123 12035 9129
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 27798 9160 27804 9172
rect 13044 9132 23796 9160
rect 27759 9132 27804 9160
rect 13044 9120 13050 9132
rect 4338 9092 4344 9104
rect 2884 9064 4344 9092
rect 2884 8965 2912 9064
rect 4338 9052 4344 9064
rect 4396 9052 4402 9104
rect 6270 9092 6276 9104
rect 6231 9064 6276 9092
rect 6270 9052 6276 9064
rect 6328 9052 6334 9104
rect 8202 9092 8208 9104
rect 6748 9064 8208 9092
rect 6748 9033 6776 9064
rect 8202 9052 8208 9064
rect 8260 9052 8266 9104
rect 17034 9092 17040 9104
rect 16995 9064 17040 9092
rect 17034 9052 17040 9064
rect 17092 9052 17098 9104
rect 21174 9092 21180 9104
rect 21135 9064 21180 9092
rect 21174 9052 21180 9064
rect 21232 9052 21238 9104
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 6733 9027 6791 9033
rect 3191 8996 4568 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 3970 8956 3976 8968
rect 3931 8928 3976 8956
rect 2869 8919 2927 8925
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4433 8959 4491 8965
rect 4433 8956 4445 8959
rect 4212 8928 4445 8956
rect 4212 8916 4218 8928
rect 4433 8925 4445 8928
rect 4479 8925 4491 8959
rect 4540 8956 4568 8996
rect 6733 8993 6745 9027
rect 6779 8993 6791 9027
rect 6733 8987 6791 8993
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 9024 6883 9027
rect 6914 9024 6920 9036
rect 6871 8996 6920 9024
rect 6871 8993 6883 8996
rect 6825 8987 6883 8993
rect 4540 8928 5028 8956
rect 4433 8919 4491 8925
rect 2774 8888 2780 8900
rect 2516 8860 2780 8888
rect 2516 8829 2544 8860
rect 2774 8848 2780 8860
rect 2832 8848 2838 8900
rect 4678 8891 4736 8897
rect 4678 8888 4690 8891
rect 4448 8860 4690 8888
rect 2501 8823 2559 8829
rect 2501 8789 2513 8823
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 2961 8823 3019 8829
rect 2961 8789 2973 8823
rect 3007 8820 3019 8823
rect 3050 8820 3056 8832
rect 3007 8792 3056 8820
rect 3007 8789 3019 8792
rect 2961 8783 3019 8789
rect 3050 8780 3056 8792
rect 3108 8780 3114 8832
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8820 3847 8823
rect 4448 8820 4476 8860
rect 4678 8857 4690 8860
rect 4724 8857 4736 8891
rect 5000 8888 5028 8928
rect 5074 8916 5080 8968
rect 5132 8956 5138 8968
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 5132 8928 6653 8956
rect 5132 8916 5138 8928
rect 6641 8925 6653 8928
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 6840 8888 6868 8987
rect 6914 8984 6920 8996
rect 6972 8984 6978 9036
rect 7282 8984 7288 9036
rect 7340 9024 7346 9036
rect 9125 9027 9183 9033
rect 9125 9024 9137 9027
rect 7340 8996 9137 9024
rect 7340 8984 7346 8996
rect 9125 8993 9137 8996
rect 9171 9024 9183 9027
rect 10502 9024 10508 9036
rect 9171 8996 10508 9024
rect 9171 8993 9183 8996
rect 9125 8987 9183 8993
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 13449 9027 13507 9033
rect 13449 8993 13461 9027
rect 13495 9024 13507 9027
rect 14642 9024 14648 9036
rect 13495 8996 14648 9024
rect 13495 8993 13507 8996
rect 13449 8987 13507 8993
rect 14642 8984 14648 8996
rect 14700 8984 14706 9036
rect 14734 8984 14740 9036
rect 14792 9024 14798 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 14792 8996 15301 9024
rect 14792 8984 14798 8996
rect 15289 8993 15301 8996
rect 15335 9024 15347 9027
rect 19702 9024 19708 9036
rect 15335 8996 18092 9024
rect 19663 8996 19708 9024
rect 15335 8993 15347 8996
rect 15289 8987 15347 8993
rect 18064 8968 18092 8996
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 20714 8984 20720 9036
rect 20772 9024 20778 9036
rect 23768 9024 23796 9132
rect 27798 9120 27804 9132
rect 27856 9120 27862 9172
rect 30374 9160 30380 9172
rect 30335 9132 30380 9160
rect 30374 9120 30380 9132
rect 30432 9120 30438 9172
rect 32766 9120 32772 9172
rect 32824 9160 32830 9172
rect 35066 9160 35072 9172
rect 32824 9132 34744 9160
rect 35027 9132 35072 9160
rect 32824 9120 32830 9132
rect 31570 9092 31576 9104
rect 30576 9064 31576 9092
rect 23845 9027 23903 9033
rect 23845 9024 23857 9027
rect 20772 8996 20944 9024
rect 23768 8996 23857 9024
rect 20772 8984 20778 8996
rect 7650 8956 7656 8968
rect 7611 8928 7656 8956
rect 7650 8916 7656 8928
rect 7708 8916 7714 8968
rect 7834 8956 7840 8968
rect 7795 8928 7840 8956
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 5000 8860 6868 8888
rect 4678 8851 4736 8857
rect 7466 8848 7472 8900
rect 7524 8888 7530 8900
rect 9416 8888 9444 8919
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 10597 8959 10655 8965
rect 10597 8956 10609 8959
rect 9732 8928 10609 8956
rect 9732 8916 9738 8928
rect 10597 8925 10609 8928
rect 10643 8956 10655 8959
rect 11698 8956 11704 8968
rect 10643 8928 11704 8956
rect 10643 8925 10655 8928
rect 10597 8919 10655 8925
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 13078 8916 13084 8968
rect 13136 8956 13142 8968
rect 13173 8959 13231 8965
rect 13173 8956 13185 8959
rect 13136 8928 13185 8956
rect 13136 8916 13142 8928
rect 13173 8925 13185 8928
rect 13219 8956 13231 8959
rect 14553 8959 14611 8965
rect 14553 8956 14565 8959
rect 13219 8928 14565 8956
rect 13219 8925 13231 8928
rect 13173 8919 13231 8925
rect 14553 8925 14565 8928
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 16666 8916 16672 8968
rect 16724 8916 16730 8968
rect 18046 8916 18052 8968
rect 18104 8956 18110 8968
rect 19242 8956 19248 8968
rect 18104 8928 19248 8956
rect 18104 8916 18110 8928
rect 19242 8916 19248 8928
rect 19300 8956 19306 8968
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19300 8928 19441 8956
rect 19300 8916 19306 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 20916 8956 20944 8996
rect 23845 8993 23857 8996
rect 23891 9024 23903 9027
rect 28718 9024 28724 9036
rect 23891 8996 28724 9024
rect 23891 8993 23903 8996
rect 23845 8987 23903 8993
rect 28718 8984 28724 8996
rect 28776 8984 28782 9036
rect 28828 8996 30052 9024
rect 24397 8959 24455 8965
rect 24397 8956 24409 8959
rect 20916 8928 24409 8956
rect 19429 8919 19487 8925
rect 24397 8925 24409 8928
rect 24443 8925 24455 8959
rect 24578 8956 24584 8968
rect 24539 8928 24584 8956
rect 24397 8919 24455 8925
rect 10410 8888 10416 8900
rect 7524 8860 10416 8888
rect 7524 8848 7530 8860
rect 10410 8848 10416 8860
rect 10468 8848 10474 8900
rect 10870 8897 10876 8900
rect 10864 8851 10876 8897
rect 10928 8888 10934 8900
rect 14461 8891 14519 8897
rect 10928 8860 10964 8888
rect 10870 8848 10876 8851
rect 10928 8848 10934 8860
rect 14461 8857 14473 8891
rect 14507 8888 14519 8891
rect 15286 8888 15292 8900
rect 14507 8860 15292 8888
rect 14507 8857 14519 8860
rect 14461 8851 14519 8857
rect 15286 8848 15292 8860
rect 15344 8848 15350 8900
rect 15562 8888 15568 8900
rect 15523 8860 15568 8888
rect 15562 8848 15568 8860
rect 15620 8848 15626 8900
rect 20930 8860 21312 8888
rect 3835 8792 4476 8820
rect 8021 8823 8079 8829
rect 3835 8789 3847 8792
rect 3789 8783 3847 8789
rect 8021 8789 8033 8823
rect 8067 8820 8079 8823
rect 8754 8820 8760 8832
rect 8067 8792 8760 8820
rect 8067 8789 8079 8792
rect 8021 8783 8079 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 12802 8820 12808 8832
rect 12763 8792 12808 8820
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 13262 8820 13268 8832
rect 13223 8792 13268 8820
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 14093 8823 14151 8829
rect 14093 8789 14105 8823
rect 14139 8820 14151 8823
rect 15470 8820 15476 8832
rect 14139 8792 15476 8820
rect 14139 8789 14151 8792
rect 14093 8783 14151 8789
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 21284 8820 21312 8860
rect 22094 8848 22100 8900
rect 22152 8888 22158 8900
rect 22152 8860 22197 8888
rect 22152 8848 22158 8860
rect 22738 8820 22744 8832
rect 21284 8792 22744 8820
rect 22738 8780 22744 8792
rect 22796 8780 22802 8832
rect 24412 8820 24440 8919
rect 24578 8916 24584 8928
rect 24636 8916 24642 8968
rect 24765 8959 24823 8965
rect 24765 8925 24777 8959
rect 24811 8956 24823 8959
rect 25409 8959 25467 8965
rect 25409 8956 25421 8959
rect 24811 8928 25421 8956
rect 24811 8925 24823 8928
rect 24765 8919 24823 8925
rect 25409 8925 25421 8928
rect 25455 8925 25467 8959
rect 25409 8919 25467 8925
rect 26053 8959 26111 8965
rect 26053 8925 26065 8959
rect 26099 8925 26111 8959
rect 26053 8919 26111 8925
rect 24486 8848 24492 8900
rect 24544 8888 24550 8900
rect 26068 8888 26096 8919
rect 27430 8916 27436 8968
rect 27488 8916 27494 8968
rect 27614 8916 27620 8968
rect 27672 8956 27678 8968
rect 28442 8956 28448 8968
rect 27672 8928 28448 8956
rect 27672 8916 27678 8928
rect 28442 8916 28448 8928
rect 28500 8956 28506 8968
rect 28828 8965 28856 8996
rect 28813 8959 28871 8965
rect 28813 8956 28825 8959
rect 28500 8928 28825 8956
rect 28500 8916 28506 8928
rect 28813 8925 28825 8928
rect 28859 8925 28871 8959
rect 28813 8919 28871 8925
rect 28997 8959 29055 8965
rect 28997 8925 29009 8959
rect 29043 8925 29055 8959
rect 28997 8919 29055 8925
rect 29733 8959 29791 8965
rect 29733 8925 29745 8959
rect 29779 8956 29791 8959
rect 29822 8956 29828 8968
rect 29779 8928 29828 8956
rect 29779 8925 29791 8928
rect 29733 8919 29791 8925
rect 26234 8888 26240 8900
rect 24544 8860 26240 8888
rect 24544 8848 24550 8860
rect 26234 8848 26240 8860
rect 26292 8848 26298 8900
rect 26326 8848 26332 8900
rect 26384 8888 26390 8900
rect 29012 8888 29040 8919
rect 29822 8916 29828 8928
rect 29880 8916 29886 8968
rect 29546 8888 29552 8900
rect 26384 8860 26429 8888
rect 27632 8860 29552 8888
rect 26384 8848 26390 8860
rect 27632 8832 27660 8860
rect 29546 8848 29552 8860
rect 29604 8848 29610 8900
rect 30024 8888 30052 8996
rect 30576 8965 30604 9064
rect 31570 9052 31576 9064
rect 31628 9052 31634 9104
rect 31662 9052 31668 9104
rect 31720 9092 31726 9104
rect 31757 9095 31815 9101
rect 31757 9092 31769 9095
rect 31720 9064 31769 9092
rect 31720 9052 31726 9064
rect 31757 9061 31769 9064
rect 31803 9061 31815 9095
rect 31757 9055 31815 9061
rect 30653 9027 30711 9033
rect 30653 8993 30665 9027
rect 30699 9024 30711 9027
rect 31849 9027 31907 9033
rect 31849 9024 31861 9027
rect 30699 8996 31861 9024
rect 30699 8993 30711 8996
rect 30653 8987 30711 8993
rect 31849 8993 31861 8996
rect 31895 9024 31907 9027
rect 31938 9024 31944 9036
rect 31895 8996 31944 9024
rect 31895 8993 31907 8996
rect 31849 8987 31907 8993
rect 31938 8984 31944 8996
rect 31996 8984 32002 9036
rect 32306 8984 32312 9036
rect 32364 9024 32370 9036
rect 32769 9027 32827 9033
rect 32769 9024 32781 9027
rect 32364 8996 32781 9024
rect 32364 8984 32370 8996
rect 32769 8993 32781 8996
rect 32815 8993 32827 9027
rect 34716 9024 34744 9132
rect 35066 9120 35072 9132
rect 35124 9120 35130 9172
rect 37369 9163 37427 9169
rect 37369 9129 37381 9163
rect 37415 9160 37427 9163
rect 38194 9160 38200 9172
rect 37415 9132 38200 9160
rect 37415 9129 37427 9132
rect 37369 9123 37427 9129
rect 38194 9120 38200 9132
rect 38252 9120 38258 9172
rect 38838 9160 38844 9172
rect 38799 9132 38844 9160
rect 38838 9120 38844 9132
rect 38896 9120 38902 9172
rect 40126 9120 40132 9172
rect 40184 9160 40190 9172
rect 40221 9163 40279 9169
rect 40221 9160 40233 9163
rect 40184 9132 40233 9160
rect 40184 9120 40190 9132
rect 40221 9129 40233 9132
rect 40267 9160 40279 9163
rect 42981 9163 43039 9169
rect 42981 9160 42993 9163
rect 40267 9132 42993 9160
rect 40267 9129 40279 9132
rect 40221 9123 40279 9129
rect 42981 9129 42993 9132
rect 43027 9129 43039 9163
rect 42981 9123 43039 9129
rect 43346 9120 43352 9172
rect 43404 9160 43410 9172
rect 43441 9163 43499 9169
rect 43441 9160 43453 9163
rect 43404 9132 43453 9160
rect 43404 9120 43410 9132
rect 43441 9129 43453 9132
rect 43487 9129 43499 9163
rect 43441 9123 43499 9129
rect 34882 9052 34888 9104
rect 34940 9092 34946 9104
rect 38381 9095 38439 9101
rect 34940 9064 38332 9092
rect 34940 9052 34946 9064
rect 34974 9024 34980 9036
rect 34716 8996 34980 9024
rect 32769 8987 32827 8993
rect 34974 8984 34980 8996
rect 35032 9024 35038 9036
rect 35161 9027 35219 9033
rect 35161 9024 35173 9027
rect 35032 8996 35173 9024
rect 35032 8984 35038 8996
rect 35161 8993 35173 8996
rect 35207 9024 35219 9027
rect 35894 9024 35900 9036
rect 35207 8996 35900 9024
rect 35207 8993 35219 8996
rect 35161 8987 35219 8993
rect 35894 8984 35900 8996
rect 35952 8984 35958 9036
rect 38304 9024 38332 9064
rect 38381 9061 38393 9095
rect 38427 9092 38439 9095
rect 39114 9092 39120 9104
rect 38427 9064 39120 9092
rect 38427 9061 38439 9064
rect 38381 9055 38439 9061
rect 39114 9052 39120 9064
rect 39172 9092 39178 9104
rect 39209 9095 39267 9101
rect 39209 9092 39221 9095
rect 39172 9064 39221 9092
rect 39172 9052 39178 9064
rect 39209 9061 39221 9064
rect 39255 9061 39267 9095
rect 39209 9055 39267 9061
rect 39850 9052 39856 9104
rect 39908 9092 39914 9104
rect 42150 9092 42156 9104
rect 39908 9064 40816 9092
rect 39908 9052 39914 9064
rect 39574 9024 39580 9036
rect 38304 8996 39580 9024
rect 39574 8984 39580 8996
rect 39632 8984 39638 9036
rect 40788 9033 40816 9064
rect 41984 9064 42156 9092
rect 40773 9027 40831 9033
rect 40773 8993 40785 9027
rect 40819 8993 40831 9027
rect 40773 8987 40831 8993
rect 30561 8959 30619 8965
rect 30561 8925 30573 8959
rect 30607 8925 30619 8959
rect 30742 8956 30748 8968
rect 30703 8928 30748 8956
rect 30561 8919 30619 8925
rect 30742 8916 30748 8928
rect 30800 8916 30806 8968
rect 30837 8959 30895 8965
rect 30837 8925 30849 8959
rect 30883 8956 30895 8959
rect 31478 8956 31484 8968
rect 30883 8928 31484 8956
rect 30883 8925 30895 8928
rect 30837 8919 30895 8925
rect 31478 8916 31484 8928
rect 31536 8916 31542 8968
rect 31570 8916 31576 8968
rect 31628 8956 31634 8968
rect 33036 8959 33094 8965
rect 31628 8928 31673 8956
rect 31628 8916 31634 8928
rect 33036 8925 33048 8959
rect 33082 8956 33094 8959
rect 34698 8956 34704 8968
rect 33082 8928 34704 8956
rect 33082 8925 33094 8928
rect 33036 8919 33094 8925
rect 34698 8916 34704 8928
rect 34756 8916 34762 8968
rect 34882 8956 34888 8968
rect 34843 8928 34888 8956
rect 34882 8916 34888 8928
rect 34940 8916 34946 8968
rect 37553 8959 37611 8965
rect 37553 8925 37565 8959
rect 37599 8956 37611 8959
rect 38562 8956 38568 8968
rect 37599 8928 38568 8956
rect 37599 8925 37611 8928
rect 37553 8919 37611 8925
rect 30760 8888 30788 8916
rect 30024 8860 30788 8888
rect 31389 8891 31447 8897
rect 31389 8857 31401 8891
rect 31435 8888 31447 8891
rect 33686 8888 33692 8900
rect 31435 8860 33692 8888
rect 31435 8857 31447 8860
rect 31389 8851 31447 8857
rect 33686 8848 33692 8860
rect 33744 8848 33750 8900
rect 34422 8848 34428 8900
rect 34480 8888 34486 8900
rect 37559 8888 37587 8919
rect 38562 8916 38568 8928
rect 38620 8916 38626 8968
rect 39022 8956 39028 8968
rect 38983 8928 39028 8956
rect 39022 8916 39028 8928
rect 39080 8916 39086 8968
rect 39301 8959 39359 8965
rect 39301 8925 39313 8959
rect 39347 8956 39359 8959
rect 39666 8956 39672 8968
rect 39347 8928 39672 8956
rect 39347 8925 39359 8928
rect 39301 8919 39359 8925
rect 39666 8916 39672 8928
rect 39724 8916 39730 8968
rect 40034 8956 40040 8968
rect 39995 8928 40040 8956
rect 40034 8916 40040 8928
rect 40092 8916 40098 8968
rect 40313 8959 40371 8965
rect 40313 8925 40325 8959
rect 40359 8925 40371 8959
rect 40313 8919 40371 8925
rect 34480 8860 37587 8888
rect 38013 8891 38071 8897
rect 34480 8848 34486 8860
rect 38013 8857 38025 8891
rect 38059 8857 38071 8891
rect 38013 8851 38071 8857
rect 38229 8891 38287 8897
rect 38229 8857 38241 8891
rect 38275 8888 38287 8891
rect 38654 8888 38660 8900
rect 38275 8860 38660 8888
rect 38275 8857 38287 8860
rect 38229 8851 38287 8857
rect 25038 8820 25044 8832
rect 24412 8792 25044 8820
rect 25038 8780 25044 8792
rect 25096 8780 25102 8832
rect 25222 8820 25228 8832
rect 25183 8792 25228 8820
rect 25222 8780 25228 8792
rect 25280 8780 25286 8832
rect 26694 8780 26700 8832
rect 26752 8820 26758 8832
rect 27614 8820 27620 8832
rect 26752 8792 27620 8820
rect 26752 8780 26758 8792
rect 27614 8780 27620 8792
rect 27672 8780 27678 8832
rect 28902 8820 28908 8832
rect 28863 8792 28908 8820
rect 28902 8780 28908 8792
rect 28960 8780 28966 8832
rect 28994 8780 29000 8832
rect 29052 8820 29058 8832
rect 29825 8823 29883 8829
rect 29825 8820 29837 8823
rect 29052 8792 29837 8820
rect 29052 8780 29058 8792
rect 29825 8789 29837 8792
rect 29871 8820 29883 8823
rect 31662 8820 31668 8832
rect 29871 8792 31668 8820
rect 29871 8789 29883 8792
rect 29825 8783 29883 8789
rect 31662 8780 31668 8792
rect 31720 8780 31726 8832
rect 32674 8780 32680 8832
rect 32732 8820 32738 8832
rect 34149 8823 34207 8829
rect 34149 8820 34161 8823
rect 32732 8792 34161 8820
rect 32732 8780 32738 8792
rect 34149 8789 34161 8792
rect 34195 8820 34207 8823
rect 34514 8820 34520 8832
rect 34195 8792 34520 8820
rect 34195 8789 34207 8792
rect 34149 8783 34207 8789
rect 34514 8780 34520 8792
rect 34572 8780 34578 8832
rect 34698 8820 34704 8832
rect 34659 8792 34704 8820
rect 34698 8780 34704 8792
rect 34756 8780 34762 8832
rect 38028 8820 38056 8851
rect 38654 8848 38660 8860
rect 38712 8888 38718 8900
rect 38712 8860 39988 8888
rect 38712 8848 38718 8860
rect 39206 8820 39212 8832
rect 38028 8792 39212 8820
rect 39206 8780 39212 8792
rect 39264 8780 39270 8832
rect 39298 8780 39304 8832
rect 39356 8820 39362 8832
rect 39853 8823 39911 8829
rect 39853 8820 39865 8823
rect 39356 8792 39865 8820
rect 39356 8780 39362 8792
rect 39853 8789 39865 8792
rect 39899 8789 39911 8823
rect 39960 8820 39988 8860
rect 40218 8848 40224 8900
rect 40276 8888 40282 8900
rect 40328 8888 40356 8919
rect 40494 8916 40500 8968
rect 40552 8956 40558 8968
rect 40552 8928 41414 8956
rect 40552 8916 40558 8928
rect 40276 8860 40356 8888
rect 40276 8848 40282 8860
rect 40770 8848 40776 8900
rect 40828 8888 40834 8900
rect 41018 8891 41076 8897
rect 41018 8888 41030 8891
rect 40828 8860 41030 8888
rect 40828 8848 40834 8860
rect 41018 8857 41030 8860
rect 41064 8857 41076 8891
rect 41386 8888 41414 8928
rect 41506 8916 41512 8968
rect 41564 8956 41570 8968
rect 41984 8956 42012 9064
rect 42150 9052 42156 9064
rect 42208 9052 42214 9104
rect 41564 8928 42012 8956
rect 42076 8996 43668 9024
rect 41564 8916 41570 8928
rect 42076 8888 42104 8996
rect 42610 8956 42616 8968
rect 42571 8928 42616 8956
rect 42610 8916 42616 8928
rect 42668 8916 42674 8968
rect 43640 8965 43668 8996
rect 42797 8959 42855 8965
rect 42797 8956 42809 8959
rect 42720 8928 42809 8956
rect 41386 8860 42104 8888
rect 41018 8851 41076 8857
rect 42720 8820 42748 8928
rect 42797 8925 42809 8928
rect 42843 8925 42855 8959
rect 42797 8919 42855 8925
rect 43625 8959 43683 8965
rect 43625 8925 43637 8959
rect 43671 8925 43683 8959
rect 43625 8919 43683 8925
rect 42794 8820 42800 8832
rect 39960 8792 42800 8820
rect 39853 8783 39911 8789
rect 42794 8780 42800 8792
rect 42852 8780 42858 8832
rect 1104 8730 45056 8752
rect 1104 8678 11898 8730
rect 11950 8678 11962 8730
rect 12014 8678 12026 8730
rect 12078 8678 12090 8730
rect 12142 8678 12154 8730
rect 12206 8678 22846 8730
rect 22898 8678 22910 8730
rect 22962 8678 22974 8730
rect 23026 8678 23038 8730
rect 23090 8678 23102 8730
rect 23154 8678 33794 8730
rect 33846 8678 33858 8730
rect 33910 8678 33922 8730
rect 33974 8678 33986 8730
rect 34038 8678 34050 8730
rect 34102 8678 44742 8730
rect 44794 8678 44806 8730
rect 44858 8678 44870 8730
rect 44922 8678 44934 8730
rect 44986 8678 44998 8730
rect 45050 8678 45056 8730
rect 1104 8656 45056 8678
rect 1397 8619 1455 8625
rect 1397 8585 1409 8619
rect 1443 8585 1455 8619
rect 3050 8616 3056 8628
rect 3011 8588 3056 8616
rect 1397 8579 1455 8585
rect 1412 8548 1440 8579
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 3142 8576 3148 8628
rect 3200 8616 3206 8628
rect 4890 8616 4896 8628
rect 3200 8588 4896 8616
rect 3200 8576 3206 8588
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 7515 8619 7573 8625
rect 7515 8585 7527 8619
rect 7561 8616 7573 8619
rect 7650 8616 7656 8628
rect 7561 8588 7656 8616
rect 7561 8585 7573 8588
rect 7515 8579 7573 8585
rect 7650 8576 7656 8588
rect 7708 8616 7714 8628
rect 9858 8616 9864 8628
rect 7708 8588 9864 8616
rect 7708 8576 7714 8588
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10594 8616 10600 8628
rect 10555 8588 10600 8616
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 13078 8616 13084 8628
rect 13039 8588 13084 8616
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 13538 8616 13544 8628
rect 13499 8588 13544 8616
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 13909 8619 13967 8625
rect 13909 8585 13921 8619
rect 13955 8616 13967 8619
rect 13955 8588 15792 8616
rect 13955 8585 13967 8588
rect 13909 8579 13967 8585
rect 14001 8551 14059 8557
rect 14001 8548 14013 8551
rect 1412 8520 14013 8548
rect 14001 8517 14013 8520
rect 14047 8517 14059 8551
rect 14001 8511 14059 8517
rect 1578 8480 1584 8492
rect 1539 8452 1584 8480
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8480 2559 8483
rect 3142 8480 3148 8492
rect 2547 8452 3148 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3234 8440 3240 8492
rect 3292 8480 3298 8492
rect 3769 8483 3827 8489
rect 3769 8480 3781 8483
rect 3292 8452 3781 8480
rect 3292 8440 3298 8452
rect 3769 8449 3781 8452
rect 3815 8449 3827 8483
rect 3769 8443 3827 8449
rect 4338 8440 4344 8492
rect 4396 8480 4402 8492
rect 5350 8480 5356 8492
rect 4396 8452 5356 8480
rect 4396 8440 4402 8452
rect 5350 8440 5356 8452
rect 5408 8480 5414 8492
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 5408 8452 5641 8480
rect 5408 8440 5414 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 6822 8480 6828 8492
rect 6595 8452 6828 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 7282 8480 7288 8492
rect 7243 8452 7288 8480
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 8754 8480 8760 8492
rect 8715 8452 8760 8480
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 9214 8480 9220 8492
rect 9175 8452 9220 8480
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 9473 8483 9531 8489
rect 9473 8480 9485 8483
rect 9364 8452 9485 8480
rect 9364 8440 9370 8452
rect 9473 8449 9485 8452
rect 9519 8449 9531 8483
rect 11698 8480 11704 8492
rect 11659 8452 11704 8480
rect 9473 8443 9531 8449
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 11957 8483 12015 8489
rect 11957 8480 11969 8483
rect 11848 8452 11969 8480
rect 11848 8440 11854 8452
rect 11957 8449 11969 8452
rect 12003 8449 12015 8483
rect 14734 8480 14740 8492
rect 14695 8452 14740 8480
rect 11957 8443 12015 8449
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 15004 8483 15062 8489
rect 15004 8449 15016 8483
rect 15050 8480 15062 8483
rect 15286 8480 15292 8492
rect 15050 8452 15292 8480
rect 15050 8449 15062 8452
rect 15004 8443 15062 8449
rect 15286 8440 15292 8452
rect 15344 8480 15350 8492
rect 15562 8480 15568 8492
rect 15344 8452 15568 8480
rect 15344 8440 15350 8452
rect 15562 8440 15568 8452
rect 15620 8440 15626 8492
rect 15764 8480 15792 8588
rect 15838 8576 15844 8628
rect 15896 8616 15902 8628
rect 16117 8619 16175 8625
rect 16117 8616 16129 8619
rect 15896 8588 16129 8616
rect 15896 8576 15902 8588
rect 16117 8585 16129 8588
rect 16163 8585 16175 8619
rect 19426 8616 19432 8628
rect 19387 8588 19432 8616
rect 16117 8579 16175 8585
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 25590 8616 25596 8628
rect 22020 8588 25596 8616
rect 16482 8508 16488 8560
rect 16540 8548 16546 8560
rect 22020 8548 22048 8588
rect 25590 8576 25596 8588
rect 25648 8576 25654 8628
rect 25869 8619 25927 8625
rect 25869 8585 25881 8619
rect 25915 8616 25927 8619
rect 27433 8619 27491 8625
rect 27433 8616 27445 8619
rect 25915 8588 27445 8616
rect 25915 8585 25927 8588
rect 25869 8579 25927 8585
rect 27433 8585 27445 8588
rect 27479 8585 27491 8619
rect 27433 8579 27491 8585
rect 27540 8588 32444 8616
rect 16540 8520 22048 8548
rect 22097 8551 22155 8557
rect 16540 8508 16546 8520
rect 22097 8517 22109 8551
rect 22143 8548 22155 8551
rect 22370 8548 22376 8560
rect 22143 8520 22376 8548
rect 22143 8517 22155 8520
rect 22097 8511 22155 8517
rect 22370 8508 22376 8520
rect 22428 8508 22434 8560
rect 27540 8548 27568 8588
rect 23616 8520 27568 8548
rect 17954 8480 17960 8492
rect 15764 8452 17960 8480
rect 17954 8440 17960 8452
rect 18012 8480 18018 8492
rect 18305 8483 18363 8489
rect 18305 8480 18317 8483
rect 18012 8452 18317 8480
rect 18012 8440 18018 8452
rect 18305 8449 18317 8452
rect 18351 8449 18363 8483
rect 18305 8443 18363 8449
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8480 20315 8483
rect 21082 8480 21088 8492
rect 20303 8452 21088 8480
rect 20303 8449 20315 8452
rect 20257 8443 20315 8449
rect 21082 8440 21088 8452
rect 21140 8440 21146 8492
rect 21266 8480 21272 8492
rect 21227 8452 21272 8480
rect 21266 8440 21272 8452
rect 21324 8440 21330 8492
rect 23198 8440 23204 8492
rect 23256 8440 23262 8492
rect 3510 8412 3516 8424
rect 3471 8384 3516 8412
rect 3510 8372 3516 8384
rect 3568 8372 3574 8424
rect 4982 8372 4988 8424
rect 5040 8412 5046 8424
rect 5445 8415 5503 8421
rect 5445 8412 5457 8415
rect 5040 8384 5457 8412
rect 5040 8372 5046 8384
rect 5445 8381 5457 8384
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8412 6423 8415
rect 7466 8412 7472 8424
rect 6411 8384 7472 8412
rect 6411 8381 6423 8384
rect 6365 8375 6423 8381
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 14182 8412 14188 8424
rect 14143 8384 14188 8412
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 18046 8412 18052 8424
rect 18007 8384 18052 8412
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 20346 8412 20352 8424
rect 20307 8384 20352 8412
rect 20346 8372 20352 8384
rect 20404 8372 20410 8424
rect 20438 8372 20444 8424
rect 20496 8421 20502 8424
rect 20496 8415 20545 8421
rect 20496 8381 20499 8415
rect 20533 8381 20545 8415
rect 21818 8412 21824 8424
rect 21779 8384 21824 8412
rect 20496 8375 20545 8381
rect 20496 8372 20502 8375
rect 21818 8372 21824 8384
rect 21876 8372 21882 8424
rect 23616 8421 23644 8520
rect 27706 8508 27712 8560
rect 27764 8548 27770 8560
rect 28261 8551 28319 8557
rect 28261 8548 28273 8551
rect 27764 8520 28273 8548
rect 27764 8508 27770 8520
rect 28261 8517 28273 8520
rect 28307 8517 28319 8551
rect 28442 8548 28448 8560
rect 28403 8520 28448 8548
rect 28261 8511 28319 8517
rect 28442 8508 28448 8520
rect 28500 8508 28506 8560
rect 28902 8508 28908 8560
rect 28960 8548 28966 8560
rect 28960 8520 30131 8548
rect 28960 8508 28966 8520
rect 24745 8483 24803 8489
rect 24745 8480 24757 8483
rect 23569 8415 23644 8421
rect 23569 8381 23581 8415
rect 23615 8384 23644 8415
rect 23676 8452 24757 8480
rect 23615 8381 23627 8384
rect 23569 8375 23627 8381
rect 5810 8344 5816 8356
rect 5771 8316 5816 8344
rect 5810 8304 5816 8316
rect 5868 8304 5874 8356
rect 6733 8347 6791 8353
rect 6733 8313 6745 8347
rect 6779 8344 6791 8347
rect 6822 8344 6828 8356
rect 6779 8316 6828 8344
rect 6779 8313 6791 8316
rect 6733 8307 6791 8313
rect 6822 8304 6828 8316
rect 6880 8304 6886 8356
rect 21085 8347 21143 8353
rect 19306 8316 20392 8344
rect 8570 8276 8576 8288
rect 8531 8248 8576 8276
rect 8570 8236 8576 8248
rect 8628 8236 8634 8288
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 13354 8276 13360 8288
rect 10836 8248 13360 8276
rect 10836 8236 10842 8248
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 19306 8276 19334 8316
rect 19886 8276 19892 8288
rect 13504 8248 19334 8276
rect 19847 8248 19892 8276
rect 13504 8236 13510 8248
rect 19886 8236 19892 8248
rect 19944 8236 19950 8288
rect 20364 8276 20392 8316
rect 21085 8313 21097 8347
rect 21131 8344 21143 8347
rect 23676 8344 23704 8452
rect 24745 8449 24757 8452
rect 24791 8449 24803 8483
rect 24745 8443 24803 8449
rect 25038 8440 25044 8492
rect 25096 8480 25102 8492
rect 27338 8480 27344 8492
rect 25096 8452 25544 8480
rect 27299 8452 27344 8480
rect 25096 8440 25102 8452
rect 24486 8412 24492 8424
rect 24447 8384 24492 8412
rect 24486 8372 24492 8384
rect 24544 8372 24550 8424
rect 21131 8316 21956 8344
rect 21131 8313 21143 8316
rect 21085 8307 21143 8313
rect 20438 8276 20444 8288
rect 20364 8248 20444 8276
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 21928 8276 21956 8316
rect 23124 8316 23704 8344
rect 25516 8344 25544 8452
rect 27338 8440 27344 8452
rect 27396 8440 27402 8492
rect 28994 8480 29000 8492
rect 27448 8452 29000 8480
rect 25590 8372 25596 8424
rect 25648 8412 25654 8424
rect 27448 8412 27476 8452
rect 28994 8440 29000 8452
rect 29052 8440 29058 8492
rect 29546 8440 29552 8492
rect 29604 8480 29610 8492
rect 29733 8483 29791 8489
rect 29733 8480 29745 8483
rect 29604 8452 29745 8480
rect 29604 8440 29610 8452
rect 29733 8449 29745 8452
rect 29779 8449 29791 8483
rect 29733 8443 29791 8449
rect 29822 8440 29828 8492
rect 29880 8489 29886 8492
rect 29880 8483 29929 8489
rect 29880 8449 29883 8483
rect 29917 8449 29929 8483
rect 30006 8480 30012 8492
rect 29967 8452 30012 8480
rect 29880 8443 29929 8449
rect 29880 8440 29886 8443
rect 30006 8440 30012 8452
rect 30064 8440 30070 8492
rect 30103 8489 30131 8520
rect 32416 8492 32444 8588
rect 33686 8576 33692 8628
rect 33744 8616 33750 8628
rect 34790 8616 34796 8628
rect 33744 8588 34796 8616
rect 33744 8576 33750 8588
rect 34790 8576 34796 8588
rect 34848 8576 34854 8628
rect 34882 8576 34888 8628
rect 34940 8616 34946 8628
rect 38473 8619 38531 8625
rect 38473 8616 38485 8619
rect 34940 8588 38485 8616
rect 34940 8576 34946 8588
rect 38473 8585 38485 8588
rect 38519 8585 38531 8619
rect 38473 8579 38531 8585
rect 38930 8576 38936 8628
rect 38988 8616 38994 8628
rect 40405 8619 40463 8625
rect 40405 8616 40417 8619
rect 38988 8588 40417 8616
rect 38988 8576 38994 8588
rect 40405 8585 40417 8588
rect 40451 8616 40463 8619
rect 40494 8616 40500 8628
rect 40451 8588 40500 8616
rect 40451 8585 40463 8588
rect 40405 8579 40463 8585
rect 40494 8576 40500 8588
rect 40552 8576 40558 8628
rect 43993 8619 44051 8625
rect 43993 8616 44005 8619
rect 41386 8588 44005 8616
rect 39850 8548 39856 8560
rect 33612 8520 39856 8548
rect 30103 8483 30183 8489
rect 30103 8450 30137 8483
rect 30125 8449 30137 8450
rect 30171 8449 30183 8483
rect 30125 8443 30183 8449
rect 31389 8483 31447 8489
rect 31389 8449 31401 8483
rect 31435 8480 31447 8483
rect 32122 8480 32128 8492
rect 31435 8452 32128 8480
rect 31435 8449 31447 8452
rect 31389 8443 31447 8449
rect 32122 8440 32128 8452
rect 32180 8440 32186 8492
rect 32398 8480 32404 8492
rect 32359 8452 32404 8480
rect 32398 8440 32404 8452
rect 32456 8440 32462 8492
rect 33042 8440 33048 8492
rect 33100 8480 33106 8492
rect 33612 8489 33640 8520
rect 33597 8483 33655 8489
rect 33597 8480 33609 8483
rect 33100 8452 33609 8480
rect 33100 8440 33106 8452
rect 33597 8449 33609 8452
rect 33643 8449 33655 8483
rect 33597 8443 33655 8449
rect 33864 8483 33922 8489
rect 33864 8449 33876 8483
rect 33910 8480 33922 8483
rect 34698 8480 34704 8492
rect 33910 8452 34704 8480
rect 33910 8449 33922 8452
rect 33864 8443 33922 8449
rect 34698 8440 34704 8452
rect 34756 8440 34762 8492
rect 37366 8480 37372 8492
rect 37327 8452 37372 8480
rect 37366 8440 37372 8452
rect 37424 8440 37430 8492
rect 38194 8440 38200 8492
rect 38252 8480 38258 8492
rect 38381 8483 38439 8489
rect 38381 8480 38393 8483
rect 38252 8452 38393 8480
rect 38252 8440 38258 8452
rect 38381 8449 38393 8452
rect 38427 8449 38439 8483
rect 38381 8443 38439 8449
rect 25648 8384 27476 8412
rect 25648 8372 25654 8384
rect 27522 8372 27528 8424
rect 27580 8412 27586 8424
rect 27580 8384 27625 8412
rect 27580 8372 27586 8384
rect 28810 8372 28816 8424
rect 28868 8412 28874 8424
rect 29181 8415 29239 8421
rect 29181 8412 29193 8415
rect 28868 8384 29193 8412
rect 28868 8372 28874 8384
rect 29181 8381 29193 8384
rect 29227 8381 29239 8415
rect 29181 8375 29239 8381
rect 31205 8415 31263 8421
rect 31205 8381 31217 8415
rect 31251 8381 31263 8415
rect 31205 8375 31263 8381
rect 32217 8415 32275 8421
rect 32217 8381 32229 8415
rect 32263 8412 32275 8415
rect 38396 8412 38424 8443
rect 38470 8440 38476 8492
rect 38528 8480 38534 8492
rect 38565 8483 38623 8489
rect 38565 8480 38577 8483
rect 38528 8452 38577 8480
rect 38528 8440 38534 8452
rect 38565 8449 38577 8452
rect 38611 8480 38623 8483
rect 38930 8480 38936 8492
rect 38611 8452 38936 8480
rect 38611 8449 38623 8452
rect 38565 8443 38623 8449
rect 38930 8440 38936 8452
rect 38988 8440 38994 8492
rect 39040 8489 39068 8520
rect 39850 8508 39856 8520
rect 39908 8508 39914 8560
rect 41386 8548 41414 8588
rect 43993 8585 44005 8588
rect 44039 8585 44051 8619
rect 43993 8579 44051 8585
rect 42794 8548 42800 8560
rect 39960 8520 41414 8548
rect 42755 8520 42800 8548
rect 39298 8489 39304 8492
rect 39025 8483 39083 8489
rect 39025 8449 39037 8483
rect 39071 8449 39083 8483
rect 39292 8480 39304 8489
rect 39259 8452 39304 8480
rect 39025 8443 39083 8449
rect 39292 8443 39304 8452
rect 39298 8440 39304 8443
rect 39356 8440 39362 8492
rect 39574 8440 39580 8492
rect 39632 8480 39638 8492
rect 39960 8480 39988 8520
rect 42794 8508 42800 8520
rect 42852 8508 42858 8560
rect 39632 8452 39988 8480
rect 40865 8483 40923 8489
rect 39632 8440 39638 8452
rect 40865 8449 40877 8483
rect 40911 8480 40923 8483
rect 41230 8480 41236 8492
rect 40911 8452 41236 8480
rect 40911 8449 40923 8452
rect 40865 8443 40923 8449
rect 41230 8440 41236 8452
rect 41288 8480 41294 8492
rect 42613 8483 42671 8489
rect 42613 8480 42625 8483
rect 41288 8452 42625 8480
rect 41288 8440 41294 8452
rect 42613 8449 42625 8452
rect 42659 8449 42671 8483
rect 43254 8480 43260 8492
rect 43215 8452 43260 8480
rect 42613 8443 42671 8449
rect 43254 8440 43260 8452
rect 43312 8440 43318 8492
rect 44174 8480 44180 8492
rect 44135 8452 44180 8480
rect 44174 8440 44180 8452
rect 44232 8440 44238 8492
rect 32263 8384 33640 8412
rect 38396 8384 39068 8412
rect 32263 8381 32275 8384
rect 32217 8375 32275 8381
rect 31220 8344 31248 8375
rect 25516 8316 31248 8344
rect 23124 8276 23152 8316
rect 31478 8304 31484 8356
rect 31536 8304 31542 8356
rect 31573 8347 31631 8353
rect 31573 8313 31585 8347
rect 31619 8344 31631 8347
rect 32490 8344 32496 8356
rect 31619 8316 32496 8344
rect 31619 8313 31631 8316
rect 31573 8307 31631 8313
rect 32490 8304 32496 8316
rect 32548 8304 32554 8356
rect 32585 8347 32643 8353
rect 32585 8313 32597 8347
rect 32631 8344 32643 8347
rect 33502 8344 33508 8356
rect 32631 8316 33508 8344
rect 32631 8313 32643 8316
rect 32585 8307 32643 8313
rect 33502 8304 33508 8316
rect 33560 8304 33566 8356
rect 26970 8276 26976 8288
rect 21928 8248 23152 8276
rect 26931 8248 26976 8276
rect 26970 8236 26976 8248
rect 27028 8236 27034 8288
rect 30282 8276 30288 8288
rect 30243 8248 30288 8276
rect 30282 8236 30288 8248
rect 30340 8236 30346 8288
rect 31496 8276 31524 8304
rect 32858 8276 32864 8288
rect 31496 8248 32864 8276
rect 32858 8236 32864 8248
rect 32916 8236 32922 8288
rect 33612 8276 33640 8384
rect 34974 8344 34980 8356
rect 34935 8316 34980 8344
rect 34974 8304 34980 8316
rect 35032 8304 35038 8356
rect 37461 8347 37519 8353
rect 37461 8313 37473 8347
rect 37507 8344 37519 8347
rect 38746 8344 38752 8356
rect 37507 8316 38752 8344
rect 37507 8313 37519 8316
rect 37461 8307 37519 8313
rect 38746 8304 38752 8316
rect 38804 8304 38810 8356
rect 34606 8276 34612 8288
rect 33612 8248 34612 8276
rect 34606 8236 34612 8248
rect 34664 8236 34670 8288
rect 39040 8276 39068 8384
rect 40402 8372 40408 8424
rect 40460 8412 40466 8424
rect 41138 8412 41144 8424
rect 40460 8384 41144 8412
rect 40460 8372 40466 8384
rect 41138 8372 41144 8384
rect 41196 8372 41202 8424
rect 41506 8372 41512 8424
rect 41564 8412 41570 8424
rect 42429 8415 42487 8421
rect 42429 8412 42441 8415
rect 41564 8384 42441 8412
rect 41564 8372 41570 8384
rect 42429 8381 42441 8384
rect 42475 8381 42487 8415
rect 42429 8375 42487 8381
rect 42518 8372 42524 8424
rect 42576 8412 42582 8424
rect 43349 8415 43407 8421
rect 43349 8412 43361 8415
rect 42576 8384 43361 8412
rect 42576 8372 42582 8384
rect 43349 8381 43361 8384
rect 43395 8381 43407 8415
rect 43349 8375 43407 8381
rect 42610 8344 42616 8356
rect 40052 8316 42616 8344
rect 40052 8276 40080 8316
rect 42610 8304 42616 8316
rect 42668 8304 42674 8356
rect 39040 8248 40080 8276
rect 1104 8186 44896 8208
rect 1104 8134 6424 8186
rect 6476 8134 6488 8186
rect 6540 8134 6552 8186
rect 6604 8134 6616 8186
rect 6668 8134 6680 8186
rect 6732 8134 17372 8186
rect 17424 8134 17436 8186
rect 17488 8134 17500 8186
rect 17552 8134 17564 8186
rect 17616 8134 17628 8186
rect 17680 8134 28320 8186
rect 28372 8134 28384 8186
rect 28436 8134 28448 8186
rect 28500 8134 28512 8186
rect 28564 8134 28576 8186
rect 28628 8134 39268 8186
rect 39320 8134 39332 8186
rect 39384 8134 39396 8186
rect 39448 8134 39460 8186
rect 39512 8134 39524 8186
rect 39576 8134 44896 8186
rect 1104 8112 44896 8134
rect 5350 8072 5356 8084
rect 5311 8044 5356 8072
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 7834 8072 7840 8084
rect 7795 8044 7840 8072
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 10781 8075 10839 8081
rect 10781 8041 10793 8075
rect 10827 8072 10839 8075
rect 10870 8072 10876 8084
rect 10827 8044 10876 8072
rect 10827 8041 10839 8044
rect 10781 8035 10839 8041
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 15562 8072 15568 8084
rect 13412 8044 15424 8072
rect 15523 8044 15568 8072
rect 13412 8032 13418 8044
rect 15396 8004 15424 8044
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 15930 8072 15936 8084
rect 15856 8044 15936 8072
rect 15856 8004 15884 8044
rect 15930 8032 15936 8044
rect 15988 8032 15994 8084
rect 18690 8032 18696 8084
rect 18748 8072 18754 8084
rect 19886 8072 19892 8084
rect 18748 8044 19892 8072
rect 18748 8032 18754 8044
rect 19886 8032 19892 8044
rect 19944 8032 19950 8084
rect 21082 8072 21088 8084
rect 21043 8044 21088 8072
rect 21082 8032 21088 8044
rect 21140 8032 21146 8084
rect 23382 8072 23388 8084
rect 22480 8044 23388 8072
rect 16022 8004 16028 8016
rect 15396 7976 15884 8004
rect 15983 7976 16028 8004
rect 16022 7964 16028 7976
rect 16080 7964 16086 8016
rect 16482 7964 16488 8016
rect 16540 7964 16546 8016
rect 21560 7976 21772 8004
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 11885 7939 11943 7945
rect 11885 7936 11897 7939
rect 11756 7908 11897 7936
rect 11756 7896 11762 7908
rect 11885 7905 11897 7908
rect 11931 7905 11943 7939
rect 16500 7936 16528 7964
rect 16577 7939 16635 7945
rect 16577 7936 16589 7939
rect 16500 7908 16589 7936
rect 11885 7899 11943 7905
rect 16577 7905 16589 7908
rect 16623 7905 16635 7939
rect 16577 7899 16635 7905
rect 17494 7896 17500 7948
rect 17552 7936 17558 7948
rect 17552 7908 19380 7936
rect 17552 7896 17558 7908
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4062 7868 4068 7880
rect 4019 7840 4068 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4062 7828 4068 7840
rect 4120 7868 4126 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 4120 7840 6469 7868
rect 4120 7828 4126 7840
rect 6457 7837 6469 7840
rect 6503 7868 6515 7871
rect 7006 7868 7012 7880
rect 6503 7840 7012 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 7006 7828 7012 7840
rect 7064 7868 7070 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 7064 7840 8953 7868
rect 7064 7828 7070 7840
rect 8941 7837 8953 7840
rect 8987 7868 8999 7871
rect 9674 7868 9680 7880
rect 8987 7840 9680 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7868 11023 7871
rect 11514 7868 11520 7880
rect 11011 7840 11520 7868
rect 11011 7837 11023 7840
rect 10965 7831 11023 7837
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 13354 7828 13360 7880
rect 13412 7868 13418 7880
rect 14185 7871 14243 7877
rect 14185 7868 14197 7871
rect 13412 7840 14197 7868
rect 13412 7828 13418 7840
rect 14185 7837 14197 7840
rect 14231 7868 14243 7871
rect 14734 7868 14740 7880
rect 14231 7840 14740 7868
rect 14231 7837 14243 7840
rect 14185 7831 14243 7837
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 15378 7828 15384 7880
rect 15436 7868 15442 7880
rect 16485 7871 16543 7877
rect 16485 7868 16497 7871
rect 15436 7840 16497 7868
rect 15436 7828 15442 7840
rect 16485 7837 16497 7840
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 16666 7828 16672 7880
rect 16724 7868 16730 7880
rect 17405 7871 17463 7877
rect 17405 7868 17417 7871
rect 16724 7840 17417 7868
rect 16724 7828 16730 7840
rect 17405 7837 17417 7840
rect 17451 7837 17463 7871
rect 18690 7868 18696 7880
rect 18651 7840 18696 7868
rect 17405 7831 17463 7837
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 19242 7868 19248 7880
rect 19203 7840 19248 7868
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 19352 7868 19380 7908
rect 21560 7868 21588 7976
rect 21744 7945 21772 7976
rect 21729 7939 21787 7945
rect 21729 7905 21741 7939
rect 21775 7936 21787 7939
rect 22370 7936 22376 7948
rect 21775 7908 22376 7936
rect 21775 7905 21787 7908
rect 21729 7899 21787 7905
rect 22370 7896 22376 7908
rect 22428 7896 22434 7948
rect 19352 7840 21588 7868
rect 22278 7828 22284 7880
rect 22336 7868 22342 7880
rect 22480 7877 22508 8044
rect 23382 8032 23388 8044
rect 23440 8072 23446 8084
rect 23845 8075 23903 8081
rect 23440 8044 23796 8072
rect 23440 8032 23446 8044
rect 22465 7871 22523 7877
rect 22465 7868 22477 7871
rect 22336 7840 22477 7868
rect 22336 7828 22342 7840
rect 22465 7837 22477 7840
rect 22511 7837 22523 7871
rect 22732 7871 22790 7877
rect 22732 7868 22744 7871
rect 22465 7831 22523 7837
rect 22664 7840 22744 7868
rect 22664 7812 22692 7840
rect 22732 7837 22744 7840
rect 22778 7837 22790 7871
rect 23768 7868 23796 8044
rect 23845 8041 23857 8075
rect 23891 8072 23903 8075
rect 24578 8072 24584 8084
rect 23891 8044 24584 8072
rect 23891 8041 23903 8044
rect 23845 8035 23903 8041
rect 24578 8032 24584 8044
rect 24636 8032 24642 8084
rect 32858 8032 32864 8084
rect 32916 8072 32922 8084
rect 33965 8075 34023 8081
rect 33965 8072 33977 8075
rect 32916 8044 33977 8072
rect 32916 8032 32922 8044
rect 33965 8041 33977 8044
rect 34011 8041 34023 8075
rect 33965 8035 34023 8041
rect 39117 8075 39175 8081
rect 39117 8041 39129 8075
rect 39163 8072 39175 8075
rect 40034 8072 40040 8084
rect 39163 8044 40040 8072
rect 39163 8041 39175 8044
rect 39117 8035 39175 8041
rect 40034 8032 40040 8044
rect 40092 8032 40098 8084
rect 41230 8072 41236 8084
rect 41191 8044 41236 8072
rect 41230 8032 41236 8044
rect 41288 8032 41294 8084
rect 42702 8032 42708 8084
rect 42760 8072 42766 8084
rect 43993 8075 44051 8081
rect 43993 8072 44005 8075
rect 42760 8044 44005 8072
rect 42760 8032 42766 8044
rect 43993 8041 44005 8044
rect 44039 8041 44051 8075
rect 43993 8035 44051 8041
rect 33226 7964 33232 8016
rect 33284 8004 33290 8016
rect 35345 8007 35403 8013
rect 35345 8004 35357 8007
rect 33284 7976 35357 8004
rect 33284 7964 33290 7976
rect 35345 7973 35357 7976
rect 35391 7973 35403 8007
rect 35345 7967 35403 7973
rect 26234 7896 26240 7948
rect 26292 7936 26298 7948
rect 26421 7939 26479 7945
rect 26421 7936 26433 7939
rect 26292 7908 26433 7936
rect 26292 7896 26298 7908
rect 26421 7905 26433 7908
rect 26467 7905 26479 7939
rect 26421 7899 26479 7905
rect 27706 7896 27712 7948
rect 27764 7936 27770 7948
rect 28810 7936 28816 7948
rect 27764 7908 28816 7936
rect 27764 7896 27770 7908
rect 28810 7896 28816 7908
rect 28868 7896 28874 7948
rect 33502 7896 33508 7948
rect 33560 7936 33566 7948
rect 33560 7908 34928 7936
rect 33560 7896 33566 7908
rect 24486 7868 24492 7880
rect 23768 7840 24492 7868
rect 22732 7831 22790 7837
rect 24486 7828 24492 7840
rect 24544 7868 24550 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24544 7840 24593 7868
rect 24544 7828 24550 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 24848 7871 24906 7877
rect 24848 7837 24860 7871
rect 24894 7868 24906 7871
rect 25222 7868 25228 7880
rect 24894 7840 25228 7868
rect 24894 7837 24906 7840
rect 24848 7831 24906 7837
rect 25222 7828 25228 7840
rect 25280 7828 25286 7880
rect 29730 7868 29736 7880
rect 29691 7840 29736 7868
rect 29730 7828 29736 7840
rect 29788 7828 29794 7880
rect 30000 7871 30058 7877
rect 30000 7837 30012 7871
rect 30046 7868 30058 7871
rect 30282 7868 30288 7880
rect 30046 7840 30288 7868
rect 30046 7837 30058 7840
rect 30000 7831 30058 7837
rect 30282 7828 30288 7840
rect 30340 7828 30346 7880
rect 32125 7871 32183 7877
rect 32125 7837 32137 7871
rect 32171 7868 32183 7871
rect 32214 7868 32220 7880
rect 32171 7840 32220 7868
rect 32171 7837 32183 7840
rect 32125 7831 32183 7837
rect 32214 7828 32220 7840
rect 32272 7828 32278 7880
rect 32392 7871 32450 7877
rect 32392 7837 32404 7871
rect 32438 7837 32450 7871
rect 32392 7831 32450 7837
rect 4240 7803 4298 7809
rect 4240 7769 4252 7803
rect 4286 7800 4298 7803
rect 5534 7800 5540 7812
rect 4286 7772 5540 7800
rect 4286 7769 4298 7772
rect 4240 7763 4298 7769
rect 5534 7760 5540 7772
rect 5592 7760 5598 7812
rect 6270 7760 6276 7812
rect 6328 7800 6334 7812
rect 6702 7803 6760 7809
rect 6702 7800 6714 7803
rect 6328 7772 6714 7800
rect 6328 7760 6334 7772
rect 6702 7769 6714 7772
rect 6748 7769 6760 7803
rect 6702 7763 6760 7769
rect 8570 7760 8576 7812
rect 8628 7800 8634 7812
rect 9186 7803 9244 7809
rect 9186 7800 9198 7803
rect 8628 7772 9198 7800
rect 8628 7760 8634 7772
rect 9186 7769 9198 7772
rect 9232 7769 9244 7803
rect 9186 7763 9244 7769
rect 11054 7760 11060 7812
rect 11112 7800 11118 7812
rect 12130 7803 12188 7809
rect 12130 7800 12142 7803
rect 11112 7772 12142 7800
rect 11112 7760 11118 7772
rect 12130 7769 12142 7772
rect 12176 7769 12188 7803
rect 12130 7763 12188 7769
rect 14452 7803 14510 7809
rect 14452 7769 14464 7803
rect 14498 7800 14510 7803
rect 19490 7803 19548 7809
rect 19490 7800 19502 7803
rect 14498 7772 17264 7800
rect 14498 7769 14510 7772
rect 14452 7763 14510 7769
rect 10321 7735 10379 7741
rect 10321 7701 10333 7735
rect 10367 7732 10379 7735
rect 11698 7732 11704 7744
rect 10367 7704 11704 7732
rect 10367 7701 10379 7704
rect 10321 7695 10379 7701
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 13262 7732 13268 7744
rect 13175 7704 13268 7732
rect 13262 7692 13268 7704
rect 13320 7732 13326 7744
rect 17236 7741 17264 7772
rect 18524 7772 19502 7800
rect 18524 7741 18552 7772
rect 19490 7769 19502 7772
rect 19536 7769 19548 7803
rect 19490 7763 19548 7769
rect 22646 7760 22652 7812
rect 22704 7760 22710 7812
rect 25884 7772 26280 7800
rect 16393 7735 16451 7741
rect 16393 7732 16405 7735
rect 13320 7704 16405 7732
rect 13320 7692 13326 7704
rect 16393 7701 16405 7704
rect 16439 7701 16451 7735
rect 16393 7695 16451 7701
rect 17221 7735 17279 7741
rect 17221 7701 17233 7735
rect 17267 7701 17279 7735
rect 17221 7695 17279 7701
rect 18509 7735 18567 7741
rect 18509 7701 18521 7735
rect 18555 7701 18567 7735
rect 18509 7695 18567 7701
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 20625 7735 20683 7741
rect 20625 7732 20637 7735
rect 19392 7704 20637 7732
rect 19392 7692 19398 7704
rect 20625 7701 20637 7704
rect 20671 7732 20683 7735
rect 21453 7735 21511 7741
rect 21453 7732 21465 7735
rect 20671 7704 21465 7732
rect 20671 7701 20683 7704
rect 20625 7695 20683 7701
rect 21453 7701 21465 7704
rect 21499 7701 21511 7735
rect 21453 7695 21511 7701
rect 21545 7735 21603 7741
rect 21545 7701 21557 7735
rect 21591 7732 21603 7735
rect 25884 7732 25912 7772
rect 21591 7704 25912 7732
rect 25961 7735 26019 7741
rect 21591 7701 21603 7704
rect 21545 7695 21603 7701
rect 25961 7701 25973 7735
rect 26007 7732 26019 7735
rect 26142 7732 26148 7744
rect 26007 7704 26148 7732
rect 26007 7701 26019 7704
rect 25961 7695 26019 7701
rect 26142 7692 26148 7704
rect 26200 7692 26206 7744
rect 26252 7732 26280 7772
rect 26326 7760 26332 7812
rect 26384 7800 26390 7812
rect 26666 7803 26724 7809
rect 26666 7800 26678 7803
rect 26384 7772 26678 7800
rect 26384 7760 26390 7772
rect 26666 7769 26678 7772
rect 26712 7769 26724 7803
rect 28629 7803 28687 7809
rect 28629 7800 28641 7803
rect 26666 7763 26724 7769
rect 27816 7772 28641 7800
rect 27816 7741 27844 7772
rect 28629 7769 28641 7772
rect 28675 7769 28687 7803
rect 28629 7763 28687 7769
rect 32306 7760 32312 7812
rect 32364 7800 32370 7812
rect 32416 7800 32444 7831
rect 33686 7828 33692 7880
rect 33744 7868 33750 7880
rect 33965 7871 34023 7877
rect 33965 7868 33977 7871
rect 33744 7840 33977 7868
rect 33744 7828 33750 7840
rect 33965 7837 33977 7840
rect 34011 7837 34023 7871
rect 33965 7831 34023 7837
rect 34149 7871 34207 7877
rect 34149 7837 34161 7871
rect 34195 7868 34207 7871
rect 34606 7868 34612 7880
rect 34195 7840 34612 7868
rect 34195 7837 34207 7840
rect 34149 7831 34207 7837
rect 34606 7828 34612 7840
rect 34664 7828 34670 7880
rect 34900 7877 34928 7908
rect 38930 7896 38936 7948
rect 38988 7936 38994 7948
rect 39850 7936 39856 7948
rect 38988 7908 39344 7936
rect 39811 7908 39856 7936
rect 38988 7896 38994 7908
rect 34885 7871 34943 7877
rect 34885 7837 34897 7871
rect 34931 7837 34943 7871
rect 34885 7831 34943 7837
rect 35529 7871 35587 7877
rect 35529 7837 35541 7871
rect 35575 7837 35587 7871
rect 39114 7868 39120 7880
rect 39075 7840 39120 7868
rect 35529 7831 35587 7837
rect 32364 7772 32444 7800
rect 32364 7760 32370 7772
rect 32490 7760 32496 7812
rect 32548 7800 32554 7812
rect 35544 7800 35572 7831
rect 39114 7828 39120 7840
rect 39172 7828 39178 7880
rect 39316 7877 39344 7908
rect 39850 7896 39856 7908
rect 39908 7896 39914 7948
rect 41138 7896 41144 7948
rect 41196 7936 41202 7948
rect 41693 7939 41751 7945
rect 41693 7936 41705 7939
rect 41196 7908 41705 7936
rect 41196 7896 41202 7908
rect 41693 7905 41705 7908
rect 41739 7905 41751 7939
rect 41693 7899 41751 7905
rect 39301 7871 39359 7877
rect 39301 7837 39313 7871
rect 39347 7868 39359 7871
rect 39390 7868 39396 7880
rect 39347 7840 39396 7868
rect 39347 7837 39359 7840
rect 39301 7831 39359 7837
rect 39390 7828 39396 7840
rect 39448 7828 39454 7880
rect 41874 7868 41880 7880
rect 41787 7840 41880 7868
rect 41874 7828 41880 7840
rect 41932 7868 41938 7880
rect 42610 7868 42616 7880
rect 41932 7840 42616 7868
rect 41932 7828 41938 7840
rect 42610 7828 42616 7840
rect 42668 7828 42674 7880
rect 44174 7868 44180 7880
rect 44135 7840 44180 7868
rect 44174 7828 44180 7840
rect 44232 7828 44238 7880
rect 32548 7772 35572 7800
rect 32548 7760 32554 7772
rect 39850 7760 39856 7812
rect 39908 7800 39914 7812
rect 40098 7803 40156 7809
rect 40098 7800 40110 7803
rect 39908 7772 40110 7800
rect 39908 7760 39914 7772
rect 40098 7769 40110 7772
rect 40144 7769 40156 7803
rect 40098 7763 40156 7769
rect 27801 7735 27859 7741
rect 27801 7732 27813 7735
rect 26252 7704 27813 7732
rect 27801 7701 27813 7704
rect 27847 7701 27859 7735
rect 28258 7732 28264 7744
rect 28219 7704 28264 7732
rect 27801 7695 27859 7701
rect 28258 7692 28264 7704
rect 28316 7692 28322 7744
rect 28721 7735 28779 7741
rect 28721 7701 28733 7735
rect 28767 7732 28779 7735
rect 28810 7732 28816 7744
rect 28767 7704 28816 7732
rect 28767 7701 28779 7704
rect 28721 7695 28779 7701
rect 28810 7692 28816 7704
rect 28868 7692 28874 7744
rect 30006 7692 30012 7744
rect 30064 7732 30070 7744
rect 31113 7735 31171 7741
rect 31113 7732 31125 7735
rect 30064 7704 31125 7732
rect 30064 7692 30070 7704
rect 31113 7701 31125 7704
rect 31159 7701 31171 7735
rect 31113 7695 31171 7701
rect 32122 7692 32128 7744
rect 32180 7732 32186 7744
rect 33505 7735 33563 7741
rect 33505 7732 33517 7735
rect 32180 7704 33517 7732
rect 32180 7692 32186 7704
rect 33505 7701 33517 7704
rect 33551 7701 33563 7735
rect 34698 7732 34704 7744
rect 34611 7704 34704 7732
rect 33505 7695 33563 7701
rect 34698 7692 34704 7704
rect 34756 7732 34762 7744
rect 40402 7732 40408 7744
rect 34756 7704 40408 7732
rect 34756 7692 34762 7704
rect 40402 7692 40408 7704
rect 40460 7692 40466 7744
rect 41138 7692 41144 7744
rect 41196 7732 41202 7744
rect 42061 7735 42119 7741
rect 42061 7732 42073 7735
rect 41196 7704 42073 7732
rect 41196 7692 41202 7704
rect 42061 7701 42073 7704
rect 42107 7701 42119 7735
rect 42061 7695 42119 7701
rect 1104 7642 45056 7664
rect 1104 7590 11898 7642
rect 11950 7590 11962 7642
rect 12014 7590 12026 7642
rect 12078 7590 12090 7642
rect 12142 7590 12154 7642
rect 12206 7590 22846 7642
rect 22898 7590 22910 7642
rect 22962 7590 22974 7642
rect 23026 7590 23038 7642
rect 23090 7590 23102 7642
rect 23154 7590 33794 7642
rect 33846 7590 33858 7642
rect 33910 7590 33922 7642
rect 33974 7590 33986 7642
rect 34038 7590 34050 7642
rect 34102 7590 44742 7642
rect 44794 7590 44806 7642
rect 44858 7590 44870 7642
rect 44922 7590 44934 7642
rect 44986 7590 44998 7642
rect 45050 7590 45056 7642
rect 1104 7568 45056 7590
rect 3510 7488 3516 7540
rect 3568 7528 3574 7540
rect 3881 7531 3939 7537
rect 3881 7528 3893 7531
rect 3568 7500 3893 7528
rect 3568 7488 3574 7500
rect 3881 7497 3893 7500
rect 3927 7497 3939 7531
rect 3881 7491 3939 7497
rect 5166 7488 5172 7540
rect 5224 7528 5230 7540
rect 10597 7531 10655 7537
rect 10597 7528 10609 7531
rect 5224 7500 10609 7528
rect 5224 7488 5230 7500
rect 10597 7497 10609 7500
rect 10643 7497 10655 7531
rect 10597 7491 10655 7497
rect 12069 7531 12127 7537
rect 12069 7497 12081 7531
rect 12115 7528 12127 7531
rect 12802 7528 12808 7540
rect 12115 7500 12808 7528
rect 12115 7497 12127 7500
rect 12069 7491 12127 7497
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 15378 7528 15384 7540
rect 14783 7500 15384 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 15565 7531 15623 7537
rect 15565 7528 15577 7531
rect 15528 7500 15577 7528
rect 15528 7488 15534 7500
rect 15565 7497 15577 7500
rect 15611 7497 15623 7531
rect 15565 7491 15623 7497
rect 17313 7531 17371 7537
rect 17313 7497 17325 7531
rect 17359 7528 17371 7531
rect 19334 7528 19340 7540
rect 17359 7500 19340 7528
rect 17359 7497 17371 7500
rect 17313 7491 17371 7497
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 19429 7531 19487 7537
rect 19429 7497 19441 7531
rect 19475 7528 19487 7531
rect 20346 7528 20352 7540
rect 19475 7500 20352 7528
rect 19475 7497 19487 7500
rect 19429 7491 19487 7497
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 22189 7531 22247 7537
rect 22189 7497 22201 7531
rect 22235 7497 22247 7531
rect 22646 7528 22652 7540
rect 22607 7500 22652 7528
rect 22189 7491 22247 7497
rect 2593 7463 2651 7469
rect 2593 7429 2605 7463
rect 2639 7460 2651 7463
rect 7374 7460 7380 7472
rect 2639 7432 7380 7460
rect 2639 7429 2651 7432
rect 2593 7423 2651 7429
rect 7374 7420 7380 7432
rect 7432 7460 7438 7472
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 7432 7432 7849 7460
rect 7432 7420 7438 7432
rect 7837 7429 7849 7432
rect 7883 7429 7895 7463
rect 9490 7460 9496 7472
rect 9451 7432 9496 7460
rect 7837 7423 7895 7429
rect 9490 7420 9496 7432
rect 9548 7460 9554 7472
rect 10413 7463 10471 7469
rect 10413 7460 10425 7463
rect 9548 7432 10425 7460
rect 9548 7420 9554 7432
rect 10413 7429 10425 7432
rect 10459 7429 10471 7463
rect 10413 7423 10471 7429
rect 10689 7463 10747 7469
rect 10689 7429 10701 7463
rect 10735 7460 10747 7463
rect 10778 7460 10784 7472
rect 10735 7432 10784 7460
rect 10735 7429 10747 7432
rect 10689 7423 10747 7429
rect 10778 7420 10784 7432
rect 10836 7420 10842 7472
rect 11698 7420 11704 7472
rect 11756 7460 11762 7472
rect 12161 7463 12219 7469
rect 12161 7460 12173 7463
rect 11756 7432 12173 7460
rect 11756 7420 11762 7432
rect 12161 7429 12173 7432
rect 12207 7429 12219 7463
rect 15396 7460 15424 7488
rect 17221 7463 17279 7469
rect 17221 7460 17233 7463
rect 15396 7432 17233 7460
rect 12161 7423 12219 7429
rect 17221 7429 17233 7432
rect 17267 7429 17279 7463
rect 17221 7423 17279 7429
rect 19242 7420 19248 7472
rect 19300 7460 19306 7472
rect 21818 7460 21824 7472
rect 19300 7432 21824 7460
rect 19300 7420 19306 7432
rect 13354 7392 13360 7404
rect 13315 7364 13360 7392
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 13624 7395 13682 7401
rect 13624 7361 13636 7395
rect 13670 7392 13682 7395
rect 14090 7392 14096 7404
rect 13670 7364 14096 7392
rect 13670 7361 13682 7364
rect 13624 7355 13682 7361
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 18322 7401 18328 7404
rect 18316 7355 18328 7401
rect 18380 7392 18386 7404
rect 19904 7401 19932 7432
rect 21818 7420 21824 7432
rect 21876 7420 21882 7472
rect 22204 7460 22232 7491
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 22738 7488 22744 7540
rect 22796 7528 22802 7540
rect 24121 7531 24179 7537
rect 24121 7528 24133 7531
rect 22796 7500 24133 7528
rect 22796 7488 22802 7500
rect 24121 7497 24133 7500
rect 24167 7497 24179 7531
rect 26142 7528 26148 7540
rect 26103 7500 26148 7528
rect 24121 7491 24179 7497
rect 26142 7488 26148 7500
rect 26200 7488 26206 7540
rect 27157 7531 27215 7537
rect 27157 7497 27169 7531
rect 27203 7528 27215 7531
rect 27338 7528 27344 7540
rect 27203 7500 27344 7528
rect 27203 7497 27215 7500
rect 27157 7491 27215 7497
rect 27338 7488 27344 7500
rect 27396 7488 27402 7540
rect 27525 7531 27583 7537
rect 27525 7497 27537 7531
rect 27571 7528 27583 7531
rect 28810 7528 28816 7540
rect 27571 7500 28816 7528
rect 27571 7497 27583 7500
rect 27525 7491 27583 7497
rect 28810 7488 28816 7500
rect 28868 7488 28874 7540
rect 29638 7488 29644 7540
rect 29696 7528 29702 7540
rect 29917 7531 29975 7537
rect 29917 7528 29929 7531
rect 29696 7500 29929 7528
rect 29696 7488 29702 7500
rect 29917 7497 29929 7500
rect 29963 7497 29975 7531
rect 29917 7491 29975 7497
rect 32582 7488 32588 7540
rect 32640 7528 32646 7540
rect 34698 7528 34704 7540
rect 32640 7500 34704 7528
rect 32640 7488 32646 7500
rect 34698 7488 34704 7500
rect 34756 7488 34762 7540
rect 39850 7528 39856 7540
rect 39811 7500 39856 7528
rect 39850 7488 39856 7500
rect 39908 7488 39914 7540
rect 40770 7528 40776 7540
rect 40731 7500 40776 7528
rect 40770 7488 40776 7500
rect 40828 7488 40834 7540
rect 26053 7463 26111 7469
rect 22204 7432 23612 7460
rect 20162 7401 20168 7404
rect 19889 7395 19947 7401
rect 18380 7364 18416 7392
rect 18322 7352 18328 7355
rect 18380 7352 18386 7364
rect 19889 7361 19901 7395
rect 19935 7361 19947 7395
rect 20156 7392 20168 7401
rect 20123 7364 20168 7392
rect 19889 7355 19947 7361
rect 20156 7355 20168 7364
rect 20162 7352 20168 7355
rect 20220 7352 20226 7404
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7392 22615 7395
rect 23290 7392 23296 7404
rect 22603 7364 23296 7392
rect 22603 7361 22615 7364
rect 22557 7355 22615 7361
rect 23290 7352 23296 7364
rect 23348 7352 23354 7404
rect 23584 7401 23612 7432
rect 26053 7429 26065 7463
rect 26099 7460 26111 7463
rect 28258 7460 28264 7472
rect 26099 7432 28264 7460
rect 26099 7429 26111 7432
rect 26053 7423 26111 7429
rect 28258 7420 28264 7432
rect 28316 7420 28322 7472
rect 30006 7460 30012 7472
rect 28552 7432 30012 7460
rect 23569 7395 23627 7401
rect 23569 7361 23581 7395
rect 23615 7361 23627 7395
rect 24026 7392 24032 7404
rect 23987 7364 24032 7392
rect 23569 7355 23627 7361
rect 24026 7352 24032 7364
rect 24084 7352 24090 7404
rect 25225 7395 25283 7401
rect 25225 7361 25237 7395
rect 25271 7392 25283 7395
rect 26970 7392 26976 7404
rect 25271 7364 26976 7392
rect 25271 7361 25283 7364
rect 25225 7355 25283 7361
rect 26970 7352 26976 7364
rect 27028 7352 27034 7404
rect 27617 7395 27675 7401
rect 27617 7361 27629 7395
rect 27663 7392 27675 7395
rect 28552 7392 28580 7432
rect 30006 7420 30012 7432
rect 30064 7420 30070 7472
rect 32306 7420 32312 7472
rect 32364 7460 32370 7472
rect 33410 7460 33416 7472
rect 32364 7432 33416 7460
rect 32364 7420 32370 7432
rect 33410 7420 33416 7432
rect 33468 7420 33474 7472
rect 35802 7460 35808 7472
rect 34546 7432 35808 7460
rect 35802 7420 35808 7432
rect 35860 7420 35866 7472
rect 39224 7432 41092 7460
rect 27663 7364 28580 7392
rect 28629 7395 28687 7401
rect 27663 7361 27675 7364
rect 27617 7355 27675 7361
rect 28629 7361 28641 7395
rect 28675 7392 28687 7395
rect 28718 7392 28724 7404
rect 28675 7364 28724 7392
rect 28675 7361 28687 7364
rect 28629 7355 28687 7361
rect 28718 7352 28724 7364
rect 28776 7392 28782 7404
rect 30374 7392 30380 7404
rect 28776 7364 30380 7392
rect 28776 7352 28782 7364
rect 30374 7352 30380 7364
rect 30432 7352 30438 7404
rect 30929 7395 30987 7401
rect 30929 7361 30941 7395
rect 30975 7361 30987 7395
rect 32122 7392 32128 7404
rect 32083 7364 32128 7392
rect 30929 7355 30987 7361
rect 12342 7324 12348 7336
rect 12303 7296 12348 7324
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 15654 7324 15660 7336
rect 15615 7296 15660 7324
rect 15654 7284 15660 7296
rect 15712 7284 15718 7336
rect 15841 7327 15899 7333
rect 15841 7293 15853 7327
rect 15887 7324 15899 7327
rect 17494 7324 17500 7336
rect 15887 7296 17356 7324
rect 17455 7296 17500 7324
rect 15887 7293 15899 7296
rect 15841 7287 15899 7293
rect 15197 7259 15255 7265
rect 15197 7225 15209 7259
rect 15243 7256 15255 7259
rect 16666 7256 16672 7268
rect 15243 7228 16672 7256
rect 15243 7225 15255 7228
rect 15197 7219 15255 7225
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 10137 7191 10195 7197
rect 10137 7157 10149 7191
rect 10183 7188 10195 7191
rect 11238 7188 11244 7200
rect 10183 7160 11244 7188
rect 10183 7157 10195 7160
rect 10137 7151 10195 7157
rect 11238 7148 11244 7160
rect 11296 7148 11302 7200
rect 11698 7188 11704 7200
rect 11659 7160 11704 7188
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 16850 7188 16856 7200
rect 16811 7160 16856 7188
rect 16850 7148 16856 7160
rect 16908 7148 16914 7200
rect 17328 7188 17356 7296
rect 17494 7284 17500 7296
rect 17552 7284 17558 7336
rect 18046 7324 18052 7336
rect 18007 7296 18052 7324
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 22833 7327 22891 7333
rect 22833 7293 22845 7327
rect 22879 7293 22891 7327
rect 22833 7287 22891 7293
rect 21358 7216 21364 7268
rect 21416 7256 21422 7268
rect 22848 7256 22876 7287
rect 26050 7284 26056 7336
rect 26108 7324 26114 7336
rect 26237 7327 26295 7333
rect 26237 7324 26249 7327
rect 26108 7296 26249 7324
rect 26108 7284 26114 7296
rect 26237 7293 26249 7296
rect 26283 7293 26295 7327
rect 27706 7324 27712 7336
rect 27667 7296 27712 7324
rect 26237 7287 26295 7293
rect 27706 7284 27712 7296
rect 27764 7284 27770 7336
rect 29914 7284 29920 7336
rect 29972 7324 29978 7336
rect 30944 7324 30972 7355
rect 32122 7352 32128 7364
rect 32180 7352 32186 7404
rect 32214 7352 32220 7404
rect 32272 7392 32278 7404
rect 32674 7392 32680 7404
rect 32272 7364 32680 7392
rect 32272 7352 32278 7364
rect 32674 7352 32680 7364
rect 32732 7392 32738 7404
rect 33042 7392 33048 7404
rect 32732 7364 33048 7392
rect 32732 7352 32738 7364
rect 33042 7352 33048 7364
rect 33100 7352 33106 7404
rect 39224 7401 39252 7432
rect 39209 7395 39267 7401
rect 39209 7361 39221 7395
rect 39255 7361 39267 7395
rect 39390 7392 39396 7404
rect 39351 7364 39396 7392
rect 39209 7355 39267 7361
rect 39390 7352 39396 7364
rect 39448 7392 39454 7404
rect 39942 7392 39948 7404
rect 39448 7364 39948 7392
rect 39448 7352 39454 7364
rect 39942 7352 39948 7364
rect 40000 7352 40006 7404
rect 40037 7395 40095 7401
rect 40037 7361 40049 7395
rect 40083 7361 40095 7395
rect 40310 7392 40316 7404
rect 40271 7364 40316 7392
rect 40037 7355 40095 7361
rect 29972 7296 30972 7324
rect 29972 7284 29978 7296
rect 31294 7284 31300 7336
rect 31352 7324 31358 7336
rect 32232 7324 32260 7352
rect 31352 7296 32260 7324
rect 33321 7327 33379 7333
rect 31352 7284 31358 7296
rect 33321 7293 33333 7327
rect 33367 7324 33379 7327
rect 35342 7324 35348 7336
rect 33367 7296 35348 7324
rect 33367 7293 33379 7296
rect 33321 7287 33379 7293
rect 35342 7284 35348 7296
rect 35400 7284 35406 7336
rect 39301 7327 39359 7333
rect 39301 7293 39313 7327
rect 39347 7324 39359 7327
rect 40052 7324 40080 7355
rect 40310 7352 40316 7364
rect 40368 7352 40374 7404
rect 40954 7392 40960 7404
rect 40915 7364 40960 7392
rect 40954 7352 40960 7364
rect 41012 7352 41018 7404
rect 41064 7392 41092 7432
rect 41138 7392 41144 7404
rect 41064 7364 41144 7392
rect 41138 7352 41144 7364
rect 41196 7352 41202 7404
rect 41233 7395 41291 7401
rect 41233 7361 41245 7395
rect 41279 7392 41291 7395
rect 41506 7392 41512 7404
rect 41279 7364 41512 7392
rect 41279 7361 41291 7364
rect 41233 7355 41291 7361
rect 41506 7352 41512 7364
rect 41564 7352 41570 7404
rect 39347 7296 40080 7324
rect 39347 7293 39359 7296
rect 39301 7287 39359 7293
rect 40402 7284 40408 7336
rect 40460 7324 40466 7336
rect 43898 7324 43904 7336
rect 40460 7296 43904 7324
rect 40460 7284 40466 7296
rect 43898 7284 43904 7296
rect 43956 7284 43962 7336
rect 21416 7228 22876 7256
rect 25041 7259 25099 7265
rect 21416 7216 21422 7228
rect 25041 7225 25053 7259
rect 25087 7256 25099 7259
rect 26142 7256 26148 7268
rect 25087 7228 26148 7256
rect 25087 7225 25099 7228
rect 25041 7219 25099 7225
rect 26142 7216 26148 7228
rect 26200 7216 26206 7268
rect 40221 7259 40279 7265
rect 40221 7225 40233 7259
rect 40267 7256 40279 7259
rect 40267 7228 41276 7256
rect 40267 7225 40279 7228
rect 40221 7219 40279 7225
rect 18690 7188 18696 7200
rect 17328 7160 18696 7188
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 20806 7148 20812 7200
rect 20864 7188 20870 7200
rect 21269 7191 21327 7197
rect 21269 7188 21281 7191
rect 20864 7160 21281 7188
rect 20864 7148 20870 7160
rect 21269 7157 21281 7160
rect 21315 7157 21327 7191
rect 21269 7151 21327 7157
rect 22370 7148 22376 7200
rect 22428 7188 22434 7200
rect 23385 7191 23443 7197
rect 23385 7188 23397 7191
rect 22428 7160 23397 7188
rect 22428 7148 22434 7160
rect 23385 7157 23397 7160
rect 23431 7157 23443 7191
rect 23385 7151 23443 7157
rect 25685 7191 25743 7197
rect 25685 7157 25697 7191
rect 25731 7188 25743 7191
rect 25774 7188 25780 7200
rect 25731 7160 25780 7188
rect 25731 7157 25743 7160
rect 25685 7151 25743 7157
rect 25774 7148 25780 7160
rect 25832 7148 25838 7200
rect 31018 7188 31024 7200
rect 30979 7160 31024 7188
rect 31018 7148 31024 7160
rect 31076 7148 31082 7200
rect 32309 7191 32367 7197
rect 32309 7157 32321 7191
rect 32355 7188 32367 7191
rect 32766 7188 32772 7200
rect 32355 7160 32772 7188
rect 32355 7157 32367 7160
rect 32309 7151 32367 7157
rect 32766 7148 32772 7160
rect 32824 7148 32830 7200
rect 34790 7188 34796 7200
rect 34751 7160 34796 7188
rect 34790 7148 34796 7160
rect 34848 7148 34854 7200
rect 41248 7188 41276 7228
rect 41874 7188 41880 7200
rect 41248 7160 41880 7188
rect 41874 7148 41880 7160
rect 41932 7148 41938 7200
rect 1104 7098 44896 7120
rect 1104 7046 6424 7098
rect 6476 7046 6488 7098
rect 6540 7046 6552 7098
rect 6604 7046 6616 7098
rect 6668 7046 6680 7098
rect 6732 7046 17372 7098
rect 17424 7046 17436 7098
rect 17488 7046 17500 7098
rect 17552 7046 17564 7098
rect 17616 7046 17628 7098
rect 17680 7046 28320 7098
rect 28372 7046 28384 7098
rect 28436 7046 28448 7098
rect 28500 7046 28512 7098
rect 28564 7046 28576 7098
rect 28628 7046 39268 7098
rect 39320 7046 39332 7098
rect 39384 7046 39396 7098
rect 39448 7046 39460 7098
rect 39512 7046 39524 7098
rect 39576 7046 44896 7098
rect 1104 7024 44896 7046
rect 8404 6956 9352 6984
rect 8404 6925 8432 6956
rect 8389 6919 8447 6925
rect 8389 6885 8401 6919
rect 8435 6885 8447 6919
rect 9217 6919 9275 6925
rect 8389 6879 8447 6885
rect 8496 6888 8800 6916
rect 7006 6848 7012 6860
rect 6967 6820 7012 6848
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 5810 6740 5816 6792
rect 5868 6780 5874 6792
rect 6549 6783 6607 6789
rect 6549 6780 6561 6783
rect 5868 6752 6561 6780
rect 5868 6740 5874 6752
rect 6549 6749 6561 6752
rect 6595 6749 6607 6783
rect 8496 6780 8524 6888
rect 8772 6848 8800 6888
rect 9217 6885 9229 6919
rect 9263 6885 9275 6919
rect 9217 6879 9275 6885
rect 9232 6848 9260 6879
rect 8772 6820 9260 6848
rect 9324 6848 9352 6956
rect 15654 6944 15660 6996
rect 15712 6984 15718 6996
rect 16025 6987 16083 6993
rect 16025 6984 16037 6987
rect 15712 6956 16037 6984
rect 15712 6944 15718 6956
rect 16025 6953 16037 6956
rect 16071 6953 16083 6987
rect 16025 6947 16083 6953
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 18509 6987 18567 6993
rect 18509 6984 18521 6987
rect 18380 6956 18521 6984
rect 18380 6944 18386 6956
rect 18509 6953 18521 6956
rect 18555 6953 18567 6987
rect 18509 6947 18567 6953
rect 18690 6944 18696 6996
rect 18748 6984 18754 6996
rect 23290 6984 23296 6996
rect 18748 6956 23152 6984
rect 23251 6956 23296 6984
rect 18748 6944 18754 6956
rect 12342 6876 12348 6928
rect 12400 6916 12406 6928
rect 12400 6888 13492 6916
rect 12400 6876 12406 6888
rect 13464 6860 13492 6888
rect 20254 6876 20260 6928
rect 20312 6916 20318 6928
rect 23124 6916 23152 6956
rect 23290 6944 23296 6956
rect 23348 6944 23354 6996
rect 26050 6944 26056 6996
rect 26108 6984 26114 6996
rect 26421 6987 26479 6993
rect 26421 6984 26433 6987
rect 26108 6956 26433 6984
rect 26108 6944 26114 6956
rect 26421 6953 26433 6956
rect 26467 6953 26479 6987
rect 27706 6984 27712 6996
rect 26421 6947 26479 6953
rect 26988 6956 27712 6984
rect 26988 6916 27016 6956
rect 27706 6944 27712 6956
rect 27764 6944 27770 6996
rect 28353 6987 28411 6993
rect 28353 6953 28365 6987
rect 28399 6984 28411 6987
rect 28810 6984 28816 6996
rect 28399 6956 28816 6984
rect 28399 6953 28411 6956
rect 28353 6947 28411 6953
rect 28810 6944 28816 6956
rect 28868 6944 28874 6996
rect 30088 6987 30146 6993
rect 30088 6953 30100 6987
rect 30134 6984 30146 6987
rect 32582 6984 32588 6996
rect 30134 6956 32588 6984
rect 30134 6953 30146 6956
rect 30088 6947 30146 6953
rect 32582 6944 32588 6956
rect 32640 6944 32646 6996
rect 40037 6987 40095 6993
rect 40037 6953 40049 6987
rect 40083 6984 40095 6987
rect 40954 6984 40960 6996
rect 40083 6956 40960 6984
rect 40083 6953 40095 6956
rect 40037 6947 40095 6953
rect 40954 6944 40960 6956
rect 41012 6944 41018 6996
rect 20312 6888 21220 6916
rect 23124 6888 27016 6916
rect 20312 6876 20318 6888
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 9324 6820 10916 6848
rect 9674 6780 9680 6792
rect 6549 6743 6607 6749
rect 7208 6752 8524 6780
rect 8772 6752 9680 6780
rect 5994 6672 6000 6724
rect 6052 6712 6058 6724
rect 7208 6712 7236 6752
rect 6052 6684 7236 6712
rect 7276 6715 7334 6721
rect 6052 6672 6058 6684
rect 7276 6681 7288 6715
rect 7322 6712 7334 6715
rect 8202 6712 8208 6724
rect 7322 6684 8208 6712
rect 7322 6681 7334 6684
rect 7276 6675 7334 6681
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 6365 6647 6423 6653
rect 6365 6613 6377 6647
rect 6411 6644 6423 6647
rect 8772 6644 8800 6752
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 9858 6780 9864 6792
rect 9819 6752 9864 6780
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10042 6780 10048 6792
rect 10003 6752 10048 6780
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 10778 6780 10784 6792
rect 10739 6752 10784 6780
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 10888 6780 10916 6820
rect 12406 6820 13277 6848
rect 12406 6780 12434 6820
rect 13265 6817 13277 6820
rect 13311 6817 13323 6851
rect 13446 6848 13452 6860
rect 13407 6820 13452 6848
rect 13265 6811 13323 6817
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 16850 6848 16856 6860
rect 15672 6820 16856 6848
rect 10888 6752 12434 6780
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6780 14703 6783
rect 14734 6780 14740 6792
rect 14691 6752 14740 6780
rect 14691 6749 14703 6752
rect 14645 6743 14703 6749
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 15672 6780 15700 6820
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 16942 6808 16948 6860
rect 17000 6848 17006 6860
rect 21192 6857 21220 6888
rect 31110 6876 31116 6928
rect 31168 6916 31174 6928
rect 31168 6888 31984 6916
rect 31168 6876 31174 6888
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 17000 6820 19257 6848
rect 17000 6808 17006 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 21177 6851 21235 6857
rect 21177 6817 21189 6851
rect 21223 6817 21235 6851
rect 21358 6848 21364 6860
rect 21319 6820 21364 6848
rect 21177 6811 21235 6817
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 26234 6808 26240 6860
rect 26292 6848 26298 6860
rect 26970 6848 26976 6860
rect 26292 6820 26976 6848
rect 26292 6808 26298 6820
rect 26970 6808 26976 6820
rect 27028 6808 27034 6860
rect 29730 6808 29736 6860
rect 29788 6848 29794 6860
rect 29825 6851 29883 6857
rect 29825 6848 29837 6851
rect 29788 6820 29837 6848
rect 29788 6808 29794 6820
rect 29825 6817 29837 6820
rect 29871 6848 29883 6851
rect 31294 6848 31300 6860
rect 29871 6820 31300 6848
rect 29871 6817 29883 6820
rect 29825 6811 29883 6817
rect 31294 6808 31300 6820
rect 31352 6808 31358 6860
rect 14844 6752 15700 6780
rect 8938 6712 8944 6724
rect 8899 6684 8944 6712
rect 8938 6672 8944 6684
rect 8996 6672 9002 6724
rect 9030 6672 9036 6724
rect 9088 6712 9094 6724
rect 10229 6715 10287 6721
rect 10229 6712 10241 6715
rect 9088 6684 10241 6712
rect 9088 6672 9094 6684
rect 10229 6681 10241 6684
rect 10275 6681 10287 6715
rect 10229 6675 10287 6681
rect 10318 6672 10324 6724
rect 10376 6712 10382 6724
rect 11026 6715 11084 6721
rect 11026 6712 11038 6715
rect 10376 6684 11038 6712
rect 10376 6672 10382 6684
rect 11026 6681 11038 6684
rect 11072 6681 11084 6715
rect 11026 6675 11084 6681
rect 13173 6715 13231 6721
rect 13173 6681 13185 6715
rect 13219 6712 13231 6715
rect 14844 6712 14872 6752
rect 15746 6740 15752 6792
rect 15804 6780 15810 6792
rect 16669 6783 16727 6789
rect 16669 6780 16681 6783
rect 15804 6752 16681 6780
rect 15804 6740 15810 6752
rect 16669 6749 16681 6752
rect 16715 6749 16727 6783
rect 16669 6743 16727 6749
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6749 18751 6783
rect 18693 6743 18751 6749
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 20806 6780 20812 6792
rect 19475 6752 20812 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 13219 6684 14872 6712
rect 14912 6715 14970 6721
rect 13219 6681 13231 6684
rect 13173 6675 13231 6681
rect 14912 6681 14924 6715
rect 14958 6712 14970 6715
rect 18708 6712 18736 6743
rect 20806 6740 20812 6752
rect 20864 6740 20870 6792
rect 21913 6783 21971 6789
rect 21913 6749 21925 6783
rect 21959 6780 21971 6783
rect 25774 6780 25780 6792
rect 21959 6752 22324 6780
rect 25735 6752 25780 6780
rect 21959 6749 21971 6752
rect 21913 6743 21971 6749
rect 22296 6724 22324 6752
rect 25774 6740 25780 6752
rect 25832 6740 25838 6792
rect 26142 6740 26148 6792
rect 26200 6780 26206 6792
rect 31956 6790 31984 6888
rect 32674 6848 32680 6860
rect 32635 6820 32680 6848
rect 32674 6808 32680 6820
rect 32732 6808 32738 6860
rect 39942 6808 39948 6860
rect 40000 6848 40006 6860
rect 40000 6820 40264 6848
rect 40000 6808 40006 6820
rect 32025 6793 32083 6799
rect 32025 6790 32037 6793
rect 27229 6783 27287 6789
rect 27229 6780 27241 6783
rect 26200 6752 27241 6780
rect 26200 6740 26206 6752
rect 27229 6749 27241 6752
rect 27275 6749 27287 6783
rect 31956 6762 32037 6790
rect 32025 6759 32037 6762
rect 32071 6759 32083 6793
rect 32025 6753 32083 6759
rect 32944 6783 33002 6789
rect 27229 6743 27287 6749
rect 32944 6749 32956 6783
rect 32990 6780 33002 6783
rect 33226 6780 33232 6792
rect 32990 6752 33232 6780
rect 32990 6749 33002 6752
rect 32944 6743 33002 6749
rect 33226 6740 33232 6752
rect 33284 6740 33290 6792
rect 40037 6783 40095 6789
rect 40037 6749 40049 6783
rect 40083 6780 40095 6783
rect 40126 6780 40132 6792
rect 40083 6752 40132 6780
rect 40083 6749 40095 6752
rect 40037 6743 40095 6749
rect 40126 6740 40132 6752
rect 40184 6740 40190 6792
rect 40236 6789 40264 6820
rect 40221 6783 40279 6789
rect 40221 6749 40233 6783
rect 40267 6749 40279 6783
rect 40221 6743 40279 6749
rect 19613 6715 19671 6721
rect 19613 6712 19625 6715
rect 14958 6684 16528 6712
rect 18708 6684 19625 6712
rect 14958 6681 14970 6684
rect 14912 6675 14970 6681
rect 6411 6616 8800 6644
rect 6411 6613 6423 6616
rect 6365 6607 6423 6613
rect 9122 6604 9128 6656
rect 9180 6644 9186 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 9180 6616 9413 6644
rect 9180 6604 9186 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9401 6607 9459 6613
rect 12161 6647 12219 6653
rect 12161 6613 12173 6647
rect 12207 6644 12219 6647
rect 12250 6644 12256 6656
rect 12207 6616 12256 6644
rect 12207 6613 12219 6616
rect 12161 6607 12219 6613
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12805 6647 12863 6653
rect 12805 6613 12817 6647
rect 12851 6644 12863 6647
rect 14274 6644 14280 6656
rect 12851 6616 14280 6644
rect 12851 6613 12863 6616
rect 12805 6607 12863 6613
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 16500 6653 16528 6684
rect 19613 6681 19625 6684
rect 19659 6681 19671 6715
rect 19613 6675 19671 6681
rect 22180 6715 22238 6721
rect 22180 6681 22192 6715
rect 22226 6681 22238 6715
rect 22180 6675 22238 6681
rect 16485 6647 16543 6653
rect 16485 6613 16497 6647
rect 16531 6613 16543 6647
rect 20714 6644 20720 6656
rect 20675 6616 20720 6644
rect 16485 6607 16543 6613
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 21082 6644 21088 6656
rect 21043 6616 21088 6644
rect 21082 6604 21088 6616
rect 21140 6604 21146 6656
rect 22204 6644 22232 6675
rect 22278 6672 22284 6724
rect 22336 6672 22342 6724
rect 26329 6715 26387 6721
rect 26329 6681 26341 6715
rect 26375 6712 26387 6715
rect 27338 6712 27344 6724
rect 26375 6684 27344 6712
rect 26375 6681 26387 6684
rect 26329 6675 26387 6681
rect 27338 6672 27344 6684
rect 27396 6672 27402 6724
rect 31326 6684 31984 6712
rect 22370 6644 22376 6656
rect 22204 6616 22376 6644
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 25593 6647 25651 6653
rect 25593 6613 25605 6647
rect 25639 6644 25651 6647
rect 26234 6644 26240 6656
rect 25639 6616 26240 6644
rect 25639 6613 25651 6616
rect 25593 6607 25651 6613
rect 26234 6604 26240 6616
rect 26292 6604 26298 6656
rect 26418 6604 26424 6656
rect 26476 6644 26482 6656
rect 29086 6644 29092 6656
rect 26476 6616 29092 6644
rect 26476 6604 26482 6616
rect 29086 6604 29092 6616
rect 29144 6604 29150 6656
rect 30466 6604 30472 6656
rect 30524 6644 30530 6656
rect 31573 6647 31631 6653
rect 31573 6644 31585 6647
rect 30524 6616 31585 6644
rect 30524 6604 30530 6616
rect 31573 6613 31585 6616
rect 31619 6613 31631 6647
rect 31956 6644 31984 6684
rect 32030 6672 32036 6724
rect 32088 6712 32094 6724
rect 32088 6684 34100 6712
rect 32088 6672 32094 6684
rect 34072 6653 34100 6684
rect 32125 6647 32183 6653
rect 32125 6644 32137 6647
rect 31956 6616 32137 6644
rect 31573 6607 31631 6613
rect 32125 6613 32137 6616
rect 32171 6613 32183 6647
rect 32125 6607 32183 6613
rect 34057 6647 34115 6653
rect 34057 6613 34069 6647
rect 34103 6613 34115 6647
rect 34057 6607 34115 6613
rect 1104 6554 45056 6576
rect 1104 6502 11898 6554
rect 11950 6502 11962 6554
rect 12014 6502 12026 6554
rect 12078 6502 12090 6554
rect 12142 6502 12154 6554
rect 12206 6502 22846 6554
rect 22898 6502 22910 6554
rect 22962 6502 22974 6554
rect 23026 6502 23038 6554
rect 23090 6502 23102 6554
rect 23154 6502 33794 6554
rect 33846 6502 33858 6554
rect 33910 6502 33922 6554
rect 33974 6502 33986 6554
rect 34038 6502 34050 6554
rect 34102 6502 44742 6554
rect 44794 6502 44806 6554
rect 44858 6502 44870 6554
rect 44922 6502 44934 6554
rect 44986 6502 44998 6554
rect 45050 6502 45056 6554
rect 1104 6480 45056 6502
rect 8202 6440 8208 6452
rect 8163 6412 8208 6440
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 8941 6443 8999 6449
rect 8941 6409 8953 6443
rect 8987 6440 8999 6443
rect 10318 6440 10324 6452
rect 8987 6412 10324 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 11517 6443 11575 6449
rect 11517 6409 11529 6443
rect 11563 6440 11575 6443
rect 11790 6440 11796 6452
rect 11563 6412 11796 6440
rect 11563 6409 11575 6412
rect 11517 6403 11575 6409
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 17497 6443 17555 6449
rect 17497 6409 17509 6443
rect 17543 6409 17555 6443
rect 17954 6440 17960 6452
rect 17915 6412 17960 6440
rect 17497 6403 17555 6409
rect 7006 6372 7012 6384
rect 6380 6344 7012 6372
rect 6380 6313 6408 6344
rect 7006 6332 7012 6344
rect 7064 6372 7070 6384
rect 10778 6372 10784 6384
rect 7064 6344 10784 6372
rect 7064 6332 7070 6344
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6621 6307 6679 6313
rect 6621 6304 6633 6307
rect 6365 6267 6423 6273
rect 6472 6276 6633 6304
rect 5994 6196 6000 6248
rect 6052 6236 6058 6248
rect 6472 6236 6500 6276
rect 6621 6273 6633 6276
rect 6667 6273 6679 6307
rect 6621 6267 6679 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6304 8447 6307
rect 9030 6304 9036 6316
rect 8435 6276 9036 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9600 6313 9628 6344
rect 10778 6332 10784 6344
rect 10836 6372 10842 6384
rect 11606 6372 11612 6384
rect 10836 6344 11612 6372
rect 10836 6332 10842 6344
rect 11606 6332 11612 6344
rect 11664 6372 11670 6384
rect 12498 6375 12556 6381
rect 12498 6372 12510 6375
rect 11664 6344 12296 6372
rect 11664 6332 11670 6344
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 9852 6307 9910 6313
rect 9852 6273 9864 6307
rect 9898 6304 9910 6307
rect 11330 6304 11336 6316
rect 9898 6276 11336 6304
rect 9898 6273 9910 6276
rect 9852 6267 9910 6273
rect 6052 6208 6500 6236
rect 6052 6196 6058 6208
rect 7745 6171 7803 6177
rect 7745 6137 7757 6171
rect 7791 6168 7803 6171
rect 8938 6168 8944 6180
rect 7791 6140 8944 6168
rect 7791 6137 7803 6140
rect 7745 6131 7803 6137
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 9140 6100 9168 6267
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 11698 6304 11704 6316
rect 11659 6276 11704 6304
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 12268 6313 12296 6344
rect 12360 6344 12510 6372
rect 12253 6307 12311 6313
rect 12253 6273 12265 6307
rect 12299 6273 12311 6307
rect 12253 6267 12311 6273
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 12360 6236 12388 6344
rect 12498 6341 12510 6344
rect 12544 6341 12556 6375
rect 12498 6335 12556 6341
rect 14820 6375 14878 6381
rect 14820 6341 14832 6375
rect 14866 6372 14878 6375
rect 15194 6372 15200 6384
rect 14866 6344 15200 6372
rect 14866 6341 14878 6344
rect 14820 6335 14878 6341
rect 15194 6332 15200 6344
rect 15252 6332 15258 6384
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6304 14611 6307
rect 14642 6304 14648 6316
rect 14599 6276 14648 6304
rect 14599 6273 14611 6276
rect 14553 6267 14611 6273
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17512 6304 17540 6403
rect 17954 6400 17960 6412
rect 18012 6400 18018 6452
rect 21085 6443 21143 6449
rect 21085 6409 21097 6443
rect 21131 6409 21143 6443
rect 21085 6403 21143 6409
rect 21100 6372 21128 6403
rect 21174 6400 21180 6452
rect 21232 6440 21238 6452
rect 21232 6412 28580 6440
rect 21232 6400 21238 6412
rect 26329 6375 26387 6381
rect 17083 6276 17540 6304
rect 17604 6344 18460 6372
rect 21100 6344 22094 6372
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17604 6236 17632 6344
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 18322 6304 18328 6316
rect 17911 6276 18328 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 11204 6208 12388 6236
rect 16316 6208 17632 6236
rect 18049 6239 18107 6245
rect 11204 6196 11210 6208
rect 16316 6168 16344 6208
rect 18049 6205 18061 6239
rect 18095 6205 18107 6239
rect 18432 6236 18460 6344
rect 20714 6264 20720 6316
rect 20772 6304 20778 6316
rect 21269 6307 21327 6313
rect 21269 6304 21281 6307
rect 20772 6276 21281 6304
rect 20772 6264 20778 6276
rect 21269 6273 21281 6276
rect 21315 6273 21327 6307
rect 21818 6304 21824 6316
rect 21779 6276 21824 6304
rect 21269 6267 21327 6273
rect 21818 6264 21824 6276
rect 21876 6264 21882 6316
rect 22066 6313 22094 6344
rect 26329 6341 26341 6375
rect 26375 6372 26387 6375
rect 28552 6372 28580 6412
rect 29822 6400 29828 6452
rect 29880 6440 29886 6452
rect 30837 6443 30895 6449
rect 30837 6440 30849 6443
rect 29880 6412 30849 6440
rect 29880 6400 29886 6412
rect 30837 6409 30849 6412
rect 30883 6409 30895 6443
rect 30837 6403 30895 6409
rect 31205 6443 31263 6449
rect 31205 6409 31217 6443
rect 31251 6440 31263 6443
rect 31846 6440 31852 6452
rect 31251 6412 31852 6440
rect 31251 6409 31263 6412
rect 31205 6403 31263 6409
rect 31846 6400 31852 6412
rect 31904 6400 31910 6452
rect 34701 6443 34759 6449
rect 34701 6440 34713 6443
rect 31956 6412 34713 6440
rect 26375 6344 27738 6372
rect 28552 6344 31432 6372
rect 26375 6341 26387 6344
rect 26329 6335 26387 6341
rect 22066 6307 22135 6313
rect 22066 6282 22089 6307
rect 22077 6273 22089 6282
rect 22123 6273 22135 6307
rect 22077 6267 22135 6273
rect 23845 6307 23903 6313
rect 23845 6273 23857 6307
rect 23891 6273 23903 6307
rect 23845 6267 23903 6273
rect 21634 6236 21640 6248
rect 18432 6208 21640 6236
rect 18049 6199 18107 6205
rect 15488 6140 16344 6168
rect 10686 6100 10692 6112
rect 9140 6072 10692 6100
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 10778 6060 10784 6112
rect 10836 6100 10842 6112
rect 10965 6103 11023 6109
rect 10965 6100 10977 6103
rect 10836 6072 10977 6100
rect 10836 6060 10842 6072
rect 10965 6069 10977 6072
rect 11011 6069 11023 6103
rect 10965 6063 11023 6069
rect 11330 6060 11336 6112
rect 11388 6100 11394 6112
rect 11790 6100 11796 6112
rect 11388 6072 11796 6100
rect 11388 6060 11394 6072
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 13170 6060 13176 6112
rect 13228 6100 13234 6112
rect 13633 6103 13691 6109
rect 13633 6100 13645 6103
rect 13228 6072 13645 6100
rect 13228 6060 13234 6072
rect 13633 6069 13645 6072
rect 13679 6100 13691 6103
rect 15488 6100 15516 6140
rect 16758 6128 16764 6180
rect 16816 6168 16822 6180
rect 18064 6168 18092 6199
rect 21634 6196 21640 6208
rect 21692 6196 21698 6248
rect 23290 6196 23296 6248
rect 23348 6236 23354 6248
rect 23753 6239 23811 6245
rect 23753 6236 23765 6239
rect 23348 6208 23765 6236
rect 23348 6196 23354 6208
rect 23753 6205 23765 6208
rect 23799 6205 23811 6239
rect 23753 6199 23811 6205
rect 19886 6168 19892 6180
rect 16816 6140 19892 6168
rect 16816 6128 16822 6140
rect 19886 6128 19892 6140
rect 19944 6168 19950 6180
rect 21358 6168 21364 6180
rect 19944 6140 21364 6168
rect 19944 6128 19950 6140
rect 21358 6128 21364 6140
rect 21416 6128 21422 6180
rect 23860 6168 23888 6267
rect 24026 6264 24032 6316
rect 24084 6304 24090 6316
rect 26237 6307 26295 6313
rect 26237 6304 26249 6307
rect 24084 6276 26249 6304
rect 24084 6264 24090 6276
rect 26237 6273 26249 6276
rect 26283 6304 26295 6307
rect 26418 6304 26424 6316
rect 26283 6276 26424 6304
rect 26283 6273 26295 6276
rect 26237 6267 26295 6273
rect 26418 6264 26424 6276
rect 26476 6264 26482 6316
rect 26970 6304 26976 6316
rect 26931 6276 26976 6304
rect 26970 6264 26976 6276
rect 27028 6264 27034 6316
rect 29549 6307 29607 6313
rect 29549 6273 29561 6307
rect 29595 6304 29607 6307
rect 30466 6304 30472 6316
rect 29595 6276 30472 6304
rect 29595 6273 29607 6276
rect 29549 6267 29607 6273
rect 30466 6264 30472 6276
rect 30524 6264 30530 6316
rect 31294 6304 31300 6316
rect 31255 6276 31300 6304
rect 31294 6264 31300 6276
rect 31352 6264 31358 6316
rect 26878 6196 26884 6248
rect 26936 6236 26942 6248
rect 27249 6239 27307 6245
rect 27249 6236 27261 6239
rect 26936 6208 27261 6236
rect 26936 6196 26942 6208
rect 27249 6205 27261 6208
rect 27295 6205 27307 6239
rect 27249 6199 27307 6205
rect 29825 6239 29883 6245
rect 29825 6205 29837 6239
rect 29871 6236 29883 6239
rect 29914 6236 29920 6248
rect 29871 6208 29920 6236
rect 29871 6205 29883 6208
rect 29825 6199 29883 6205
rect 29914 6196 29920 6208
rect 29972 6196 29978 6248
rect 31404 6245 31432 6344
rect 31570 6332 31576 6384
rect 31628 6372 31634 6384
rect 31956 6372 31984 6412
rect 34701 6409 34713 6412
rect 34747 6409 34759 6443
rect 34701 6403 34759 6409
rect 35802 6400 35808 6452
rect 35860 6440 35866 6452
rect 35897 6443 35955 6449
rect 35897 6440 35909 6443
rect 35860 6412 35909 6440
rect 35860 6400 35866 6412
rect 35897 6409 35909 6412
rect 35943 6409 35955 6443
rect 35897 6403 35955 6409
rect 35253 6375 35311 6381
rect 35253 6372 35265 6375
rect 31628 6344 31984 6372
rect 34454 6344 35265 6372
rect 31628 6332 31634 6344
rect 35253 6341 35265 6344
rect 35299 6341 35311 6375
rect 35253 6335 35311 6341
rect 32122 6264 32128 6316
rect 32180 6304 32186 6316
rect 32309 6307 32367 6313
rect 32180 6276 32225 6304
rect 32180 6264 32186 6276
rect 32309 6273 32321 6307
rect 32355 6304 32367 6307
rect 32582 6304 32588 6316
rect 32355 6276 32588 6304
rect 32355 6273 32367 6276
rect 32309 6267 32367 6273
rect 32582 6264 32588 6276
rect 32640 6264 32646 6316
rect 32674 6264 32680 6316
rect 32732 6304 32738 6316
rect 32953 6307 33011 6313
rect 32953 6304 32965 6307
rect 32732 6276 32965 6304
rect 32732 6264 32738 6276
rect 32953 6273 32965 6276
rect 32999 6273 33011 6307
rect 32953 6267 33011 6273
rect 34514 6264 34520 6316
rect 34572 6304 34578 6316
rect 35161 6307 35219 6313
rect 35161 6304 35173 6307
rect 34572 6276 35173 6304
rect 34572 6264 34578 6276
rect 35161 6273 35173 6276
rect 35207 6304 35219 6307
rect 35710 6304 35716 6316
rect 35207 6276 35716 6304
rect 35207 6273 35219 6276
rect 35161 6267 35219 6273
rect 35710 6264 35716 6276
rect 35768 6304 35774 6316
rect 35805 6307 35863 6313
rect 35805 6304 35817 6307
rect 35768 6276 35817 6304
rect 35768 6264 35774 6276
rect 35805 6273 35817 6276
rect 35851 6273 35863 6307
rect 35805 6267 35863 6273
rect 31389 6239 31447 6245
rect 31389 6205 31401 6239
rect 31435 6205 31447 6239
rect 31389 6199 31447 6205
rect 33229 6239 33287 6245
rect 33229 6205 33241 6239
rect 33275 6236 33287 6239
rect 34698 6236 34704 6248
rect 33275 6208 34704 6236
rect 33275 6205 33287 6208
rect 33229 6199 33287 6205
rect 34698 6196 34704 6208
rect 34756 6196 34762 6248
rect 30006 6168 30012 6180
rect 23860 6140 26832 6168
rect 13679 6072 15516 6100
rect 13679 6069 13691 6072
rect 13633 6063 13691 6069
rect 15562 6060 15568 6112
rect 15620 6100 15626 6112
rect 15933 6103 15991 6109
rect 15933 6100 15945 6103
rect 15620 6072 15945 6100
rect 15620 6060 15626 6072
rect 15933 6069 15945 6072
rect 15979 6069 15991 6103
rect 16850 6100 16856 6112
rect 16811 6072 16856 6100
rect 15933 6063 15991 6069
rect 16850 6060 16856 6072
rect 16908 6060 16914 6112
rect 21082 6060 21088 6112
rect 21140 6100 21146 6112
rect 22922 6100 22928 6112
rect 21140 6072 22928 6100
rect 21140 6060 21146 6072
rect 22922 6060 22928 6072
rect 22980 6100 22986 6112
rect 23201 6103 23259 6109
rect 23201 6100 23213 6103
rect 22980 6072 23213 6100
rect 22980 6060 22986 6072
rect 23201 6069 23213 6072
rect 23247 6069 23259 6103
rect 23201 6063 23259 6069
rect 24213 6103 24271 6109
rect 24213 6069 24225 6103
rect 24259 6100 24271 6103
rect 24394 6100 24400 6112
rect 24259 6072 24400 6100
rect 24259 6069 24271 6072
rect 24213 6063 24271 6069
rect 24394 6060 24400 6072
rect 24452 6060 24458 6112
rect 26804 6100 26832 6140
rect 28644 6140 30012 6168
rect 28644 6100 28672 6140
rect 30006 6128 30012 6140
rect 30064 6128 30070 6180
rect 26804 6072 28672 6100
rect 28721 6103 28779 6109
rect 28721 6069 28733 6103
rect 28767 6100 28779 6103
rect 28994 6100 29000 6112
rect 28767 6072 29000 6100
rect 28767 6069 28779 6072
rect 28721 6063 28779 6069
rect 28994 6060 29000 6072
rect 29052 6060 29058 6112
rect 29086 6060 29092 6112
rect 29144 6100 29150 6112
rect 31110 6100 31116 6112
rect 29144 6072 31116 6100
rect 29144 6060 29150 6072
rect 31110 6060 31116 6072
rect 31168 6060 31174 6112
rect 32493 6103 32551 6109
rect 32493 6069 32505 6103
rect 32539 6100 32551 6103
rect 33594 6100 33600 6112
rect 32539 6072 33600 6100
rect 32539 6069 32551 6072
rect 32493 6063 32551 6069
rect 33594 6060 33600 6072
rect 33652 6060 33658 6112
rect 1104 6010 44896 6032
rect 1104 5958 6424 6010
rect 6476 5958 6488 6010
rect 6540 5958 6552 6010
rect 6604 5958 6616 6010
rect 6668 5958 6680 6010
rect 6732 5958 17372 6010
rect 17424 5958 17436 6010
rect 17488 5958 17500 6010
rect 17552 5958 17564 6010
rect 17616 5958 17628 6010
rect 17680 5958 28320 6010
rect 28372 5958 28384 6010
rect 28436 5958 28448 6010
rect 28500 5958 28512 6010
rect 28564 5958 28576 6010
rect 28628 5958 39268 6010
rect 39320 5958 39332 6010
rect 39384 5958 39396 6010
rect 39448 5958 39460 6010
rect 39512 5958 39524 6010
rect 39576 5958 44896 6010
rect 1104 5936 44896 5958
rect 8297 5899 8355 5905
rect 8297 5865 8309 5899
rect 8343 5896 8355 5899
rect 10042 5896 10048 5908
rect 8343 5868 10048 5896
rect 8343 5865 8355 5868
rect 8297 5859 8355 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 11701 5899 11759 5905
rect 11701 5896 11713 5899
rect 11664 5868 11713 5896
rect 11664 5856 11670 5868
rect 11701 5865 11713 5868
rect 11747 5865 11759 5899
rect 11701 5859 11759 5865
rect 11790 5856 11796 5908
rect 11848 5896 11854 5908
rect 12618 5896 12624 5908
rect 11848 5868 12624 5896
rect 11848 5856 11854 5868
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 15746 5896 15752 5908
rect 15707 5868 15752 5896
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 18322 5896 18328 5908
rect 18283 5868 18328 5896
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 23474 5856 23480 5908
rect 23532 5896 23538 5908
rect 24397 5899 24455 5905
rect 24397 5896 24409 5899
rect 23532 5868 24409 5896
rect 23532 5856 23538 5868
rect 24397 5865 24409 5868
rect 24443 5865 24455 5899
rect 26786 5896 26792 5908
rect 24397 5859 24455 5865
rect 26344 5868 26792 5896
rect 9769 5831 9827 5837
rect 9769 5797 9781 5831
rect 9815 5828 9827 5831
rect 11054 5828 11060 5840
rect 9815 5800 11060 5828
rect 9815 5797 9827 5800
rect 9769 5791 9827 5797
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 11330 5788 11336 5840
rect 11388 5828 11394 5840
rect 12805 5831 12863 5837
rect 12805 5828 12817 5831
rect 11388 5800 12817 5828
rect 11388 5788 11394 5800
rect 12805 5797 12817 5800
rect 12851 5797 12863 5831
rect 14737 5831 14795 5837
rect 14737 5828 14749 5831
rect 12805 5791 12863 5797
rect 13372 5800 14749 5828
rect 8938 5720 8944 5772
rect 8996 5760 9002 5772
rect 13372 5769 13400 5800
rect 14737 5797 14749 5800
rect 14783 5828 14795 5831
rect 16758 5828 16764 5840
rect 14783 5800 16764 5828
rect 14783 5797 14795 5800
rect 14737 5791 14795 5797
rect 16758 5788 16764 5800
rect 16816 5788 16822 5840
rect 16942 5788 16948 5840
rect 17000 5788 17006 5840
rect 13357 5763 13415 5769
rect 8996 5732 13308 5760
rect 8996 5720 9002 5732
rect 6917 5695 6975 5701
rect 6917 5661 6929 5695
rect 6963 5692 6975 5695
rect 7006 5692 7012 5704
rect 6963 5664 7012 5692
rect 6963 5661 6975 5664
rect 6917 5655 6975 5661
rect 7006 5652 7012 5664
rect 7064 5652 7070 5704
rect 9122 5692 9128 5704
rect 9083 5664 9128 5692
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 12986 5692 12992 5704
rect 10459 5664 12992 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 7184 5627 7242 5633
rect 7184 5593 7196 5627
rect 7230 5624 7242 5627
rect 8202 5624 8208 5636
rect 7230 5596 8208 5624
rect 7230 5593 7242 5596
rect 7184 5587 7242 5593
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 9968 5624 9996 5655
rect 12986 5652 12992 5664
rect 13044 5652 13050 5704
rect 13170 5692 13176 5704
rect 13131 5664 13176 5692
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 11790 5624 11796 5636
rect 9968 5596 11796 5624
rect 11790 5584 11796 5596
rect 11848 5584 11854 5636
rect 13280 5624 13308 5732
rect 13357 5729 13369 5763
rect 13403 5729 13415 5763
rect 13357 5723 13415 5729
rect 13446 5720 13452 5772
rect 13504 5760 13510 5772
rect 15381 5763 15439 5769
rect 15381 5760 15393 5763
rect 13504 5732 15393 5760
rect 13504 5720 13510 5732
rect 15381 5729 15393 5732
rect 15427 5760 15439 5763
rect 16960 5760 16988 5788
rect 15427 5732 16988 5760
rect 18340 5760 18368 5856
rect 26344 5828 26372 5868
rect 26786 5856 26792 5868
rect 26844 5856 26850 5908
rect 26878 5856 26884 5908
rect 26936 5896 26942 5908
rect 30926 5896 30932 5908
rect 26936 5868 26981 5896
rect 27080 5868 30932 5896
rect 26936 5856 26942 5868
rect 27080 5828 27108 5868
rect 30926 5856 30932 5868
rect 30984 5856 30990 5908
rect 31110 5856 31116 5908
rect 31168 5896 31174 5908
rect 34514 5896 34520 5908
rect 31168 5868 34520 5896
rect 31168 5856 31174 5868
rect 34514 5856 34520 5868
rect 34572 5856 34578 5908
rect 34698 5896 34704 5908
rect 34659 5868 34704 5896
rect 34698 5856 34704 5868
rect 34756 5856 34762 5908
rect 35342 5896 35348 5908
rect 35303 5868 35348 5896
rect 35342 5856 35348 5868
rect 35400 5856 35406 5908
rect 28350 5828 28356 5840
rect 23032 5800 26372 5828
rect 26436 5800 27108 5828
rect 27724 5800 28356 5828
rect 19337 5763 19395 5769
rect 19337 5760 19349 5763
rect 18340 5732 19349 5760
rect 15427 5729 15439 5732
rect 15381 5723 15439 5729
rect 19337 5729 19349 5732
rect 19383 5729 19395 5763
rect 19337 5723 19395 5729
rect 19797 5763 19855 5769
rect 19797 5729 19809 5763
rect 19843 5760 19855 5763
rect 20530 5760 20536 5772
rect 19843 5732 20536 5760
rect 19843 5729 19855 5732
rect 19797 5723 19855 5729
rect 20530 5720 20536 5732
rect 20588 5720 20594 5772
rect 22922 5760 22928 5772
rect 22883 5732 22928 5760
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 15562 5692 15568 5704
rect 15523 5664 15568 5692
rect 15562 5652 15568 5664
rect 15620 5652 15626 5704
rect 16945 5695 17003 5701
rect 16945 5661 16957 5695
rect 16991 5692 17003 5695
rect 17494 5692 17500 5704
rect 16991 5664 17500 5692
rect 16991 5661 17003 5664
rect 16945 5655 17003 5661
rect 17494 5652 17500 5664
rect 17552 5692 17558 5704
rect 18046 5692 18052 5704
rect 17552 5664 18052 5692
rect 17552 5652 17558 5664
rect 18046 5652 18052 5664
rect 18104 5652 18110 5704
rect 19429 5695 19487 5701
rect 19429 5661 19441 5695
rect 19475 5661 19487 5695
rect 19429 5655 19487 5661
rect 14550 5624 14556 5636
rect 13280 5596 13400 5624
rect 14511 5596 14556 5624
rect 8938 5556 8944 5568
rect 8899 5528 8944 5556
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 12710 5516 12716 5568
rect 12768 5556 12774 5568
rect 13265 5559 13323 5565
rect 13265 5556 13277 5559
rect 12768 5528 13277 5556
rect 12768 5516 12774 5528
rect 13265 5525 13277 5528
rect 13311 5525 13323 5559
rect 13372 5556 13400 5596
rect 14550 5584 14556 5596
rect 14608 5584 14614 5636
rect 16850 5584 16856 5636
rect 16908 5624 16914 5636
rect 17190 5627 17248 5633
rect 17190 5624 17202 5627
rect 16908 5596 17202 5624
rect 16908 5584 16914 5596
rect 17190 5593 17202 5596
rect 17236 5593 17248 5627
rect 19444 5624 19472 5655
rect 21726 5652 21732 5704
rect 21784 5692 21790 5704
rect 23032 5701 23060 5800
rect 23385 5763 23443 5769
rect 23385 5729 23397 5763
rect 23431 5760 23443 5763
rect 24489 5763 24547 5769
rect 24489 5760 24501 5763
rect 23431 5732 24501 5760
rect 23431 5729 23443 5732
rect 23385 5723 23443 5729
rect 24489 5729 24501 5732
rect 24535 5729 24547 5763
rect 24489 5723 24547 5729
rect 26436 5704 26464 5800
rect 27724 5760 27752 5800
rect 28350 5788 28356 5800
rect 28408 5828 28414 5840
rect 28994 5828 29000 5840
rect 28408 5800 29000 5828
rect 28408 5788 28414 5800
rect 28994 5788 29000 5800
rect 29052 5788 29058 5840
rect 29638 5788 29644 5840
rect 29696 5828 29702 5840
rect 31018 5828 31024 5840
rect 29696 5800 31024 5828
rect 29696 5788 29702 5800
rect 31018 5788 31024 5800
rect 31076 5828 31082 5840
rect 31076 5800 33640 5828
rect 31076 5788 31082 5800
rect 29733 5763 29791 5769
rect 29733 5760 29745 5763
rect 26528 5732 27752 5760
rect 21821 5695 21879 5701
rect 21821 5692 21833 5695
rect 21784 5664 21833 5692
rect 21784 5652 21790 5664
rect 21821 5661 21833 5664
rect 21867 5661 21879 5695
rect 21821 5655 21879 5661
rect 23017 5695 23075 5701
rect 23017 5661 23029 5695
rect 23063 5661 23075 5695
rect 24394 5692 24400 5704
rect 24355 5664 24400 5692
rect 23017 5655 23075 5661
rect 24394 5652 24400 5664
rect 24452 5652 24458 5704
rect 24670 5692 24676 5704
rect 24631 5664 24676 5692
rect 24670 5652 24676 5664
rect 24728 5652 24734 5704
rect 26418 5692 26424 5704
rect 26379 5664 26424 5692
rect 26418 5652 26424 5664
rect 26476 5652 26482 5704
rect 26528 5624 26556 5732
rect 27065 5695 27123 5701
rect 27065 5661 27077 5695
rect 27111 5692 27123 5695
rect 27614 5692 27620 5704
rect 27111 5664 27620 5692
rect 27111 5661 27123 5664
rect 27065 5655 27123 5661
rect 27614 5652 27620 5664
rect 27672 5652 27678 5704
rect 27724 5701 27752 5732
rect 28736 5732 29745 5760
rect 27709 5695 27767 5701
rect 27709 5661 27721 5695
rect 27755 5661 27767 5695
rect 27709 5655 27767 5661
rect 27798 5652 27804 5704
rect 27856 5692 27862 5704
rect 27856 5664 27901 5692
rect 27856 5652 27862 5664
rect 28350 5652 28356 5704
rect 28408 5692 28414 5704
rect 28736 5701 28764 5732
rect 29733 5729 29745 5732
rect 29779 5760 29791 5763
rect 29779 5732 31754 5760
rect 29779 5729 29791 5732
rect 29733 5723 29791 5729
rect 28445 5695 28503 5701
rect 28445 5692 28457 5695
rect 28408 5664 28457 5692
rect 28408 5652 28414 5664
rect 28445 5661 28457 5664
rect 28491 5661 28503 5695
rect 28445 5655 28503 5661
rect 28721 5695 28779 5701
rect 28721 5661 28733 5695
rect 28767 5661 28779 5695
rect 28721 5655 28779 5661
rect 19444 5596 26556 5624
rect 27525 5627 27583 5633
rect 17190 5587 17248 5593
rect 27525 5593 27537 5627
rect 27571 5624 27583 5627
rect 28736 5624 28764 5655
rect 28994 5652 29000 5704
rect 29052 5692 29058 5704
rect 29822 5692 29828 5704
rect 29052 5664 29828 5692
rect 29052 5652 29058 5664
rect 29822 5652 29828 5664
rect 29880 5652 29886 5704
rect 29917 5695 29975 5701
rect 29917 5661 29929 5695
rect 29963 5661 29975 5695
rect 29917 5655 29975 5661
rect 29638 5624 29644 5636
rect 27571 5596 28764 5624
rect 29472 5596 29644 5624
rect 27571 5593 27583 5596
rect 27525 5587 27583 5593
rect 21174 5556 21180 5568
rect 13372 5528 21180 5556
rect 13265 5519 13323 5525
rect 21174 5516 21180 5528
rect 21232 5516 21238 5568
rect 22005 5559 22063 5565
rect 22005 5525 22017 5559
rect 22051 5556 22063 5559
rect 24026 5556 24032 5568
rect 22051 5528 24032 5556
rect 22051 5525 22063 5528
rect 22005 5519 22063 5525
rect 24026 5516 24032 5528
rect 24084 5516 24090 5568
rect 24302 5516 24308 5568
rect 24360 5556 24366 5568
rect 24857 5559 24915 5565
rect 24857 5556 24869 5559
rect 24360 5528 24869 5556
rect 24360 5516 24366 5528
rect 24857 5525 24869 5528
rect 24903 5525 24915 5559
rect 24857 5519 24915 5525
rect 26237 5559 26295 5565
rect 26237 5525 26249 5559
rect 26283 5556 26295 5559
rect 27540 5556 27568 5587
rect 26283 5528 27568 5556
rect 27801 5559 27859 5565
rect 26283 5525 26295 5528
rect 26237 5519 26295 5525
rect 27801 5525 27813 5559
rect 27847 5556 27859 5559
rect 28166 5556 28172 5568
rect 27847 5528 28172 5556
rect 27847 5525 27859 5528
rect 27801 5519 27859 5525
rect 28166 5516 28172 5528
rect 28224 5516 28230 5568
rect 28261 5559 28319 5565
rect 28261 5525 28273 5559
rect 28307 5556 28319 5559
rect 28534 5556 28540 5568
rect 28307 5528 28540 5556
rect 28307 5525 28319 5528
rect 28261 5519 28319 5525
rect 28534 5516 28540 5528
rect 28592 5516 28598 5568
rect 28626 5516 28632 5568
rect 28684 5556 28690 5568
rect 29472 5556 29500 5596
rect 29638 5584 29644 5596
rect 29696 5624 29702 5636
rect 29932 5624 29960 5655
rect 30006 5652 30012 5704
rect 30064 5692 30070 5704
rect 30064 5664 30109 5692
rect 30064 5652 30070 5664
rect 30374 5652 30380 5704
rect 30432 5692 30438 5704
rect 31205 5695 31263 5701
rect 31205 5692 31217 5695
rect 30432 5664 31217 5692
rect 30432 5652 30438 5664
rect 31205 5661 31217 5664
rect 31251 5661 31263 5695
rect 31726 5692 31754 5732
rect 32674 5720 32680 5772
rect 32732 5760 32738 5772
rect 32769 5763 32827 5769
rect 32769 5760 32781 5763
rect 32732 5732 32781 5760
rect 32732 5720 32738 5732
rect 32769 5729 32781 5732
rect 32815 5729 32827 5763
rect 32769 5723 32827 5729
rect 32122 5692 32128 5704
rect 31726 5664 32128 5692
rect 31205 5655 31263 5661
rect 32122 5652 32128 5664
rect 32180 5692 32186 5704
rect 33612 5701 33640 5800
rect 33686 5720 33692 5772
rect 33744 5760 33750 5772
rect 33744 5732 35572 5760
rect 33744 5720 33750 5732
rect 35544 5701 35572 5732
rect 33413 5695 33471 5701
rect 33413 5692 33425 5695
rect 32180 5664 33425 5692
rect 32180 5652 32186 5664
rect 33413 5661 33425 5664
rect 33459 5661 33471 5695
rect 33413 5655 33471 5661
rect 33597 5695 33655 5701
rect 33597 5661 33609 5695
rect 33643 5661 33655 5695
rect 33597 5655 33655 5661
rect 34885 5695 34943 5701
rect 34885 5661 34897 5695
rect 34931 5661 34943 5695
rect 34885 5655 34943 5661
rect 35529 5695 35587 5701
rect 35529 5661 35541 5695
rect 35575 5661 35587 5695
rect 35529 5655 35587 5661
rect 29696 5596 29960 5624
rect 30024 5624 30052 5652
rect 30742 5624 30748 5636
rect 30024 5596 30748 5624
rect 29696 5584 29702 5596
rect 30742 5584 30748 5596
rect 30800 5624 30806 5636
rect 31570 5624 31576 5636
rect 30800 5596 31576 5624
rect 30800 5584 30806 5596
rect 31570 5584 31576 5596
rect 31628 5584 31634 5636
rect 33134 5584 33140 5636
rect 33192 5624 33198 5636
rect 34900 5624 34928 5655
rect 35618 5652 35624 5704
rect 35676 5692 35682 5704
rect 36173 5695 36231 5701
rect 36173 5692 36185 5695
rect 35676 5664 36185 5692
rect 35676 5652 35682 5664
rect 36173 5661 36185 5664
rect 36219 5661 36231 5695
rect 43898 5692 43904 5704
rect 43859 5664 43904 5692
rect 36173 5655 36231 5661
rect 43898 5652 43904 5664
rect 43956 5652 43962 5704
rect 33192 5596 34928 5624
rect 33192 5584 33198 5596
rect 28684 5528 29500 5556
rect 29549 5559 29607 5565
rect 28684 5516 28690 5528
rect 29549 5525 29561 5559
rect 29595 5556 29607 5559
rect 31386 5556 31392 5568
rect 29595 5528 31392 5556
rect 29595 5525 29607 5528
rect 29549 5519 29607 5525
rect 31386 5516 31392 5528
rect 31444 5516 31450 5568
rect 33502 5556 33508 5568
rect 33463 5528 33508 5556
rect 33502 5516 33508 5528
rect 33560 5516 33566 5568
rect 35434 5516 35440 5568
rect 35492 5556 35498 5568
rect 35989 5559 36047 5565
rect 35989 5556 36001 5559
rect 35492 5528 36001 5556
rect 35492 5516 35498 5528
rect 35989 5525 36001 5528
rect 36035 5525 36047 5559
rect 44082 5556 44088 5568
rect 44043 5528 44088 5556
rect 35989 5519 36047 5525
rect 44082 5516 44088 5528
rect 44140 5516 44146 5568
rect 1104 5466 45056 5488
rect 1104 5414 11898 5466
rect 11950 5414 11962 5466
rect 12014 5414 12026 5466
rect 12078 5414 12090 5466
rect 12142 5414 12154 5466
rect 12206 5414 22846 5466
rect 22898 5414 22910 5466
rect 22962 5414 22974 5466
rect 23026 5414 23038 5466
rect 23090 5414 23102 5466
rect 23154 5414 33794 5466
rect 33846 5414 33858 5466
rect 33910 5414 33922 5466
rect 33974 5414 33986 5466
rect 34038 5414 34050 5466
rect 34102 5414 44742 5466
rect 44794 5414 44806 5466
rect 44858 5414 44870 5466
rect 44922 5414 44934 5466
rect 44986 5414 44998 5466
rect 45050 5414 45056 5466
rect 1104 5392 45056 5414
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 10965 5355 11023 5361
rect 10965 5352 10977 5355
rect 10744 5324 10977 5352
rect 10744 5312 10750 5324
rect 10965 5321 10977 5324
rect 11011 5321 11023 5355
rect 11790 5352 11796 5364
rect 11751 5324 11796 5352
rect 10965 5315 11023 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 12250 5352 12256 5364
rect 12211 5324 12256 5352
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 13630 5312 13636 5364
rect 13688 5352 13694 5364
rect 18785 5355 18843 5361
rect 13688 5324 18736 5352
rect 13688 5312 13694 5324
rect 8012 5287 8070 5293
rect 8012 5253 8024 5287
rect 8058 5284 8070 5287
rect 8938 5284 8944 5296
rect 8058 5256 8944 5284
rect 8058 5253 8070 5256
rect 8012 5247 8070 5253
rect 8938 5244 8944 5256
rect 8996 5244 9002 5296
rect 11330 5284 11336 5296
rect 10152 5256 11336 5284
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 10152 5225 10180 5256
rect 11330 5244 11336 5256
rect 11388 5244 11394 5296
rect 12986 5284 12992 5296
rect 12947 5256 12992 5284
rect 12986 5244 12992 5256
rect 13044 5244 13050 5296
rect 16022 5284 16028 5296
rect 14200 5256 16028 5284
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7064 5188 7757 5216
rect 7064 5176 7070 5188
rect 7745 5185 7757 5188
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5185 10195 5219
rect 10778 5216 10784 5228
rect 10739 5188 10784 5216
rect 10137 5179 10195 5185
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5216 12219 5219
rect 14200 5216 14228 5256
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 17672 5287 17730 5293
rect 17672 5253 17684 5287
rect 17718 5284 17730 5287
rect 17770 5284 17776 5296
rect 17718 5256 17776 5284
rect 17718 5253 17730 5256
rect 17672 5247 17730 5253
rect 17770 5244 17776 5256
rect 17828 5244 17834 5296
rect 18708 5284 18736 5324
rect 18785 5321 18797 5355
rect 18831 5352 18843 5355
rect 19334 5352 19340 5364
rect 18831 5324 19340 5352
rect 18831 5321 18843 5324
rect 18785 5315 18843 5321
rect 19334 5312 19340 5324
rect 19392 5352 19398 5364
rect 19613 5355 19671 5361
rect 19613 5352 19625 5355
rect 19392 5324 19625 5352
rect 19392 5312 19398 5324
rect 19613 5321 19625 5324
rect 19659 5321 19671 5355
rect 19613 5315 19671 5321
rect 19705 5355 19763 5361
rect 19705 5321 19717 5355
rect 19751 5352 19763 5355
rect 19794 5352 19800 5364
rect 19751 5324 19800 5352
rect 19751 5321 19763 5324
rect 19705 5315 19763 5321
rect 19794 5312 19800 5324
rect 19852 5312 19858 5364
rect 19904 5324 41414 5352
rect 19904 5284 19932 5324
rect 23937 5287 23995 5293
rect 18708 5256 19932 5284
rect 22112 5256 23796 5284
rect 12207 5188 14228 5216
rect 12207 5185 12219 5188
rect 12161 5179 12219 5185
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 15381 5219 15439 5225
rect 15381 5216 15393 5219
rect 14884 5188 15393 5216
rect 14884 5176 14890 5188
rect 15381 5185 15393 5188
rect 15427 5185 15439 5219
rect 15381 5179 15439 5185
rect 17218 5176 17224 5228
rect 17276 5216 17282 5228
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 17276 5188 17417 5216
rect 17276 5176 17282 5188
rect 17405 5185 17417 5188
rect 17451 5216 17463 5219
rect 17494 5216 17500 5228
rect 17451 5188 17500 5216
rect 17451 5185 17463 5188
rect 17405 5179 17463 5185
rect 17494 5176 17500 5188
rect 17552 5176 17558 5228
rect 20438 5216 20444 5228
rect 20399 5188 20444 5216
rect 20438 5176 20444 5188
rect 20496 5176 20502 5228
rect 20714 5216 20720 5228
rect 20675 5188 20720 5216
rect 20714 5176 20720 5188
rect 20772 5176 20778 5228
rect 22112 5225 22140 5256
rect 22097 5219 22155 5225
rect 22097 5185 22109 5219
rect 22143 5185 22155 5219
rect 23106 5216 23112 5228
rect 23067 5188 23112 5216
rect 22097 5179 22155 5185
rect 23106 5176 23112 5188
rect 23164 5176 23170 5228
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5148 1731 5151
rect 6270 5148 6276 5160
rect 1719 5120 6276 5148
rect 1719 5117 1731 5120
rect 1673 5111 1731 5117
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 9858 5108 9864 5160
rect 9916 5148 9922 5160
rect 10597 5151 10655 5157
rect 10597 5148 10609 5151
rect 9916 5120 10609 5148
rect 9916 5108 9922 5120
rect 10597 5117 10609 5120
rect 10643 5148 10655 5151
rect 12342 5148 12348 5160
rect 10643 5120 12204 5148
rect 12303 5120 12348 5148
rect 10643 5117 10655 5120
rect 10597 5111 10655 5117
rect 9953 5083 10011 5089
rect 9953 5049 9965 5083
rect 9999 5080 10011 5083
rect 11146 5080 11152 5092
rect 9999 5052 11152 5080
rect 9999 5049 10011 5052
rect 9953 5043 10011 5049
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 12176 5080 12204 5120
rect 12342 5108 12348 5120
rect 12400 5108 12406 5160
rect 14734 5148 14740 5160
rect 14647 5120 14740 5148
rect 14734 5108 14740 5120
rect 14792 5148 14798 5160
rect 15746 5148 15752 5160
rect 14792 5120 15752 5148
rect 14792 5108 14798 5120
rect 15746 5108 15752 5120
rect 15804 5148 15810 5160
rect 17236 5148 17264 5176
rect 19886 5148 19892 5160
rect 15804 5120 17264 5148
rect 19847 5120 19892 5148
rect 15804 5108 15810 5120
rect 19886 5108 19892 5120
rect 19944 5108 19950 5160
rect 20530 5148 20536 5160
rect 20491 5120 20536 5148
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 22189 5151 22247 5157
rect 22189 5117 22201 5151
rect 22235 5148 22247 5151
rect 22278 5148 22284 5160
rect 22235 5120 22284 5148
rect 22235 5117 22247 5120
rect 22189 5111 22247 5117
rect 22278 5108 22284 5120
rect 22336 5108 22342 5160
rect 23017 5151 23075 5157
rect 23017 5148 23029 5151
rect 22388 5120 23029 5148
rect 13446 5080 13452 5092
rect 12176 5052 13452 5080
rect 13446 5040 13452 5052
rect 13504 5040 13510 5092
rect 21634 5040 21640 5092
rect 21692 5080 21698 5092
rect 22388 5080 22416 5120
rect 23017 5117 23029 5120
rect 23063 5117 23075 5151
rect 23474 5148 23480 5160
rect 23435 5120 23480 5148
rect 23017 5111 23075 5117
rect 23474 5108 23480 5120
rect 23532 5108 23538 5160
rect 23768 5148 23796 5256
rect 23937 5253 23949 5287
rect 23983 5284 23995 5287
rect 25409 5287 25467 5293
rect 23983 5256 25084 5284
rect 23983 5253 23995 5256
rect 23937 5247 23995 5253
rect 25056 5228 25084 5256
rect 25409 5253 25421 5287
rect 25455 5284 25467 5287
rect 27522 5284 27528 5296
rect 25455 5256 27528 5284
rect 25455 5253 25467 5256
rect 25409 5247 25467 5253
rect 27522 5244 27528 5256
rect 27580 5284 27586 5296
rect 27985 5287 28043 5293
rect 27985 5284 27997 5287
rect 27580 5256 27997 5284
rect 27580 5244 27586 5256
rect 27985 5253 27997 5256
rect 28031 5253 28043 5287
rect 28442 5284 28448 5296
rect 28403 5256 28448 5284
rect 27985 5247 28043 5253
rect 28442 5244 28448 5256
rect 28500 5244 28506 5296
rect 28534 5244 28540 5296
rect 28592 5284 28598 5296
rect 28645 5287 28703 5293
rect 28645 5284 28657 5287
rect 28592 5256 28657 5284
rect 28592 5244 28598 5256
rect 28645 5253 28657 5256
rect 28691 5253 28703 5287
rect 28645 5247 28703 5253
rect 30466 5244 30472 5296
rect 30524 5284 30530 5296
rect 30561 5287 30619 5293
rect 30561 5284 30573 5287
rect 30524 5256 30573 5284
rect 30524 5244 30530 5256
rect 30561 5253 30573 5256
rect 30607 5253 30619 5287
rect 30837 5287 30895 5293
rect 30837 5284 30849 5287
rect 30561 5247 30619 5253
rect 30668 5256 30849 5284
rect 23842 5176 23848 5228
rect 23900 5216 23906 5228
rect 24121 5219 24179 5225
rect 24121 5216 24133 5219
rect 23900 5188 24133 5216
rect 23900 5176 23906 5188
rect 24121 5185 24133 5188
rect 24167 5185 24179 5219
rect 25038 5216 25044 5228
rect 24951 5188 25044 5216
rect 24121 5179 24179 5185
rect 25038 5176 25044 5188
rect 25096 5176 25102 5228
rect 25130 5176 25136 5228
rect 25188 5216 25194 5228
rect 25314 5216 25320 5228
rect 25188 5188 25233 5216
rect 25275 5188 25320 5216
rect 25188 5176 25194 5188
rect 25314 5176 25320 5188
rect 25372 5176 25378 5228
rect 25498 5176 25504 5228
rect 25556 5216 25562 5228
rect 27065 5219 27123 5225
rect 27065 5216 27077 5219
rect 25556 5188 27077 5216
rect 25556 5176 25562 5188
rect 27065 5185 27077 5188
rect 27111 5185 27123 5219
rect 27065 5179 27123 5185
rect 27249 5219 27307 5225
rect 27249 5185 27261 5219
rect 27295 5216 27307 5219
rect 27338 5216 27344 5228
rect 27295 5188 27344 5216
rect 27295 5185 27307 5188
rect 27249 5179 27307 5185
rect 27338 5176 27344 5188
rect 27396 5216 27402 5228
rect 27801 5219 27859 5225
rect 27801 5216 27813 5219
rect 27396 5188 27813 5216
rect 27396 5176 27402 5188
rect 27801 5185 27813 5188
rect 27847 5216 27859 5219
rect 27847 5188 29684 5216
rect 27847 5185 27859 5188
rect 27801 5179 27859 5185
rect 24854 5148 24860 5160
rect 23768 5120 24860 5148
rect 24854 5108 24860 5120
rect 24912 5108 24918 5160
rect 27157 5151 27215 5157
rect 27157 5117 27169 5151
rect 27203 5148 27215 5151
rect 28442 5148 28448 5160
rect 27203 5120 28448 5148
rect 27203 5117 27215 5120
rect 27157 5111 27215 5117
rect 28442 5108 28448 5120
rect 28500 5148 28506 5160
rect 29270 5148 29276 5160
rect 28500 5120 29276 5148
rect 28500 5108 28506 5120
rect 29270 5108 29276 5120
rect 29328 5108 29334 5160
rect 29362 5108 29368 5160
rect 29420 5148 29426 5160
rect 29549 5151 29607 5157
rect 29549 5148 29561 5151
rect 29420 5120 29561 5148
rect 29420 5108 29426 5120
rect 29549 5117 29561 5120
rect 29595 5117 29607 5151
rect 29656 5148 29684 5188
rect 29822 5176 29828 5228
rect 29880 5216 29886 5228
rect 30668 5216 30696 5256
rect 30837 5253 30849 5256
rect 30883 5253 30895 5287
rect 30837 5247 30895 5253
rect 30926 5244 30932 5296
rect 30984 5284 30990 5296
rect 31113 5287 31171 5293
rect 30984 5256 31029 5284
rect 30984 5244 30990 5256
rect 31113 5253 31125 5287
rect 31159 5284 31171 5287
rect 31754 5284 31760 5296
rect 31159 5256 31760 5284
rect 31159 5253 31171 5256
rect 31113 5247 31171 5253
rect 31754 5244 31760 5256
rect 31812 5284 31818 5296
rect 31938 5284 31944 5296
rect 31812 5256 31944 5284
rect 31812 5244 31818 5256
rect 31938 5244 31944 5256
rect 31996 5244 32002 5296
rect 32309 5287 32367 5293
rect 32309 5284 32321 5287
rect 32048 5256 32321 5284
rect 29880 5188 30696 5216
rect 29880 5176 29886 5188
rect 30742 5176 30748 5228
rect 30800 5216 30806 5228
rect 32048 5216 32076 5256
rect 32309 5253 32321 5256
rect 32355 5253 32367 5287
rect 35805 5287 35863 5293
rect 35805 5284 35817 5287
rect 34914 5256 35817 5284
rect 32309 5247 32367 5253
rect 35805 5253 35817 5256
rect 35851 5253 35863 5287
rect 35805 5247 35863 5253
rect 30800 5188 30845 5216
rect 31726 5188 32076 5216
rect 30800 5176 30806 5188
rect 29914 5148 29920 5160
rect 29656 5120 29920 5148
rect 29549 5111 29607 5117
rect 29914 5108 29920 5120
rect 29972 5148 29978 5160
rect 31726 5148 31754 5188
rect 32122 5176 32128 5228
rect 32180 5216 32186 5228
rect 32180 5188 32225 5216
rect 32180 5176 32186 5188
rect 32674 5176 32680 5228
rect 32732 5216 32738 5228
rect 33413 5219 33471 5225
rect 33413 5216 33425 5219
rect 32732 5188 33425 5216
rect 32732 5176 32738 5188
rect 33413 5185 33425 5188
rect 33459 5185 33471 5219
rect 35710 5216 35716 5228
rect 35671 5188 35716 5216
rect 33413 5179 33471 5185
rect 35710 5176 35716 5188
rect 35768 5176 35774 5228
rect 41386 5216 41414 5324
rect 42981 5219 43039 5225
rect 42981 5216 42993 5219
rect 41386 5188 42993 5216
rect 42981 5185 42993 5188
rect 43027 5216 43039 5219
rect 43257 5219 43315 5225
rect 43257 5216 43269 5219
rect 43027 5188 43269 5216
rect 43027 5185 43039 5188
rect 42981 5179 43039 5185
rect 43257 5185 43269 5188
rect 43303 5185 43315 5219
rect 43257 5179 43315 5185
rect 29972 5120 31754 5148
rect 33689 5151 33747 5157
rect 29972 5108 29978 5120
rect 33689 5117 33701 5151
rect 33735 5148 33747 5151
rect 35434 5148 35440 5160
rect 33735 5120 35440 5148
rect 33735 5117 33747 5120
rect 33689 5111 33747 5117
rect 35434 5108 35440 5120
rect 35492 5108 35498 5160
rect 21692 5052 22416 5080
rect 22465 5083 22523 5089
rect 21692 5040 21698 5052
rect 22465 5049 22477 5083
rect 22511 5080 22523 5083
rect 24670 5080 24676 5092
rect 22511 5052 24676 5080
rect 22511 5049 22523 5052
rect 22465 5043 22523 5049
rect 24670 5040 24676 5052
rect 24728 5040 24734 5092
rect 27614 5040 27620 5092
rect 27672 5080 27678 5092
rect 28813 5083 28871 5089
rect 28813 5080 28825 5083
rect 27672 5052 28825 5080
rect 27672 5040 27678 5052
rect 28813 5049 28825 5052
rect 28859 5049 28871 5083
rect 28813 5043 28871 5049
rect 30926 5040 30932 5092
rect 30984 5080 30990 5092
rect 33318 5080 33324 5092
rect 30984 5052 33324 5080
rect 30984 5040 30990 5052
rect 33318 5040 33324 5052
rect 33376 5040 33382 5092
rect 9122 5012 9128 5024
rect 9083 4984 9128 5012
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 15010 4972 15016 5024
rect 15068 5012 15074 5024
rect 15197 5015 15255 5021
rect 15197 5012 15209 5015
rect 15068 4984 15209 5012
rect 15068 4972 15074 4984
rect 15197 4981 15209 4984
rect 15243 4981 15255 5015
rect 15197 4975 15255 4981
rect 18046 4972 18052 5024
rect 18104 5012 18110 5024
rect 19245 5015 19303 5021
rect 19245 5012 19257 5015
rect 18104 4984 19257 5012
rect 18104 4972 18110 4984
rect 19245 4981 19257 4984
rect 19291 4981 19303 5015
rect 19245 4975 19303 4981
rect 19426 4972 19432 5024
rect 19484 5012 19490 5024
rect 20441 5015 20499 5021
rect 20441 5012 20453 5015
rect 19484 4984 20453 5012
rect 19484 4972 19490 4984
rect 20441 4981 20453 4984
rect 20487 4981 20499 5015
rect 20441 4975 20499 4981
rect 20901 5015 20959 5021
rect 20901 4981 20913 5015
rect 20947 5012 20959 5015
rect 22738 5012 22744 5024
rect 20947 4984 22744 5012
rect 20947 4981 20959 4984
rect 20901 4975 20959 4981
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 23566 4972 23572 5024
rect 23624 5012 23630 5024
rect 24305 5015 24363 5021
rect 24305 5012 24317 5015
rect 23624 4984 24317 5012
rect 23624 4972 23630 4984
rect 24305 4981 24317 4984
rect 24351 4981 24363 5015
rect 24305 4975 24363 4981
rect 24394 4972 24400 5024
rect 24452 5012 24458 5024
rect 25041 5015 25099 5021
rect 25041 5012 25053 5015
rect 24452 4984 25053 5012
rect 24452 4972 24458 4984
rect 25041 4981 25053 4984
rect 25087 4981 25099 5015
rect 25041 4975 25099 4981
rect 28166 4972 28172 5024
rect 28224 5012 28230 5024
rect 28629 5015 28687 5021
rect 28629 5012 28641 5015
rect 28224 4984 28641 5012
rect 28224 4972 28230 4984
rect 28629 4981 28641 4984
rect 28675 4981 28687 5015
rect 28629 4975 28687 4981
rect 31938 4972 31944 5024
rect 31996 5012 32002 5024
rect 32493 5015 32551 5021
rect 32493 5012 32505 5015
rect 31996 4984 32505 5012
rect 31996 4972 32002 4984
rect 32493 4981 32505 4984
rect 32539 4981 32551 5015
rect 32493 4975 32551 4981
rect 32582 4972 32588 5024
rect 32640 5012 32646 5024
rect 35161 5015 35219 5021
rect 35161 5012 35173 5015
rect 32640 4984 35173 5012
rect 32640 4972 32646 4984
rect 35161 4981 35173 4984
rect 35207 4981 35219 5015
rect 42794 5012 42800 5024
rect 42755 4984 42800 5012
rect 35161 4975 35219 4981
rect 42794 4972 42800 4984
rect 42852 4972 42858 5024
rect 1104 4922 44896 4944
rect 1104 4870 6424 4922
rect 6476 4870 6488 4922
rect 6540 4870 6552 4922
rect 6604 4870 6616 4922
rect 6668 4870 6680 4922
rect 6732 4870 17372 4922
rect 17424 4870 17436 4922
rect 17488 4870 17500 4922
rect 17552 4870 17564 4922
rect 17616 4870 17628 4922
rect 17680 4870 28320 4922
rect 28372 4870 28384 4922
rect 28436 4870 28448 4922
rect 28500 4870 28512 4922
rect 28564 4870 28576 4922
rect 28628 4870 39268 4922
rect 39320 4870 39332 4922
rect 39384 4870 39396 4922
rect 39448 4870 39460 4922
rect 39512 4870 39524 4922
rect 39576 4870 44896 4922
rect 1104 4848 44896 4870
rect 11698 4768 11704 4820
rect 11756 4808 11762 4820
rect 12342 4808 12348 4820
rect 11756 4780 12348 4808
rect 11756 4768 11762 4780
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 14090 4808 14096 4820
rect 14051 4780 14096 4808
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 17497 4811 17555 4817
rect 17497 4777 17509 4811
rect 17543 4808 17555 4811
rect 17770 4808 17776 4820
rect 17543 4780 17776 4808
rect 17543 4777 17555 4780
rect 17497 4771 17555 4777
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 19797 4811 19855 4817
rect 19797 4777 19809 4811
rect 19843 4808 19855 4811
rect 20438 4808 20444 4820
rect 19843 4780 20444 4808
rect 19843 4777 19855 4780
rect 19797 4771 19855 4777
rect 20438 4768 20444 4780
rect 20496 4768 20502 4820
rect 22084 4811 22142 4817
rect 22084 4777 22096 4811
rect 22130 4808 22142 4811
rect 24394 4808 24400 4820
rect 22130 4780 24400 4808
rect 22130 4777 22142 4780
rect 22084 4771 22142 4777
rect 24394 4768 24400 4780
rect 24452 4768 24458 4820
rect 24854 4808 24860 4820
rect 24815 4780 24860 4808
rect 24854 4768 24860 4780
rect 24912 4768 24918 4820
rect 25038 4808 25044 4820
rect 24999 4780 25044 4808
rect 25038 4768 25044 4780
rect 25096 4768 25102 4820
rect 25130 4768 25136 4820
rect 25188 4808 25194 4820
rect 25593 4811 25651 4817
rect 25593 4808 25605 4811
rect 25188 4780 25605 4808
rect 25188 4768 25194 4780
rect 25593 4777 25605 4780
rect 25639 4777 25651 4811
rect 25593 4771 25651 4777
rect 26142 4768 26148 4820
rect 26200 4808 26206 4820
rect 26789 4811 26847 4817
rect 26789 4808 26801 4811
rect 26200 4780 26801 4808
rect 26200 4768 26206 4780
rect 26789 4777 26801 4780
rect 26835 4777 26847 4811
rect 26789 4771 26847 4777
rect 26878 4768 26884 4820
rect 26936 4808 26942 4820
rect 28629 4811 28687 4817
rect 28629 4808 28641 4811
rect 26936 4780 28641 4808
rect 26936 4768 26942 4780
rect 28629 4777 28641 4780
rect 28675 4808 28687 4811
rect 29086 4808 29092 4820
rect 28675 4780 29092 4808
rect 28675 4777 28687 4780
rect 28629 4771 28687 4777
rect 29086 4768 29092 4780
rect 29144 4768 29150 4820
rect 29454 4768 29460 4820
rect 29512 4808 29518 4820
rect 31297 4811 31355 4817
rect 31297 4808 31309 4811
rect 29512 4780 31309 4808
rect 29512 4768 29518 4780
rect 31297 4777 31309 4780
rect 31343 4777 31355 4811
rect 31297 4771 31355 4777
rect 31941 4811 31999 4817
rect 31941 4777 31953 4811
rect 31987 4777 31999 4811
rect 31941 4771 31999 4777
rect 32125 4811 32183 4817
rect 32125 4777 32137 4811
rect 32171 4808 32183 4811
rect 32766 4808 32772 4820
rect 32171 4780 32628 4808
rect 32727 4780 32772 4808
rect 32171 4777 32183 4780
rect 32125 4771 32183 4777
rect 10321 4743 10379 4749
rect 10321 4709 10333 4743
rect 10367 4740 10379 4743
rect 11790 4740 11796 4752
rect 10367 4712 11796 4740
rect 10367 4709 10379 4712
rect 10321 4703 10379 4709
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 18693 4743 18751 4749
rect 18693 4709 18705 4743
rect 18739 4740 18751 4743
rect 20714 4740 20720 4752
rect 18739 4712 20720 4740
rect 18739 4709 18751 4712
rect 18693 4703 18751 4709
rect 20714 4700 20720 4712
rect 20772 4700 20778 4752
rect 29270 4700 29276 4752
rect 29328 4740 29334 4752
rect 31956 4740 31984 4771
rect 32600 4740 32628 4780
rect 32766 4768 32772 4780
rect 32824 4768 32830 4820
rect 32953 4811 33011 4817
rect 32953 4777 32965 4811
rect 32999 4808 33011 4811
rect 33134 4808 33140 4820
rect 32999 4780 33140 4808
rect 32999 4777 33011 4780
rect 32953 4771 33011 4777
rect 33134 4768 33140 4780
rect 33192 4768 33198 4820
rect 33226 4768 33232 4820
rect 33284 4808 33290 4820
rect 33597 4811 33655 4817
rect 33597 4808 33609 4811
rect 33284 4780 33609 4808
rect 33284 4768 33290 4780
rect 33597 4777 33609 4780
rect 33643 4777 33655 4811
rect 33597 4771 33655 4777
rect 33781 4811 33839 4817
rect 33781 4777 33793 4811
rect 33827 4808 33839 4811
rect 35618 4808 35624 4820
rect 33827 4780 35624 4808
rect 33827 4777 33839 4780
rect 33781 4771 33839 4777
rect 35618 4768 35624 4780
rect 35676 4768 35682 4820
rect 33686 4740 33692 4752
rect 29328 4712 29684 4740
rect 31956 4712 32260 4740
rect 32600 4712 33692 4740
rect 29328 4700 29334 4712
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 9180 4644 11529 4672
rect 9180 4632 9186 4644
rect 11517 4641 11529 4644
rect 11563 4641 11575 4675
rect 11517 4635 11575 4641
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4604 10563 4607
rect 11422 4604 11428 4616
rect 10551 4576 11428 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 11532 4604 11560 4635
rect 11606 4632 11612 4684
rect 11664 4672 11670 4684
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 11664 4644 12173 4672
rect 11664 4632 11670 4644
rect 12161 4641 12173 4644
rect 12207 4641 12219 4675
rect 14734 4672 14740 4684
rect 14695 4644 14740 4672
rect 12161 4635 12219 4641
rect 14734 4632 14740 4644
rect 14792 4632 14798 4684
rect 18233 4675 18291 4681
rect 18233 4641 18245 4675
rect 18279 4641 18291 4675
rect 19334 4672 19340 4684
rect 19295 4644 19340 4672
rect 18233 4635 18291 4641
rect 12710 4604 12716 4616
rect 11532 4576 12716 4604
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 15010 4613 15016 4616
rect 15004 4604 15016 4613
rect 14971 4576 15016 4604
rect 15004 4567 15016 4576
rect 15010 4564 15016 4567
rect 15068 4564 15074 4616
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4604 17739 4607
rect 18046 4604 18052 4616
rect 17727 4576 18052 4604
rect 17727 4573 17739 4576
rect 17681 4567 17739 4573
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 6270 4496 6276 4548
rect 6328 4536 6334 4548
rect 12434 4545 12440 4548
rect 11333 4539 11391 4545
rect 6328 4508 11284 4536
rect 6328 4496 6334 4508
rect 10965 4471 11023 4477
rect 10965 4437 10977 4471
rect 11011 4468 11023 4471
rect 11146 4468 11152 4480
rect 11011 4440 11152 4468
rect 11011 4437 11023 4440
rect 10965 4431 11023 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 11256 4468 11284 4508
rect 11333 4505 11345 4539
rect 11379 4536 11391 4539
rect 11379 4508 11928 4536
rect 11379 4505 11391 4508
rect 11333 4499 11391 4505
rect 11425 4471 11483 4477
rect 11425 4468 11437 4471
rect 11256 4440 11437 4468
rect 11425 4437 11437 4440
rect 11471 4468 11483 4471
rect 11698 4468 11704 4480
rect 11471 4440 11704 4468
rect 11471 4437 11483 4440
rect 11425 4431 11483 4437
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 11900 4468 11928 4508
rect 12428 4499 12440 4545
rect 12492 4536 12498 4548
rect 18248 4536 18276 4635
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 21821 4675 21879 4681
rect 21821 4641 21833 4675
rect 21867 4672 21879 4675
rect 22186 4672 22192 4684
rect 21867 4644 22192 4672
rect 21867 4641 21879 4644
rect 21821 4635 21879 4641
rect 22186 4632 22192 4644
rect 22244 4632 22250 4684
rect 23106 4632 23112 4684
rect 23164 4672 23170 4684
rect 29546 4672 29552 4684
rect 23164 4644 28212 4672
rect 29507 4644 29552 4672
rect 23164 4632 23170 4644
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4604 18383 4607
rect 19429 4607 19487 4613
rect 18371 4576 19334 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 12492 4508 12528 4536
rect 13556 4508 18276 4536
rect 12434 4496 12440 4499
rect 12492 4496 12498 4508
rect 13556 4477 13584 4508
rect 13541 4471 13599 4477
rect 13541 4468 13553 4471
rect 11900 4440 13553 4468
rect 13541 4437 13553 4440
rect 13587 4437 13599 4471
rect 13541 4431 13599 4437
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 16117 4471 16175 4477
rect 16117 4468 16129 4471
rect 15160 4440 16129 4468
rect 15160 4428 15166 4440
rect 16117 4437 16129 4440
rect 16163 4468 16175 4471
rect 18138 4468 18144 4480
rect 16163 4440 18144 4468
rect 16163 4437 16175 4440
rect 16117 4431 16175 4437
rect 18138 4428 18144 4440
rect 18196 4428 18202 4480
rect 19306 4468 19334 4576
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 20622 4604 20628 4616
rect 19475 4576 20628 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 23198 4564 23204 4616
rect 23256 4564 23262 4616
rect 25501 4607 25559 4613
rect 25501 4604 25513 4607
rect 24688 4576 25513 4604
rect 24688 4545 24716 4576
rect 25501 4573 25513 4576
rect 25547 4573 25559 4607
rect 25501 4567 25559 4573
rect 26050 4564 26056 4616
rect 26108 4604 26114 4616
rect 27433 4607 27491 4613
rect 27433 4604 27445 4607
rect 26108 4576 27445 4604
rect 26108 4564 26114 4576
rect 27433 4573 27445 4576
rect 27479 4604 27491 4607
rect 27479 4576 27936 4604
rect 27479 4573 27491 4576
rect 27433 4567 27491 4573
rect 24673 4539 24731 4545
rect 24673 4505 24685 4539
rect 24719 4505 24731 4539
rect 24673 4499 24731 4505
rect 24889 4539 24947 4545
rect 24889 4505 24901 4539
rect 24935 4536 24947 4539
rect 26068 4536 26096 4564
rect 26602 4536 26608 4548
rect 24935 4508 26096 4536
rect 26563 4508 26608 4536
rect 24935 4505 24947 4508
rect 24889 4499 24947 4505
rect 23569 4471 23627 4477
rect 23569 4468 23581 4471
rect 19306 4440 23581 4468
rect 23569 4437 23581 4440
rect 23615 4468 23627 4471
rect 24688 4468 24716 4499
rect 26602 4496 26608 4508
rect 26660 4496 26666 4548
rect 26821 4539 26879 4545
rect 26821 4505 26833 4539
rect 26867 4536 26879 4539
rect 27614 4536 27620 4548
rect 26867 4508 27384 4536
rect 27575 4508 27620 4536
rect 26867 4505 26879 4508
rect 26821 4499 26879 4505
rect 23615 4440 24716 4468
rect 26973 4471 27031 4477
rect 23615 4437 23627 4440
rect 23569 4431 23627 4437
rect 26973 4437 26985 4471
rect 27019 4468 27031 4471
rect 27246 4468 27252 4480
rect 27019 4440 27252 4468
rect 27019 4437 27031 4440
rect 26973 4431 27031 4437
rect 27246 4428 27252 4440
rect 27304 4428 27310 4480
rect 27356 4468 27384 4508
rect 27614 4496 27620 4508
rect 27672 4496 27678 4548
rect 27801 4471 27859 4477
rect 27801 4468 27813 4471
rect 27356 4440 27813 4468
rect 27801 4437 27813 4440
rect 27847 4437 27859 4471
rect 27908 4468 27936 4576
rect 28184 4536 28212 4644
rect 29546 4632 29552 4644
rect 29604 4632 29610 4684
rect 29656 4672 29684 4712
rect 29656 4644 32076 4672
rect 29454 4604 29460 4616
rect 28460 4576 29460 4604
rect 28460 4545 28488 4576
rect 29454 4564 29460 4576
rect 29512 4564 29518 4616
rect 30926 4564 30932 4616
rect 30984 4564 30990 4616
rect 28445 4539 28503 4545
rect 28445 4536 28457 4539
rect 28184 4508 28457 4536
rect 28445 4505 28457 4508
rect 28491 4505 28503 4539
rect 28445 4499 28503 4505
rect 28661 4539 28719 4545
rect 28661 4505 28673 4539
rect 28707 4536 28719 4539
rect 29822 4536 29828 4548
rect 28707 4508 29684 4536
rect 29783 4508 29828 4536
rect 28707 4505 28719 4508
rect 28661 4499 28719 4505
rect 28813 4471 28871 4477
rect 28813 4468 28825 4471
rect 27908 4440 28825 4468
rect 27801 4431 27859 4437
rect 28813 4437 28825 4440
rect 28859 4468 28871 4471
rect 29178 4468 29184 4480
rect 28859 4440 29184 4468
rect 28859 4437 28871 4440
rect 28813 4431 28871 4437
rect 29178 4428 29184 4440
rect 29236 4428 29242 4480
rect 29656 4468 29684 4508
rect 29822 4496 29828 4508
rect 29880 4496 29886 4548
rect 31772 4545 31800 4644
rect 31757 4539 31815 4545
rect 31757 4505 31769 4539
rect 31803 4505 31815 4539
rect 31757 4499 31815 4505
rect 31938 4496 31944 4548
rect 31996 4545 32002 4548
rect 31996 4539 32015 4545
rect 32003 4505 32015 4539
rect 32048 4536 32076 4644
rect 32232 4604 32260 4712
rect 33686 4700 33692 4712
rect 33744 4700 33750 4752
rect 32232 4576 32904 4604
rect 32585 4539 32643 4545
rect 32585 4536 32597 4539
rect 32048 4508 32597 4536
rect 31996 4499 32015 4505
rect 32585 4505 32597 4508
rect 32631 4505 32643 4539
rect 32585 4499 32643 4505
rect 31996 4496 32002 4499
rect 30006 4468 30012 4480
rect 29656 4440 30012 4468
rect 30006 4428 30012 4440
rect 30064 4428 30070 4480
rect 31386 4428 31392 4480
rect 31444 4468 31450 4480
rect 32785 4471 32843 4477
rect 32785 4468 32797 4471
rect 31444 4440 32797 4468
rect 31444 4428 31450 4440
rect 32785 4437 32797 4440
rect 32831 4437 32843 4471
rect 32876 4468 32904 4576
rect 33318 4564 33324 4616
rect 33376 4604 33382 4616
rect 34790 4604 34796 4616
rect 33376 4576 34796 4604
rect 33376 4564 33382 4576
rect 34790 4564 34796 4576
rect 34848 4564 34854 4616
rect 42794 4564 42800 4616
rect 42852 4604 42858 4616
rect 43901 4607 43959 4613
rect 43901 4604 43913 4607
rect 42852 4576 43913 4604
rect 42852 4564 42858 4576
rect 43901 4573 43913 4576
rect 43947 4573 43959 4607
rect 43901 4567 43959 4573
rect 33410 4536 33416 4548
rect 33371 4508 33416 4536
rect 33410 4496 33416 4508
rect 33468 4496 33474 4548
rect 33594 4496 33600 4548
rect 33652 4545 33658 4548
rect 33652 4539 33671 4545
rect 33659 4505 33671 4539
rect 33652 4499 33671 4505
rect 33652 4496 33658 4499
rect 33502 4468 33508 4480
rect 32876 4440 33508 4468
rect 32785 4431 32843 4437
rect 33502 4428 33508 4440
rect 33560 4428 33566 4480
rect 44082 4468 44088 4480
rect 44043 4440 44088 4468
rect 44082 4428 44088 4440
rect 44140 4428 44146 4480
rect 1104 4378 45056 4400
rect 1104 4326 11898 4378
rect 11950 4326 11962 4378
rect 12014 4326 12026 4378
rect 12078 4326 12090 4378
rect 12142 4326 12154 4378
rect 12206 4326 22846 4378
rect 22898 4326 22910 4378
rect 22962 4326 22974 4378
rect 23026 4326 23038 4378
rect 23090 4326 23102 4378
rect 23154 4326 33794 4378
rect 33846 4326 33858 4378
rect 33910 4326 33922 4378
rect 33974 4326 33986 4378
rect 34038 4326 34050 4378
rect 34102 4326 44742 4378
rect 44794 4326 44806 4378
rect 44858 4326 44870 4378
rect 44922 4326 44934 4378
rect 44986 4326 44998 4378
rect 45050 4326 45056 4378
rect 1104 4304 45056 4326
rect 14737 4267 14795 4273
rect 14737 4233 14749 4267
rect 14783 4264 14795 4267
rect 14826 4264 14832 4276
rect 14783 4236 14832 4264
rect 14783 4233 14795 4236
rect 14737 4227 14795 4233
rect 14826 4224 14832 4236
rect 14884 4224 14890 4276
rect 15102 4264 15108 4276
rect 15063 4236 15108 4264
rect 15102 4224 15108 4236
rect 15160 4224 15166 4276
rect 15194 4224 15200 4276
rect 15252 4264 15258 4276
rect 15252 4236 15297 4264
rect 15252 4224 15258 4236
rect 25314 4224 25320 4276
rect 25372 4264 25378 4276
rect 26142 4264 26148 4276
rect 25372 4236 26148 4264
rect 25372 4224 25378 4236
rect 26142 4224 26148 4236
rect 26200 4224 26206 4276
rect 29086 4224 29092 4276
rect 29144 4264 29150 4276
rect 29917 4267 29975 4273
rect 29917 4264 29929 4267
rect 29144 4236 29929 4264
rect 29144 4224 29150 4236
rect 29917 4233 29929 4236
rect 29963 4264 29975 4267
rect 30558 4264 30564 4276
rect 29963 4236 30564 4264
rect 29963 4233 29975 4236
rect 29917 4227 29975 4233
rect 30558 4224 30564 4236
rect 30616 4224 30622 4276
rect 33410 4264 33416 4276
rect 31864 4236 33416 4264
rect 11790 4156 11796 4208
rect 11848 4196 11854 4208
rect 22278 4196 22284 4208
rect 11848 4168 12020 4196
rect 11848 4156 11854 4168
rect 11606 4088 11612 4140
rect 11664 4128 11670 4140
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11664 4100 11897 4128
rect 11664 4088 11670 4100
rect 11885 4097 11897 4100
rect 11931 4097 11943 4131
rect 11992 4128 12020 4168
rect 17420 4168 19104 4196
rect 12141 4131 12199 4137
rect 12141 4128 12153 4131
rect 11992 4100 12153 4128
rect 11885 4091 11943 4097
rect 12141 4097 12153 4100
rect 12187 4097 12199 4131
rect 12141 4091 12199 4097
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 12768 4100 12940 4128
rect 12768 4088 12774 4100
rect 12912 4060 12940 4100
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 17420 4137 17448 4168
rect 17405 4131 17463 4137
rect 17405 4128 17417 4131
rect 17276 4100 17417 4128
rect 17276 4088 17282 4100
rect 17405 4097 17417 4100
rect 17451 4097 17463 4131
rect 17405 4091 17463 4097
rect 18230 4088 18236 4140
rect 18288 4128 18294 4140
rect 19076 4137 19104 4168
rect 21928 4168 22284 4196
rect 19061 4131 19119 4137
rect 18288 4100 18333 4128
rect 18288 4088 18294 4100
rect 19061 4097 19073 4131
rect 19107 4097 19119 4131
rect 19061 4091 19119 4097
rect 14550 4060 14556 4072
rect 12912 4032 14556 4060
rect 14550 4020 14556 4032
rect 14608 4060 14614 4072
rect 15381 4063 15439 4069
rect 15381 4060 15393 4063
rect 14608 4032 15393 4060
rect 14608 4020 14614 4032
rect 15381 4029 15393 4032
rect 15427 4029 15439 4063
rect 18138 4060 18144 4072
rect 18099 4032 18144 4060
rect 15381 4023 15439 4029
rect 18138 4020 18144 4032
rect 18196 4020 18202 4072
rect 18601 4063 18659 4069
rect 18601 4029 18613 4063
rect 18647 4060 18659 4063
rect 19426 4060 19432 4072
rect 18647 4032 19432 4060
rect 18647 4029 18659 4032
rect 18601 4023 18659 4029
rect 19426 4020 19432 4032
rect 19484 4020 19490 4072
rect 13265 3995 13323 4001
rect 13265 3961 13277 3995
rect 13311 3961 13323 3995
rect 21928 3992 21956 4168
rect 22278 4156 22284 4168
rect 22336 4156 22342 4208
rect 24394 4196 24400 4208
rect 23598 4168 24400 4196
rect 24394 4156 24400 4168
rect 24452 4156 24458 4208
rect 24854 4156 24860 4208
rect 24912 4196 24918 4208
rect 27614 4196 27620 4208
rect 24912 4168 27620 4196
rect 24912 4156 24918 4168
rect 24302 4128 24308 4140
rect 24263 4100 24308 4128
rect 24302 4088 24308 4100
rect 24360 4088 24366 4140
rect 24489 4131 24547 4137
rect 24489 4097 24501 4131
rect 24535 4097 24547 4131
rect 24489 4091 24547 4097
rect 24949 4131 25007 4137
rect 24949 4097 24961 4131
rect 24995 4128 25007 4131
rect 25038 4128 25044 4140
rect 24995 4100 25044 4128
rect 24995 4097 25007 4100
rect 24949 4091 25007 4097
rect 22097 4063 22155 4069
rect 22097 4029 22109 4063
rect 22143 4029 22155 4063
rect 22097 4023 22155 4029
rect 22373 4063 22431 4069
rect 22373 4029 22385 4063
rect 22419 4060 22431 4063
rect 23382 4060 23388 4072
rect 22419 4032 23388 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 13265 3955 13323 3961
rect 15948 3964 21956 3992
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 13280 3924 13308 3955
rect 15948 3924 15976 3964
rect 12584 3896 15976 3924
rect 12584 3884 12590 3896
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 16816 3896 16957 3924
rect 16816 3884 16822 3896
rect 16945 3893 16957 3896
rect 16991 3893 17003 3927
rect 16945 3887 17003 3893
rect 17497 3927 17555 3933
rect 17497 3893 17509 3927
rect 17543 3924 17555 3927
rect 17770 3924 17776 3936
rect 17543 3896 17776 3924
rect 17543 3893 17555 3896
rect 17497 3887 17555 3893
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 19153 3927 19211 3933
rect 19153 3893 19165 3927
rect 19199 3924 19211 3927
rect 19242 3924 19248 3936
rect 19199 3896 19248 3924
rect 19199 3893 19211 3896
rect 19153 3887 19211 3893
rect 19242 3884 19248 3896
rect 19300 3884 19306 3936
rect 22112 3924 22140 4023
rect 23382 4020 23388 4032
rect 23440 4020 23446 4072
rect 24504 3992 24532 4091
rect 25038 4088 25044 4100
rect 25096 4088 25102 4140
rect 25133 4131 25191 4137
rect 25133 4097 25145 4131
rect 25179 4097 25191 4131
rect 26050 4128 26056 4140
rect 26011 4100 26056 4128
rect 25133 4091 25191 4097
rect 24762 4020 24768 4072
rect 24820 4060 24826 4072
rect 25148 4060 25176 4091
rect 26050 4088 26056 4100
rect 26108 4088 26114 4140
rect 26252 4137 26280 4168
rect 27614 4156 27620 4168
rect 27672 4156 27678 4208
rect 28074 4156 28080 4208
rect 28132 4156 28138 4208
rect 31754 4196 31760 4208
rect 30024 4168 31760 4196
rect 30024 4140 30052 4168
rect 31754 4156 31760 4168
rect 31812 4156 31818 4208
rect 26237 4131 26295 4137
rect 26237 4097 26249 4131
rect 26283 4097 26295 4131
rect 26237 4091 26295 4097
rect 26970 4088 26976 4140
rect 27028 4128 27034 4140
rect 27249 4131 27307 4137
rect 27249 4128 27261 4131
rect 27028 4100 27261 4128
rect 27028 4088 27034 4100
rect 27249 4097 27261 4100
rect 27295 4097 27307 4131
rect 27249 4091 27307 4097
rect 29454 4088 29460 4140
rect 29512 4128 29518 4140
rect 29733 4131 29791 4137
rect 29733 4128 29745 4131
rect 29512 4100 29745 4128
rect 29512 4088 29518 4100
rect 29733 4097 29745 4100
rect 29779 4097 29791 4131
rect 29733 4091 29791 4097
rect 30006 4088 30012 4140
rect 30064 4128 30070 4140
rect 31205 4131 31263 4137
rect 30064 4100 30109 4128
rect 30064 4088 30070 4100
rect 31205 4097 31217 4131
rect 31251 4128 31263 4131
rect 31294 4128 31300 4140
rect 31251 4100 31300 4128
rect 31251 4097 31263 4100
rect 31205 4091 31263 4097
rect 31294 4088 31300 4100
rect 31352 4088 31358 4140
rect 31864 4128 31892 4236
rect 33410 4224 33416 4236
rect 33468 4224 33474 4276
rect 32674 4196 32680 4208
rect 32140 4168 32680 4196
rect 32140 4137 32168 4168
rect 32674 4156 32680 4168
rect 32732 4156 32738 4208
rect 32858 4156 32864 4208
rect 32916 4156 32922 4208
rect 31404 4100 31892 4128
rect 32125 4131 32183 4137
rect 27522 4060 27528 4072
rect 24820 4032 25176 4060
rect 27483 4032 27528 4060
rect 24820 4020 24826 4032
rect 27522 4020 27528 4032
rect 27580 4020 27586 4072
rect 27614 4020 27620 4072
rect 27672 4060 27678 4072
rect 28997 4063 29055 4069
rect 28997 4060 29009 4063
rect 27672 4032 29009 4060
rect 27672 4020 27678 4032
rect 28997 4029 29009 4032
rect 29043 4029 29055 4063
rect 28997 4023 29055 4029
rect 29362 4020 29368 4072
rect 29420 4060 29426 4072
rect 31113 4063 31171 4069
rect 31113 4060 31125 4063
rect 29420 4032 31125 4060
rect 29420 4020 29426 4032
rect 31113 4029 31125 4032
rect 31159 4060 31171 4063
rect 31404 4060 31432 4100
rect 32125 4097 32137 4131
rect 32171 4097 32183 4131
rect 32125 4091 32183 4097
rect 32401 4063 32459 4069
rect 32401 4060 32413 4063
rect 31159 4032 31432 4060
rect 31726 4032 32413 4060
rect 31159 4029 31171 4032
rect 31113 4023 31171 4029
rect 25498 3992 25504 4004
rect 23400 3964 24532 3992
rect 24872 3964 25504 3992
rect 22186 3924 22192 3936
rect 22112 3896 22192 3924
rect 22186 3884 22192 3896
rect 22244 3884 22250 3936
rect 22738 3884 22744 3936
rect 22796 3924 22802 3936
rect 23400 3924 23428 3964
rect 23842 3924 23848 3936
rect 22796 3896 23428 3924
rect 23803 3896 23848 3924
rect 22796 3884 22802 3896
rect 23842 3884 23848 3896
rect 23900 3884 23906 3936
rect 24305 3927 24363 3933
rect 24305 3893 24317 3927
rect 24351 3924 24363 3927
rect 24872 3924 24900 3964
rect 25498 3952 25504 3964
rect 25556 3952 25562 4004
rect 31573 3995 31631 4001
rect 31573 3961 31585 3995
rect 31619 3992 31631 3995
rect 31726 3992 31754 4032
rect 32401 4029 32413 4032
rect 32447 4029 32459 4063
rect 32401 4023 32459 4029
rect 31619 3964 31754 3992
rect 31619 3961 31631 3964
rect 31573 3955 31631 3961
rect 25038 3924 25044 3936
rect 24351 3896 24900 3924
rect 24999 3896 25044 3924
rect 24351 3893 24363 3896
rect 24305 3887 24363 3893
rect 25038 3884 25044 3896
rect 25096 3884 25102 3936
rect 29086 3884 29092 3936
rect 29144 3924 29150 3936
rect 29549 3927 29607 3933
rect 29549 3924 29561 3927
rect 29144 3896 29561 3924
rect 29144 3884 29150 3896
rect 29549 3893 29561 3896
rect 29595 3893 29607 3927
rect 29549 3887 29607 3893
rect 31294 3884 31300 3936
rect 31352 3924 31358 3936
rect 33873 3927 33931 3933
rect 33873 3924 33885 3927
rect 31352 3896 33885 3924
rect 31352 3884 31358 3896
rect 33873 3893 33885 3896
rect 33919 3924 33931 3927
rect 43898 3924 43904 3936
rect 33919 3896 43904 3924
rect 33919 3893 33931 3896
rect 33873 3887 33931 3893
rect 43898 3884 43904 3896
rect 43956 3884 43962 3936
rect 1104 3834 44896 3856
rect 1104 3782 6424 3834
rect 6476 3782 6488 3834
rect 6540 3782 6552 3834
rect 6604 3782 6616 3834
rect 6668 3782 6680 3834
rect 6732 3782 17372 3834
rect 17424 3782 17436 3834
rect 17488 3782 17500 3834
rect 17552 3782 17564 3834
rect 17616 3782 17628 3834
rect 17680 3782 28320 3834
rect 28372 3782 28384 3834
rect 28436 3782 28448 3834
rect 28500 3782 28512 3834
rect 28564 3782 28576 3834
rect 28628 3782 39268 3834
rect 39320 3782 39332 3834
rect 39384 3782 39396 3834
rect 39448 3782 39460 3834
rect 39512 3782 39524 3834
rect 39576 3782 44896 3834
rect 1104 3760 44896 3782
rect 11517 3723 11575 3729
rect 11517 3689 11529 3723
rect 11563 3720 11575 3723
rect 12434 3720 12440 3732
rect 11563 3692 12440 3720
rect 11563 3689 11575 3692
rect 11517 3683 11575 3689
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 18230 3680 18236 3732
rect 18288 3720 18294 3732
rect 23566 3720 23572 3732
rect 18288 3692 22094 3720
rect 23527 3692 23572 3720
rect 18288 3680 18294 3692
rect 11422 3612 11428 3664
rect 11480 3652 11486 3664
rect 12161 3655 12219 3661
rect 12161 3652 12173 3655
rect 11480 3624 12173 3652
rect 11480 3612 11486 3624
rect 12161 3621 12173 3624
rect 12207 3621 12219 3655
rect 22066 3652 22094 3692
rect 23566 3680 23572 3692
rect 23624 3680 23630 3732
rect 23750 3720 23756 3732
rect 23711 3692 23756 3720
rect 23750 3680 23756 3692
rect 23808 3680 23814 3732
rect 24394 3680 24400 3732
rect 24452 3720 24458 3732
rect 24489 3723 24547 3729
rect 24489 3720 24501 3723
rect 24452 3692 24501 3720
rect 24452 3680 24458 3692
rect 24489 3689 24501 3692
rect 24535 3689 24547 3723
rect 24489 3683 24547 3689
rect 27249 3723 27307 3729
rect 27249 3689 27261 3723
rect 27295 3720 27307 3723
rect 27522 3720 27528 3732
rect 27295 3692 27528 3720
rect 27295 3689 27307 3692
rect 27249 3683 27307 3689
rect 27522 3680 27528 3692
rect 27580 3680 27586 3732
rect 28074 3720 28080 3732
rect 28035 3692 28080 3720
rect 28074 3680 28080 3692
rect 28132 3680 28138 3732
rect 28813 3723 28871 3729
rect 28813 3689 28825 3723
rect 28859 3720 28871 3723
rect 29549 3723 29607 3729
rect 29549 3720 29561 3723
rect 28859 3692 29561 3720
rect 28859 3689 28871 3692
rect 28813 3683 28871 3689
rect 29549 3689 29561 3692
rect 29595 3689 29607 3723
rect 29549 3683 29607 3689
rect 29822 3680 29828 3732
rect 29880 3720 29886 3732
rect 30285 3723 30343 3729
rect 30285 3720 30297 3723
rect 29880 3692 30297 3720
rect 29880 3680 29886 3692
rect 30285 3689 30297 3692
rect 30331 3689 30343 3723
rect 30285 3683 30343 3689
rect 30926 3680 30932 3732
rect 30984 3720 30990 3732
rect 31021 3723 31079 3729
rect 31021 3720 31033 3723
rect 30984 3692 31033 3720
rect 30984 3680 30990 3692
rect 31021 3689 31033 3692
rect 31067 3689 31079 3723
rect 31021 3683 31079 3689
rect 31849 3723 31907 3729
rect 31849 3689 31861 3723
rect 31895 3720 31907 3723
rect 33226 3720 33232 3732
rect 31895 3692 33232 3720
rect 31895 3689 31907 3692
rect 31849 3683 31907 3689
rect 33226 3680 33232 3692
rect 33284 3680 33290 3732
rect 23842 3652 23848 3664
rect 22066 3624 23848 3652
rect 12161 3615 12219 3621
rect 23842 3612 23848 3624
rect 23900 3652 23906 3664
rect 24762 3652 24768 3664
rect 23900 3624 24768 3652
rect 23900 3612 23906 3624
rect 24762 3612 24768 3624
rect 24820 3612 24826 3664
rect 28997 3655 29055 3661
rect 28997 3621 29009 3655
rect 29043 3652 29055 3655
rect 29043 3624 30328 3652
rect 29043 3621 29055 3624
rect 28997 3615 29055 3621
rect 12618 3584 12624 3596
rect 12579 3556 12624 3584
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 16758 3584 16764 3596
rect 12768 3556 12813 3584
rect 16719 3556 16764 3584
rect 12768 3544 12774 3556
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 19242 3584 19248 3596
rect 19203 3556 19248 3584
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 22094 3544 22100 3596
rect 22152 3584 22158 3596
rect 30300 3584 30328 3624
rect 22152 3556 30052 3584
rect 30300 3556 30420 3584
rect 22152 3544 22158 3556
rect 1578 3516 1584 3528
rect 1539 3488 1584 3516
rect 1578 3476 1584 3488
rect 1636 3476 1642 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11204 3488 11713 3516
rect 11204 3476 11210 3488
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 12526 3516 12532 3528
rect 12487 3488 12532 3516
rect 11701 3479 11759 3485
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 12636 3516 12664 3544
rect 12986 3516 12992 3528
rect 12636 3488 12992 3516
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 15746 3516 15752 3528
rect 15707 3488 15752 3516
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3516 15899 3519
rect 16393 3519 16451 3525
rect 16393 3516 16405 3519
rect 15887 3488 16405 3516
rect 15887 3485 15899 3488
rect 15841 3479 15899 3485
rect 16393 3485 16405 3488
rect 16439 3485 16451 3519
rect 19610 3516 19616 3528
rect 19571 3488 19616 3516
rect 16393 3479 16451 3485
rect 19610 3476 19616 3488
rect 19668 3476 19674 3528
rect 21039 3519 21097 3525
rect 21039 3485 21051 3519
rect 21085 3516 21097 3519
rect 21726 3516 21732 3528
rect 21085 3488 21732 3516
rect 21085 3485 21097 3488
rect 21039 3479 21097 3485
rect 21726 3476 21732 3488
rect 21784 3516 21790 3528
rect 22189 3519 22247 3525
rect 22189 3516 22201 3519
rect 21784 3488 22201 3516
rect 21784 3476 21790 3488
rect 22189 3485 22201 3488
rect 22235 3485 22247 3519
rect 22738 3516 22744 3528
rect 22189 3479 22247 3485
rect 22388 3488 22744 3516
rect 17126 3408 17132 3460
rect 17184 3408 17190 3460
rect 20162 3408 20168 3460
rect 20220 3408 20226 3460
rect 18138 3340 18144 3392
rect 18196 3389 18202 3392
rect 22388 3389 22416 3488
rect 22738 3476 22744 3488
rect 22796 3516 22802 3528
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 22796 3488 24409 3516
rect 22796 3476 22802 3488
rect 24397 3485 24409 3488
rect 24443 3516 24455 3519
rect 24443 3488 26648 3516
rect 24443 3485 24455 3488
rect 24397 3479 24455 3485
rect 23385 3451 23443 3457
rect 23385 3417 23397 3451
rect 23431 3417 23443 3451
rect 23385 3411 23443 3417
rect 23601 3451 23659 3457
rect 23601 3417 23613 3451
rect 23647 3448 23659 3451
rect 25038 3448 25044 3460
rect 23647 3420 25044 3448
rect 23647 3417 23659 3420
rect 23601 3411 23659 3417
rect 18196 3383 18245 3389
rect 18196 3349 18199 3383
rect 18233 3349 18245 3383
rect 18196 3343 18245 3349
rect 22373 3383 22431 3389
rect 22373 3349 22385 3383
rect 22419 3349 22431 3383
rect 23400 3380 23428 3411
rect 25038 3408 25044 3420
rect 25096 3408 25102 3460
rect 26620 3448 26648 3488
rect 27246 3476 27252 3528
rect 27304 3516 27310 3528
rect 27433 3519 27491 3525
rect 27433 3516 27445 3519
rect 27304 3488 27445 3516
rect 27304 3476 27310 3488
rect 27433 3485 27445 3488
rect 27479 3485 27491 3519
rect 27982 3516 27988 3528
rect 27943 3488 27988 3516
rect 27433 3479 27491 3485
rect 27982 3476 27988 3488
rect 28040 3476 28046 3528
rect 29086 3516 29092 3528
rect 28920 3488 29092 3516
rect 28000 3448 28028 3476
rect 26620 3420 28028 3448
rect 28629 3451 28687 3457
rect 28629 3417 28641 3451
rect 28675 3417 28687 3451
rect 28629 3411 28687 3417
rect 28834 3451 28892 3457
rect 28834 3417 28846 3451
rect 28880 3448 28892 3451
rect 28920 3448 28948 3488
rect 29086 3476 29092 3488
rect 29144 3476 29150 3528
rect 29178 3476 29184 3528
rect 29236 3516 29242 3528
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 29236 3488 29561 3516
rect 29236 3476 29242 3488
rect 29549 3485 29561 3488
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 28880 3420 28948 3448
rect 28880 3417 28892 3420
rect 28834 3411 28892 3417
rect 26602 3380 26608 3392
rect 23400 3352 26608 3380
rect 22373 3343 22431 3349
rect 18196 3340 18202 3343
rect 26602 3340 26608 3352
rect 26660 3380 26666 3392
rect 28644 3380 28672 3411
rect 29362 3380 29368 3392
rect 26660 3352 29368 3380
rect 26660 3340 26666 3352
rect 29362 3340 29368 3352
rect 29420 3340 29426 3392
rect 30024 3380 30052 3556
rect 30392 3512 30420 3556
rect 30558 3544 30564 3596
rect 30616 3584 30622 3596
rect 30616 3556 31984 3584
rect 30616 3544 30622 3556
rect 30461 3515 30519 3521
rect 30926 3516 30932 3528
rect 30461 3512 30473 3515
rect 30392 3484 30473 3512
rect 30461 3481 30473 3484
rect 30507 3481 30519 3515
rect 30887 3488 30932 3516
rect 30461 3475 30519 3481
rect 30926 3476 30932 3488
rect 30984 3476 30990 3528
rect 31754 3476 31760 3528
rect 31812 3516 31818 3528
rect 31956 3525 31984 3556
rect 31941 3519 31999 3525
rect 31812 3488 31857 3516
rect 31812 3476 31818 3488
rect 31941 3485 31953 3519
rect 31987 3516 31999 3519
rect 32582 3516 32588 3528
rect 31987 3488 32588 3516
rect 31987 3485 31999 3488
rect 31941 3479 31999 3485
rect 32582 3476 32588 3488
rect 32640 3476 32646 3528
rect 44174 3516 44180 3528
rect 44135 3488 44180 3516
rect 44174 3476 44180 3488
rect 44232 3476 44238 3528
rect 33502 3380 33508 3392
rect 30024 3352 33508 3380
rect 33502 3340 33508 3352
rect 33560 3340 33566 3392
rect 1104 3290 45056 3312
rect 1104 3238 11898 3290
rect 11950 3238 11962 3290
rect 12014 3238 12026 3290
rect 12078 3238 12090 3290
rect 12142 3238 12154 3290
rect 12206 3238 22846 3290
rect 22898 3238 22910 3290
rect 22962 3238 22974 3290
rect 23026 3238 23038 3290
rect 23090 3238 23102 3290
rect 23154 3238 33794 3290
rect 33846 3238 33858 3290
rect 33910 3238 33922 3290
rect 33974 3238 33986 3290
rect 34038 3238 34050 3290
rect 34102 3238 44742 3290
rect 44794 3238 44806 3290
rect 44858 3238 44870 3290
rect 44922 3238 44934 3290
rect 44986 3238 44998 3290
rect 45050 3238 45056 3290
rect 1104 3216 45056 3238
rect 16025 3179 16083 3185
rect 16025 3145 16037 3179
rect 16071 3176 16083 3179
rect 17126 3176 17132 3188
rect 16071 3148 17132 3176
rect 16071 3145 16083 3148
rect 16025 3139 16083 3145
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 19610 3185 19616 3188
rect 17221 3179 17279 3185
rect 17221 3145 17233 3179
rect 17267 3176 17279 3179
rect 19567 3179 19616 3185
rect 17267 3148 18460 3176
rect 17267 3145 17279 3148
rect 17221 3139 17279 3145
rect 18432 3108 18460 3148
rect 19567 3145 19579 3179
rect 19613 3145 19616 3179
rect 19567 3139 19616 3145
rect 19610 3136 19616 3139
rect 19668 3136 19674 3188
rect 20162 3176 20168 3188
rect 20123 3148 20168 3176
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 23017 3179 23075 3185
rect 23017 3145 23029 3179
rect 23063 3176 23075 3179
rect 23198 3176 23204 3188
rect 23063 3148 23204 3176
rect 23063 3145 23075 3148
rect 23017 3139 23075 3145
rect 23198 3136 23204 3148
rect 23256 3136 23262 3188
rect 23382 3136 23388 3188
rect 23440 3176 23446 3188
rect 23569 3179 23627 3185
rect 23569 3176 23581 3179
rect 23440 3148 23581 3176
rect 23440 3136 23446 3148
rect 23569 3145 23581 3148
rect 23615 3145 23627 3179
rect 23569 3139 23627 3145
rect 31389 3179 31447 3185
rect 31389 3145 31401 3179
rect 31435 3176 31447 3179
rect 32858 3176 32864 3188
rect 31435 3148 32864 3176
rect 31435 3145 31447 3148
rect 31389 3139 31447 3145
rect 32858 3136 32864 3148
rect 32916 3136 32922 3188
rect 34057 3179 34115 3185
rect 34057 3145 34069 3179
rect 34103 3176 34115 3179
rect 34146 3176 34152 3188
rect 34103 3148 34152 3176
rect 34103 3145 34115 3148
rect 34057 3139 34115 3145
rect 34146 3136 34152 3148
rect 34204 3136 34210 3188
rect 43254 3176 43260 3188
rect 43215 3148 43260 3176
rect 43254 3136 43260 3148
rect 43312 3136 43318 3188
rect 43438 3136 43444 3188
rect 43496 3176 43502 3188
rect 43901 3179 43959 3185
rect 43901 3176 43913 3179
rect 43496 3148 43913 3176
rect 43496 3136 43502 3148
rect 43901 3145 43913 3148
rect 43947 3145 43959 3179
rect 43901 3139 43959 3145
rect 18432 3080 18538 3108
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6822 3040 6828 3052
rect 6595 3012 6828 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 12897 3043 12955 3049
rect 12897 3040 12909 3043
rect 11296 3012 12909 3040
rect 11296 3000 11302 3012
rect 12897 3009 12909 3012
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 17129 3043 17187 3049
rect 17129 3040 17141 3043
rect 15979 3012 17141 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 17129 3009 17141 3012
rect 17175 3009 17187 3043
rect 17770 3040 17776 3052
rect 17731 3012 17776 3040
rect 17129 3003 17187 3009
rect 17144 2972 17172 3003
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 18138 3040 18144 3052
rect 18099 3012 18144 3040
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 20073 3043 20131 3049
rect 20073 3009 20085 3043
rect 20119 3009 20131 3043
rect 20073 3003 20131 3009
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3040 22155 3043
rect 22462 3040 22468 3052
rect 22143 3012 22468 3040
rect 22143 3009 22155 3012
rect 22097 3003 22155 3009
rect 20088 2972 20116 3003
rect 22462 3000 22468 3012
rect 22520 3000 22526 3052
rect 22738 3000 22744 3052
rect 22796 3040 22802 3052
rect 22925 3043 22983 3049
rect 22925 3040 22937 3043
rect 22796 3012 22937 3040
rect 22796 3000 22802 3012
rect 22925 3009 22937 3012
rect 22971 3009 22983 3043
rect 23750 3040 23756 3052
rect 23711 3012 23756 3040
rect 22925 3003 22983 3009
rect 23750 3000 23756 3012
rect 23808 3000 23814 3052
rect 27982 3000 27988 3052
rect 28040 3040 28046 3052
rect 30926 3040 30932 3052
rect 28040 3012 30932 3040
rect 28040 3000 28046 3012
rect 30926 3000 30932 3012
rect 30984 3040 30990 3052
rect 31297 3043 31355 3049
rect 31297 3040 31309 3043
rect 30984 3012 31309 3040
rect 30984 3000 30990 3012
rect 31297 3009 31309 3012
rect 31343 3009 31355 3043
rect 34164 3040 34192 3136
rect 34517 3043 34575 3049
rect 34517 3040 34529 3043
rect 34164 3012 34529 3040
rect 31297 3003 31355 3009
rect 34517 3009 34529 3012
rect 34563 3009 34575 3043
rect 34517 3003 34575 3009
rect 43441 3043 43499 3049
rect 43441 3009 43453 3043
rect 43487 3009 43499 3043
rect 43441 3003 43499 3009
rect 17144 2944 20116 2972
rect 43456 2972 43484 3003
rect 43806 3000 43812 3052
rect 43864 3040 43870 3052
rect 44085 3043 44143 3049
rect 44085 3040 44097 3043
rect 43864 3012 44097 3040
rect 43864 3000 43870 3012
rect 44085 3009 44097 3012
rect 44131 3009 44143 3043
rect 44085 3003 44143 3009
rect 45094 2972 45100 2984
rect 43456 2944 45100 2972
rect 17788 2916 17816 2944
rect 45094 2932 45100 2944
rect 45152 2932 45158 2984
rect 17770 2864 17776 2916
rect 17828 2864 17834 2916
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 6270 2796 6276 2848
rect 6328 2836 6334 2848
rect 6365 2839 6423 2845
rect 6365 2836 6377 2839
rect 6328 2808 6377 2836
rect 6328 2796 6334 2808
rect 6365 2805 6377 2808
rect 6411 2805 6423 2839
rect 6365 2799 6423 2805
rect 13081 2839 13139 2845
rect 13081 2805 13093 2839
rect 13127 2836 13139 2839
rect 14458 2836 14464 2848
rect 13127 2808 14464 2836
rect 13127 2805 13139 2808
rect 13081 2799 13139 2805
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 21913 2839 21971 2845
rect 21913 2805 21925 2839
rect 21959 2836 21971 2839
rect 22646 2836 22652 2848
rect 21959 2808 22652 2836
rect 21959 2805 21971 2808
rect 21913 2799 21971 2805
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 34333 2839 34391 2845
rect 34333 2805 34345 2839
rect 34379 2836 34391 2839
rect 35526 2836 35532 2848
rect 34379 2808 35532 2836
rect 34379 2805 34391 2808
rect 34333 2799 34391 2805
rect 35526 2796 35532 2808
rect 35584 2796 35590 2848
rect 1104 2746 44896 2768
rect 1104 2694 6424 2746
rect 6476 2694 6488 2746
rect 6540 2694 6552 2746
rect 6604 2694 6616 2746
rect 6668 2694 6680 2746
rect 6732 2694 17372 2746
rect 17424 2694 17436 2746
rect 17488 2694 17500 2746
rect 17552 2694 17564 2746
rect 17616 2694 17628 2746
rect 17680 2694 28320 2746
rect 28372 2694 28384 2746
rect 28436 2694 28448 2746
rect 28500 2694 28512 2746
rect 28564 2694 28576 2746
rect 28628 2694 39268 2746
rect 39320 2694 39332 2746
rect 39384 2694 39396 2746
rect 39448 2694 39460 2746
rect 39512 2694 39524 2746
rect 39576 2694 44896 2746
rect 1104 2672 44896 2694
rect 12986 2632 12992 2644
rect 12947 2604 12992 2632
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 25869 2635 25927 2641
rect 25869 2601 25881 2635
rect 25915 2632 25927 2635
rect 35986 2632 35992 2644
rect 25915 2604 35992 2632
rect 25915 2601 25927 2604
rect 25869 2595 25927 2601
rect 35986 2592 35992 2604
rect 36044 2592 36050 2644
rect 37277 2635 37335 2641
rect 37277 2601 37289 2635
rect 37323 2632 37335 2635
rect 37366 2632 37372 2644
rect 37323 2604 37372 2632
rect 37323 2601 37335 2604
rect 37277 2595 37335 2601
rect 37366 2592 37372 2604
rect 37424 2592 37430 2644
rect 15102 2524 15108 2576
rect 15160 2564 15166 2576
rect 43073 2567 43131 2573
rect 43073 2564 43085 2567
rect 15160 2536 43085 2564
rect 15160 2524 15166 2536
rect 43073 2533 43085 2536
rect 43119 2533 43131 2567
rect 43073 2527 43131 2533
rect 14 2456 20 2508
rect 72 2496 78 2508
rect 2225 2499 2283 2505
rect 2225 2496 2237 2499
rect 72 2468 2237 2496
rect 72 2456 78 2468
rect 2225 2465 2237 2468
rect 2271 2465 2283 2499
rect 17770 2496 17776 2508
rect 17731 2468 17776 2496
rect 2225 2459 2283 2465
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1360 2400 1593 2428
rect 1360 2388 1366 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3292 2400 3985 2428
rect 3292 2388 3298 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4580 2400 4813 2428
rect 4580 2388 4586 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 6270 2388 6276 2440
rect 6328 2428 6334 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6328 2400 6561 2428
rect 6328 2388 6334 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7800 2400 8033 2428
rect 7800 2388 7806 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 8021 2391 8079 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11020 2400 11713 2428
rect 11020 2388 11026 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 12952 2400 13185 2428
rect 12952 2388 12958 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 14458 2428 14464 2440
rect 14419 2400 14464 2428
rect 13173 2391 13231 2397
rect 14458 2388 14464 2400
rect 14516 2388 14522 2440
rect 15473 2431 15531 2437
rect 15473 2397 15485 2431
rect 15519 2428 15531 2431
rect 16114 2428 16120 2440
rect 15519 2400 16120 2428
rect 15519 2397 15531 2400
rect 15473 2391 15531 2397
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17460 2400 17509 2428
rect 17460 2388 17466 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20680 2400 20913 2428
rect 20680 2388 20686 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 22646 2428 22652 2440
rect 22607 2400 22652 2428
rect 20901 2391 20959 2397
rect 22646 2388 22652 2400
rect 22704 2388 22710 2440
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23900 2400 24593 2428
rect 23900 2388 23906 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 25832 2400 26065 2428
rect 25832 2388 25838 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 26053 2391 26111 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 27120 2400 27169 2428
rect 27120 2388 27126 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29052 2400 29745 2428
rect 29052 2388 29058 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30282 2388 30288 2440
rect 30340 2428 30346 2440
rect 30561 2431 30619 2437
rect 30561 2428 30573 2431
rect 30340 2400 30573 2428
rect 30340 2388 30346 2400
rect 30561 2397 30573 2400
rect 30607 2397 30619 2431
rect 35526 2428 35532 2440
rect 35487 2400 35532 2428
rect 30561 2391 30619 2397
rect 35526 2388 35532 2400
rect 35584 2388 35590 2440
rect 36722 2388 36728 2440
rect 36780 2428 36786 2440
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 36780 2400 37473 2428
rect 36780 2388 36786 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 38654 2388 38660 2440
rect 38712 2428 38718 2440
rect 38933 2431 38991 2437
rect 38933 2428 38945 2431
rect 38712 2400 38945 2428
rect 38712 2388 38718 2400
rect 38933 2397 38945 2400
rect 38979 2397 38991 2431
rect 38933 2391 38991 2397
rect 39942 2388 39948 2440
rect 40000 2428 40006 2440
rect 40221 2431 40279 2437
rect 40221 2428 40233 2431
rect 40000 2400 40233 2428
rect 40000 2388 40006 2400
rect 40221 2397 40233 2400
rect 40267 2397 40279 2431
rect 43898 2428 43904 2440
rect 43859 2400 43904 2428
rect 40221 2391 40279 2397
rect 43898 2388 43904 2400
rect 43956 2388 43962 2440
rect 19702 2320 19708 2372
rect 19760 2360 19766 2372
rect 19760 2332 31248 2360
rect 19760 2320 19766 2332
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9953 2295 10011 2301
rect 9953 2292 9965 2295
rect 9732 2264 9965 2292
rect 9732 2252 9738 2264
rect 9953 2261 9965 2264
rect 9999 2261 10011 2295
rect 9953 2255 10011 2261
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 14240 2264 14289 2292
rect 14240 2252 14246 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22833 2295 22891 2301
rect 22833 2292 22845 2295
rect 22612 2264 22845 2292
rect 22612 2252 22618 2264
rect 22833 2261 22845 2264
rect 22879 2261 22891 2295
rect 22833 2255 22891 2261
rect 27341 2295 27399 2301
rect 27341 2261 27353 2295
rect 27387 2292 27399 2295
rect 27430 2292 27436 2304
rect 27387 2264 27436 2292
rect 27387 2261 27399 2264
rect 27341 2255 27399 2261
rect 27430 2252 27436 2264
rect 27488 2252 27494 2304
rect 31220 2292 31248 2332
rect 32214 2320 32220 2372
rect 32272 2360 32278 2372
rect 32585 2363 32643 2369
rect 32585 2360 32597 2363
rect 32272 2332 32597 2360
rect 32272 2320 32278 2332
rect 32585 2329 32597 2332
rect 32631 2329 32643 2363
rect 32585 2323 32643 2329
rect 41874 2320 41880 2372
rect 41932 2360 41938 2372
rect 42889 2363 42947 2369
rect 42889 2360 42901 2363
rect 41932 2332 42901 2360
rect 41932 2320 41938 2332
rect 42889 2329 42901 2332
rect 42935 2329 42947 2363
rect 42889 2323 42947 2329
rect 32306 2292 32312 2304
rect 31220 2264 32312 2292
rect 32306 2252 32312 2264
rect 32364 2292 32370 2304
rect 32677 2295 32735 2301
rect 32677 2292 32689 2295
rect 32364 2264 32689 2292
rect 32364 2252 32370 2264
rect 32677 2261 32689 2264
rect 32723 2261 32735 2295
rect 32677 2255 32735 2261
rect 35434 2252 35440 2304
rect 35492 2292 35498 2304
rect 35713 2295 35771 2301
rect 35713 2292 35725 2295
rect 35492 2264 35725 2292
rect 35492 2252 35498 2264
rect 35713 2261 35725 2264
rect 35759 2261 35771 2295
rect 44082 2292 44088 2304
rect 44043 2264 44088 2292
rect 35713 2255 35771 2261
rect 44082 2252 44088 2264
rect 44140 2252 44146 2304
rect 1104 2202 45056 2224
rect 1104 2150 11898 2202
rect 11950 2150 11962 2202
rect 12014 2150 12026 2202
rect 12078 2150 12090 2202
rect 12142 2150 12154 2202
rect 12206 2150 22846 2202
rect 22898 2150 22910 2202
rect 22962 2150 22974 2202
rect 23026 2150 23038 2202
rect 23090 2150 23102 2202
rect 23154 2150 33794 2202
rect 33846 2150 33858 2202
rect 33910 2150 33922 2202
rect 33974 2150 33986 2202
rect 34038 2150 34050 2202
rect 34102 2150 44742 2202
rect 44794 2150 44806 2202
rect 44858 2150 44870 2202
rect 44922 2150 44934 2202
rect 44986 2150 44998 2202
rect 45050 2150 45056 2202
rect 1104 2128 45056 2150
<< via1 >>
rect 11898 17382 11950 17434
rect 11962 17382 12014 17434
rect 12026 17382 12078 17434
rect 12090 17382 12142 17434
rect 12154 17382 12206 17434
rect 22846 17382 22898 17434
rect 22910 17382 22962 17434
rect 22974 17382 23026 17434
rect 23038 17382 23090 17434
rect 23102 17382 23154 17434
rect 33794 17382 33846 17434
rect 33858 17382 33910 17434
rect 33922 17382 33974 17434
rect 33986 17382 34038 17434
rect 34050 17382 34102 17434
rect 44742 17382 44794 17434
rect 44806 17382 44858 17434
rect 44870 17382 44922 17434
rect 44934 17382 44986 17434
rect 44998 17382 45050 17434
rect 17408 17280 17460 17332
rect 20720 17280 20772 17332
rect 37280 17280 37332 17332
rect 40592 17280 40644 17332
rect 44088 17323 44140 17332
rect 44088 17289 44097 17323
rect 44097 17289 44131 17323
rect 44131 17289 44140 17323
rect 44088 17280 44140 17289
rect 1308 17212 1360 17264
rect 3240 17212 3292 17264
rect 38660 17212 38712 17264
rect 2228 17187 2280 17196
rect 2228 17153 2237 17187
rect 2237 17153 2271 17187
rect 2271 17153 2280 17187
rect 2228 17144 2280 17153
rect 4528 17144 4580 17196
rect 6460 17144 6512 17196
rect 7748 17144 7800 17196
rect 9680 17144 9732 17196
rect 11060 17144 11112 17196
rect 12900 17144 12952 17196
rect 14188 17144 14240 17196
rect 16120 17144 16172 17196
rect 16764 17144 16816 17196
rect 19340 17144 19392 17196
rect 4896 17119 4948 17128
rect 4160 17051 4212 17060
rect 4160 17017 4169 17051
rect 4169 17017 4203 17051
rect 4203 17017 4212 17051
rect 4160 17008 4212 17017
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 17224 17076 17276 17128
rect 17960 17076 18012 17128
rect 22560 17144 22612 17196
rect 23848 17144 23900 17196
rect 25780 17144 25832 17196
rect 27712 17144 27764 17196
rect 29000 17144 29052 17196
rect 30932 17144 30984 17196
rect 32220 17144 32272 17196
rect 34152 17144 34204 17196
rect 35440 17144 35492 17196
rect 37372 17144 37424 17196
rect 40684 17187 40736 17196
rect 40684 17153 40693 17187
rect 40693 17153 40727 17187
rect 40727 17153 40736 17187
rect 40684 17144 40736 17153
rect 41880 17144 41932 17196
rect 43904 17187 43956 17196
rect 43904 17153 43913 17187
rect 43913 17153 43947 17187
rect 43947 17153 43956 17187
rect 43904 17144 43956 17153
rect 32588 17119 32640 17128
rect 32588 17085 32597 17119
rect 32597 17085 32631 17119
rect 32631 17085 32640 17119
rect 32588 17076 32640 17085
rect 45100 17076 45152 17128
rect 42524 17008 42576 17060
rect 3056 16983 3108 16992
rect 3056 16949 3065 16983
rect 3065 16949 3099 16983
rect 3099 16949 3108 16983
rect 3056 16940 3108 16949
rect 9680 16940 9732 16992
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 23572 16940 23624 16992
rect 34152 16940 34204 16992
rect 38936 16983 38988 16992
rect 38936 16949 38945 16983
rect 38945 16949 38979 16983
rect 38979 16949 38988 16983
rect 38936 16940 38988 16949
rect 6424 16838 6476 16890
rect 6488 16838 6540 16890
rect 6552 16838 6604 16890
rect 6616 16838 6668 16890
rect 6680 16838 6732 16890
rect 17372 16838 17424 16890
rect 17436 16838 17488 16890
rect 17500 16838 17552 16890
rect 17564 16838 17616 16890
rect 17628 16838 17680 16890
rect 28320 16838 28372 16890
rect 28384 16838 28436 16890
rect 28448 16838 28500 16890
rect 28512 16838 28564 16890
rect 28576 16838 28628 16890
rect 39268 16838 39320 16890
rect 39332 16838 39384 16890
rect 39396 16838 39448 16890
rect 39460 16838 39512 16890
rect 39524 16838 39576 16890
rect 3976 16779 4028 16788
rect 3976 16745 3985 16779
rect 3985 16745 4019 16779
rect 4019 16745 4028 16779
rect 3976 16736 4028 16745
rect 4896 16736 4948 16788
rect 11704 16736 11756 16788
rect 16856 16736 16908 16788
rect 33692 16736 33744 16788
rect 43444 16779 43496 16788
rect 43444 16745 43453 16779
rect 43453 16745 43487 16779
rect 43487 16745 43496 16779
rect 43444 16736 43496 16745
rect 43812 16736 43864 16788
rect 10692 16668 10744 16720
rect 20 16532 72 16584
rect 15660 16532 15712 16584
rect 17132 16575 17184 16584
rect 17132 16541 17141 16575
rect 17141 16541 17175 16575
rect 17175 16541 17184 16575
rect 17132 16532 17184 16541
rect 40040 16575 40092 16584
rect 40040 16541 40049 16575
rect 40049 16541 40083 16575
rect 40083 16541 40092 16575
rect 40040 16532 40092 16541
rect 16764 16396 16816 16448
rect 17960 16396 18012 16448
rect 40684 16396 40736 16448
rect 11898 16294 11950 16346
rect 11962 16294 12014 16346
rect 12026 16294 12078 16346
rect 12090 16294 12142 16346
rect 12154 16294 12206 16346
rect 22846 16294 22898 16346
rect 22910 16294 22962 16346
rect 22974 16294 23026 16346
rect 23038 16294 23090 16346
rect 23102 16294 23154 16346
rect 33794 16294 33846 16346
rect 33858 16294 33910 16346
rect 33922 16294 33974 16346
rect 33986 16294 34038 16346
rect 34050 16294 34102 16346
rect 44742 16294 44794 16346
rect 44806 16294 44858 16346
rect 44870 16294 44922 16346
rect 44934 16294 44986 16346
rect 44998 16294 45050 16346
rect 44180 15895 44232 15904
rect 44180 15861 44189 15895
rect 44189 15861 44223 15895
rect 44223 15861 44232 15895
rect 44180 15852 44232 15861
rect 6424 15750 6476 15802
rect 6488 15750 6540 15802
rect 6552 15750 6604 15802
rect 6616 15750 6668 15802
rect 6680 15750 6732 15802
rect 17372 15750 17424 15802
rect 17436 15750 17488 15802
rect 17500 15750 17552 15802
rect 17564 15750 17616 15802
rect 17628 15750 17680 15802
rect 28320 15750 28372 15802
rect 28384 15750 28436 15802
rect 28448 15750 28500 15802
rect 28512 15750 28564 15802
rect 28576 15750 28628 15802
rect 39268 15750 39320 15802
rect 39332 15750 39384 15802
rect 39396 15750 39448 15802
rect 39460 15750 39512 15802
rect 39524 15750 39576 15802
rect 3148 15444 3200 15496
rect 18604 15444 18656 15496
rect 19156 15444 19208 15496
rect 34888 15487 34940 15496
rect 34888 15453 34897 15487
rect 34897 15453 34931 15487
rect 34931 15453 34940 15487
rect 34888 15444 34940 15453
rect 19248 15419 19300 15428
rect 19248 15385 19257 15419
rect 19257 15385 19291 15419
rect 19291 15385 19300 15419
rect 19248 15376 19300 15385
rect 19432 15419 19484 15428
rect 19432 15385 19441 15419
rect 19441 15385 19475 15419
rect 19475 15385 19484 15419
rect 19432 15376 19484 15385
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 18052 15308 18104 15360
rect 19156 15308 19208 15360
rect 19524 15351 19576 15360
rect 19524 15317 19533 15351
rect 19533 15317 19567 15351
rect 19567 15317 19576 15351
rect 19524 15308 19576 15317
rect 43904 15308 43956 15360
rect 11898 15206 11950 15258
rect 11962 15206 12014 15258
rect 12026 15206 12078 15258
rect 12090 15206 12142 15258
rect 12154 15206 12206 15258
rect 22846 15206 22898 15258
rect 22910 15206 22962 15258
rect 22974 15206 23026 15258
rect 23038 15206 23090 15258
rect 23102 15206 23154 15258
rect 33794 15206 33846 15258
rect 33858 15206 33910 15258
rect 33922 15206 33974 15258
rect 33986 15206 34038 15258
rect 34050 15206 34102 15258
rect 44742 15206 44794 15258
rect 44806 15206 44858 15258
rect 44870 15206 44922 15258
rect 44934 15206 44986 15258
rect 44998 15206 45050 15258
rect 8760 14832 8812 14884
rect 12256 14968 12308 15020
rect 9588 14900 9640 14952
rect 12900 15011 12952 15020
rect 12900 14977 12909 15011
rect 12909 14977 12943 15011
rect 12943 14977 12952 15011
rect 13084 15011 13136 15020
rect 12900 14968 12952 14977
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 18696 15104 18748 15156
rect 19156 15104 19208 15156
rect 18052 15079 18104 15088
rect 18052 15045 18061 15079
rect 18061 15045 18095 15079
rect 18095 15045 18104 15079
rect 18052 15036 18104 15045
rect 19248 15036 19300 15088
rect 16120 14968 16172 15020
rect 18788 14968 18840 15020
rect 19800 14968 19852 15020
rect 19432 14900 19484 14952
rect 9128 14832 9180 14884
rect 8944 14807 8996 14816
rect 8944 14773 8953 14807
rect 8953 14773 8987 14807
rect 8987 14773 8996 14807
rect 8944 14764 8996 14773
rect 11796 14764 11848 14816
rect 13268 14764 13320 14816
rect 13544 14807 13596 14816
rect 13544 14773 13553 14807
rect 13553 14773 13587 14807
rect 13587 14773 13596 14807
rect 13544 14764 13596 14773
rect 15752 14764 15804 14816
rect 18420 14764 18472 14816
rect 18604 14832 18656 14884
rect 23296 14900 23348 14952
rect 23388 14832 23440 14884
rect 19340 14764 19392 14816
rect 20536 14764 20588 14816
rect 6424 14662 6476 14714
rect 6488 14662 6540 14714
rect 6552 14662 6604 14714
rect 6616 14662 6668 14714
rect 6680 14662 6732 14714
rect 17372 14662 17424 14714
rect 17436 14662 17488 14714
rect 17500 14662 17552 14714
rect 17564 14662 17616 14714
rect 17628 14662 17680 14714
rect 28320 14662 28372 14714
rect 28384 14662 28436 14714
rect 28448 14662 28500 14714
rect 28512 14662 28564 14714
rect 28576 14662 28628 14714
rect 39268 14662 39320 14714
rect 39332 14662 39384 14714
rect 39396 14662 39448 14714
rect 39460 14662 39512 14714
rect 39524 14662 39576 14714
rect 8392 14560 8444 14612
rect 19524 14560 19576 14612
rect 9220 14492 9272 14544
rect 9496 14424 9548 14476
rect 19156 14492 19208 14544
rect 9772 14356 9824 14408
rect 12532 14424 12584 14476
rect 12716 14424 12768 14476
rect 12900 14356 12952 14408
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 19800 14467 19852 14476
rect 19800 14433 19809 14467
rect 19809 14433 19843 14467
rect 19843 14433 19852 14467
rect 23940 14560 23992 14612
rect 19800 14424 19852 14433
rect 13268 14399 13320 14408
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 13268 14356 13320 14365
rect 8760 14288 8812 14340
rect 9128 14331 9180 14340
rect 9128 14297 9153 14331
rect 9153 14297 9180 14331
rect 9128 14288 9180 14297
rect 12624 14288 12676 14340
rect 13544 14356 13596 14408
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 16672 14356 16724 14408
rect 19248 14356 19300 14408
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 20168 14356 20220 14408
rect 15568 14288 15620 14340
rect 15752 14331 15804 14340
rect 15752 14297 15786 14331
rect 15786 14297 15804 14331
rect 15752 14288 15804 14297
rect 17592 14331 17644 14340
rect 17592 14297 17626 14331
rect 17626 14297 17644 14331
rect 17592 14288 17644 14297
rect 19800 14288 19852 14340
rect 20536 14331 20588 14340
rect 20536 14297 20561 14331
rect 20561 14297 20588 14331
rect 24676 14356 24728 14408
rect 42984 14399 43036 14408
rect 42984 14365 42993 14399
rect 42993 14365 43027 14399
rect 43027 14365 43036 14399
rect 42984 14356 43036 14365
rect 20536 14288 20588 14297
rect 7380 14263 7432 14272
rect 7380 14229 7389 14263
rect 7389 14229 7423 14263
rect 7423 14229 7432 14263
rect 7380 14220 7432 14229
rect 8024 14263 8076 14272
rect 8024 14229 8033 14263
rect 8033 14229 8067 14263
rect 8067 14229 8076 14263
rect 8024 14220 8076 14229
rect 8576 14220 8628 14272
rect 12348 14263 12400 14272
rect 12348 14229 12357 14263
rect 12357 14229 12391 14263
rect 12391 14229 12400 14263
rect 12348 14220 12400 14229
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 16856 14263 16908 14272
rect 16856 14229 16865 14263
rect 16865 14229 16899 14263
rect 16899 14229 16908 14263
rect 16856 14220 16908 14229
rect 18604 14220 18656 14272
rect 18788 14220 18840 14272
rect 19984 14220 20036 14272
rect 21272 14220 21324 14272
rect 21364 14220 21416 14272
rect 23848 14220 23900 14272
rect 44088 14263 44140 14272
rect 44088 14229 44097 14263
rect 44097 14229 44131 14263
rect 44131 14229 44140 14263
rect 44088 14220 44140 14229
rect 11898 14118 11950 14170
rect 11962 14118 12014 14170
rect 12026 14118 12078 14170
rect 12090 14118 12142 14170
rect 12154 14118 12206 14170
rect 22846 14118 22898 14170
rect 22910 14118 22962 14170
rect 22974 14118 23026 14170
rect 23038 14118 23090 14170
rect 23102 14118 23154 14170
rect 33794 14118 33846 14170
rect 33858 14118 33910 14170
rect 33922 14118 33974 14170
rect 33986 14118 34038 14170
rect 34050 14118 34102 14170
rect 44742 14118 44794 14170
rect 44806 14118 44858 14170
rect 44870 14118 44922 14170
rect 44934 14118 44986 14170
rect 44998 14118 45050 14170
rect 3148 14059 3200 14068
rect 3148 14025 3157 14059
rect 3157 14025 3191 14059
rect 3191 14025 3200 14059
rect 3148 14016 3200 14025
rect 8392 14016 8444 14068
rect 12256 14059 12308 14068
rect 3332 13923 3384 13932
rect 3332 13889 3341 13923
rect 3341 13889 3375 13923
rect 3375 13889 3384 13923
rect 3332 13880 3384 13889
rect 4436 13948 4488 14000
rect 7380 13948 7432 14000
rect 9588 13991 9640 14000
rect 9588 13957 9597 13991
rect 9597 13957 9631 13991
rect 9631 13957 9640 13991
rect 9588 13948 9640 13957
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 12716 14016 12768 14068
rect 12992 14016 13044 14068
rect 13084 14016 13136 14068
rect 15016 14016 15068 14068
rect 16120 14059 16172 14068
rect 16120 14025 16129 14059
rect 16129 14025 16163 14059
rect 16163 14025 16172 14059
rect 16120 14016 16172 14025
rect 17592 14059 17644 14068
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 7104 13812 7156 13864
rect 8944 13880 8996 13932
rect 12624 13880 12676 13932
rect 15476 13948 15528 14000
rect 15568 13948 15620 14000
rect 19800 14016 19852 14068
rect 20168 14059 20220 14068
rect 20168 14025 20177 14059
rect 20177 14025 20211 14059
rect 20211 14025 20220 14059
rect 20168 14016 20220 14025
rect 23388 14059 23440 14068
rect 12808 13880 12860 13932
rect 18512 13948 18564 14000
rect 18696 13948 18748 14000
rect 21364 13948 21416 14000
rect 23388 14025 23397 14059
rect 23397 14025 23431 14059
rect 23431 14025 23440 14059
rect 23388 14016 23440 14025
rect 34888 14016 34940 14068
rect 9680 13812 9732 13864
rect 9220 13787 9272 13796
rect 3056 13676 3108 13728
rect 5356 13719 5408 13728
rect 5356 13685 5365 13719
rect 5365 13685 5399 13719
rect 5399 13685 5408 13719
rect 5356 13676 5408 13685
rect 9220 13753 9229 13787
rect 9229 13753 9263 13787
rect 9263 13753 9272 13787
rect 9220 13744 9272 13753
rect 8668 13676 8720 13728
rect 8760 13719 8812 13728
rect 8760 13685 8769 13719
rect 8769 13685 8803 13719
rect 8803 13685 8812 13719
rect 11152 13744 11204 13796
rect 16856 13880 16908 13932
rect 18604 13880 18656 13932
rect 19340 13880 19392 13932
rect 21272 13923 21324 13932
rect 21272 13889 21281 13923
rect 21281 13889 21315 13923
rect 21315 13889 21324 13923
rect 21272 13880 21324 13889
rect 23388 13880 23440 13932
rect 16304 13812 16356 13864
rect 20628 13812 20680 13864
rect 23204 13812 23256 13864
rect 23940 13855 23992 13864
rect 23940 13821 23949 13855
rect 23949 13821 23983 13855
rect 23983 13821 23992 13855
rect 23940 13812 23992 13821
rect 33692 13991 33744 14000
rect 33692 13957 33701 13991
rect 33701 13957 33735 13991
rect 33735 13957 33744 13991
rect 33692 13948 33744 13957
rect 42984 13948 43036 14000
rect 24216 13880 24268 13932
rect 33232 13880 33284 13932
rect 8760 13676 8812 13685
rect 9772 13719 9824 13728
rect 9772 13685 9781 13719
rect 9781 13685 9815 13719
rect 9815 13685 9824 13719
rect 9772 13676 9824 13685
rect 12348 13676 12400 13728
rect 16396 13744 16448 13796
rect 16856 13676 16908 13728
rect 18420 13719 18472 13728
rect 18420 13685 18429 13719
rect 18429 13685 18463 13719
rect 18463 13685 18472 13719
rect 18420 13676 18472 13685
rect 18604 13719 18656 13728
rect 18604 13685 18613 13719
rect 18613 13685 18647 13719
rect 18647 13685 18656 13719
rect 18604 13676 18656 13685
rect 19984 13719 20036 13728
rect 19984 13685 19993 13719
rect 19993 13685 20027 13719
rect 20027 13685 20036 13719
rect 19984 13676 20036 13685
rect 23480 13676 23532 13728
rect 25412 13744 25464 13796
rect 33232 13676 33284 13728
rect 34520 13812 34572 13864
rect 33692 13744 33744 13796
rect 38936 13676 38988 13728
rect 6424 13574 6476 13626
rect 6488 13574 6540 13626
rect 6552 13574 6604 13626
rect 6616 13574 6668 13626
rect 6680 13574 6732 13626
rect 17372 13574 17424 13626
rect 17436 13574 17488 13626
rect 17500 13574 17552 13626
rect 17564 13574 17616 13626
rect 17628 13574 17680 13626
rect 28320 13574 28372 13626
rect 28384 13574 28436 13626
rect 28448 13574 28500 13626
rect 28512 13574 28564 13626
rect 28576 13574 28628 13626
rect 39268 13574 39320 13626
rect 39332 13574 39384 13626
rect 39396 13574 39448 13626
rect 39460 13574 39512 13626
rect 39524 13574 39576 13626
rect 8392 13515 8444 13524
rect 8392 13481 8401 13515
rect 8401 13481 8435 13515
rect 8435 13481 8444 13515
rect 8392 13472 8444 13481
rect 9036 13472 9088 13524
rect 9496 13515 9548 13524
rect 9496 13481 9505 13515
rect 9505 13481 9539 13515
rect 9539 13481 9548 13515
rect 9496 13472 9548 13481
rect 8944 13447 8996 13456
rect 8944 13413 8953 13447
rect 8953 13413 8987 13447
rect 8987 13413 8996 13447
rect 8944 13404 8996 13413
rect 8668 13336 8720 13388
rect 12992 13404 13044 13456
rect 16028 13404 16080 13456
rect 14464 13336 14516 13388
rect 18512 13404 18564 13456
rect 19432 13404 19484 13456
rect 20260 13404 20312 13456
rect 20996 13404 21048 13456
rect 18788 13336 18840 13388
rect 4436 13268 4488 13320
rect 7104 13268 7156 13320
rect 8852 13268 8904 13320
rect 11152 13311 11204 13320
rect 11152 13277 11161 13311
rect 11161 13277 11195 13311
rect 11195 13277 11204 13311
rect 11152 13268 11204 13277
rect 8024 13200 8076 13252
rect 9588 13200 9640 13252
rect 10784 13200 10836 13252
rect 11888 13268 11940 13320
rect 12532 13268 12584 13320
rect 15292 13268 15344 13320
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 16304 13311 16356 13320
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 17868 13268 17920 13320
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 11520 13132 11572 13184
rect 12900 13132 12952 13184
rect 16212 13243 16264 13252
rect 16212 13209 16221 13243
rect 16221 13209 16255 13243
rect 16255 13209 16264 13243
rect 16212 13200 16264 13209
rect 18420 13200 18472 13252
rect 19156 13268 19208 13320
rect 20628 13336 20680 13388
rect 22744 13404 22796 13456
rect 25412 13404 25464 13456
rect 22192 13336 22244 13388
rect 22284 13336 22336 13388
rect 21364 13268 21416 13320
rect 23296 13268 23348 13320
rect 24216 13268 24268 13320
rect 19340 13200 19392 13252
rect 15016 13175 15068 13184
rect 15016 13141 15025 13175
rect 15025 13141 15059 13175
rect 15059 13141 15068 13175
rect 15016 13132 15068 13141
rect 16488 13175 16540 13184
rect 16488 13141 16497 13175
rect 16497 13141 16531 13175
rect 16531 13141 16540 13175
rect 16488 13132 16540 13141
rect 22744 13200 22796 13252
rect 32588 13336 32640 13388
rect 37280 13379 37332 13388
rect 26332 13311 26384 13320
rect 26332 13277 26341 13311
rect 26341 13277 26375 13311
rect 26375 13277 26384 13311
rect 26332 13268 26384 13277
rect 26792 13311 26844 13320
rect 26792 13277 26801 13311
rect 26801 13277 26835 13311
rect 26835 13277 26844 13311
rect 26792 13268 26844 13277
rect 30288 13311 30340 13320
rect 30288 13277 30297 13311
rect 30297 13277 30331 13311
rect 30331 13277 30340 13311
rect 30288 13268 30340 13277
rect 32312 13268 32364 13320
rect 37280 13345 37289 13379
rect 37289 13345 37323 13379
rect 37323 13345 37332 13379
rect 37280 13336 37332 13345
rect 38936 13336 38988 13388
rect 33324 13268 33376 13320
rect 37648 13268 37700 13320
rect 38292 13311 38344 13320
rect 38292 13277 38301 13311
rect 38301 13277 38335 13311
rect 38335 13277 38344 13311
rect 38292 13268 38344 13277
rect 38384 13311 38436 13320
rect 38384 13277 38393 13311
rect 38393 13277 38427 13311
rect 38427 13277 38436 13311
rect 40960 13404 41012 13456
rect 42616 13404 42668 13456
rect 38384 13268 38436 13277
rect 39672 13268 39724 13320
rect 22376 13132 22428 13184
rect 22652 13132 22704 13184
rect 23296 13132 23348 13184
rect 27804 13200 27856 13252
rect 33232 13200 33284 13252
rect 38476 13200 38528 13252
rect 41972 13200 42024 13252
rect 28724 13132 28776 13184
rect 30472 13132 30524 13184
rect 35624 13132 35676 13184
rect 38568 13175 38620 13184
rect 38568 13141 38577 13175
rect 38577 13141 38611 13175
rect 38611 13141 38620 13175
rect 38568 13132 38620 13141
rect 40224 13132 40276 13184
rect 40500 13175 40552 13184
rect 40500 13141 40509 13175
rect 40509 13141 40543 13175
rect 40543 13141 40552 13175
rect 40500 13132 40552 13141
rect 11898 13030 11950 13082
rect 11962 13030 12014 13082
rect 12026 13030 12078 13082
rect 12090 13030 12142 13082
rect 12154 13030 12206 13082
rect 22846 13030 22898 13082
rect 22910 13030 22962 13082
rect 22974 13030 23026 13082
rect 23038 13030 23090 13082
rect 23102 13030 23154 13082
rect 33794 13030 33846 13082
rect 33858 13030 33910 13082
rect 33922 13030 33974 13082
rect 33986 13030 34038 13082
rect 34050 13030 34102 13082
rect 44742 13030 44794 13082
rect 44806 13030 44858 13082
rect 44870 13030 44922 13082
rect 44934 13030 44986 13082
rect 44998 13030 45050 13082
rect 22284 12971 22336 12980
rect 5356 12860 5408 12912
rect 8576 12860 8628 12912
rect 9036 12903 9088 12912
rect 9036 12869 9045 12903
rect 9045 12869 9079 12903
rect 9079 12869 9088 12903
rect 9036 12860 9088 12869
rect 4436 12835 4488 12844
rect 4436 12801 4445 12835
rect 4445 12801 4479 12835
rect 4479 12801 4488 12835
rect 4436 12792 4488 12801
rect 8760 12792 8812 12844
rect 10508 12792 10560 12844
rect 8392 12724 8444 12776
rect 12532 12860 12584 12912
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 13912 12792 13964 12844
rect 14464 12835 14516 12844
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 14648 12835 14700 12844
rect 14648 12801 14657 12835
rect 14657 12801 14691 12835
rect 14691 12801 14700 12835
rect 14648 12792 14700 12801
rect 15292 12860 15344 12912
rect 15936 12860 15988 12912
rect 17776 12860 17828 12912
rect 22284 12937 22293 12971
rect 22293 12937 22327 12971
rect 22327 12937 22336 12971
rect 22284 12928 22336 12937
rect 22376 12971 22428 12980
rect 22376 12937 22385 12971
rect 22385 12937 22419 12971
rect 22419 12937 22428 12971
rect 23296 12971 23348 12980
rect 22376 12928 22428 12937
rect 23296 12937 23305 12971
rect 23305 12937 23339 12971
rect 23339 12937 23348 12971
rect 23296 12928 23348 12937
rect 23848 12971 23900 12980
rect 23848 12937 23857 12971
rect 23857 12937 23891 12971
rect 23891 12937 23900 12971
rect 23848 12928 23900 12937
rect 24032 12971 24084 12980
rect 24032 12937 24041 12971
rect 24041 12937 24075 12971
rect 24075 12937 24084 12971
rect 24032 12928 24084 12937
rect 16212 12792 16264 12844
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 17868 12792 17920 12844
rect 15292 12724 15344 12776
rect 16304 12724 16356 12776
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 2780 12588 2832 12640
rect 6000 12588 6052 12640
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 12164 12588 12216 12640
rect 13360 12588 13412 12640
rect 15844 12588 15896 12640
rect 20260 12767 20312 12776
rect 20260 12733 20269 12767
rect 20269 12733 20303 12767
rect 20303 12733 20312 12767
rect 20260 12724 20312 12733
rect 25136 12860 25188 12912
rect 20996 12767 21048 12776
rect 20996 12733 21005 12767
rect 21005 12733 21039 12767
rect 21039 12733 21048 12767
rect 20996 12724 21048 12733
rect 21088 12767 21140 12776
rect 21088 12733 21097 12767
rect 21097 12733 21131 12767
rect 21131 12733 21140 12767
rect 21088 12724 21140 12733
rect 22100 12724 22152 12776
rect 21364 12656 21416 12708
rect 23388 12835 23440 12844
rect 22468 12767 22520 12776
rect 22468 12733 22477 12767
rect 22477 12733 22511 12767
rect 22511 12733 22520 12767
rect 23388 12801 23397 12835
rect 23397 12801 23431 12835
rect 23431 12801 23440 12835
rect 23388 12792 23440 12801
rect 22468 12724 22520 12733
rect 23480 12724 23532 12776
rect 23020 12656 23072 12708
rect 23388 12656 23440 12708
rect 24216 12792 24268 12844
rect 27988 12860 28040 12912
rect 30472 12860 30524 12912
rect 35624 12971 35676 12980
rect 35624 12937 35633 12971
rect 35633 12937 35667 12971
rect 35667 12937 35676 12971
rect 35624 12928 35676 12937
rect 38384 12928 38436 12980
rect 39120 12928 39172 12980
rect 30748 12792 30800 12844
rect 25320 12724 25372 12776
rect 24584 12656 24636 12708
rect 27252 12767 27304 12776
rect 20904 12588 20956 12640
rect 22284 12588 22336 12640
rect 25044 12588 25096 12640
rect 26700 12656 26752 12708
rect 26516 12588 26568 12640
rect 26792 12588 26844 12640
rect 27252 12733 27261 12767
rect 27261 12733 27295 12767
rect 27295 12733 27304 12767
rect 27252 12724 27304 12733
rect 29460 12767 29512 12776
rect 29460 12733 29469 12767
rect 29469 12733 29503 12767
rect 29503 12733 29512 12767
rect 29460 12724 29512 12733
rect 30196 12724 30248 12776
rect 29092 12588 29144 12640
rect 34520 12860 34572 12912
rect 34336 12835 34388 12844
rect 34336 12801 34345 12835
rect 34345 12801 34379 12835
rect 34379 12801 34388 12835
rect 34336 12792 34388 12801
rect 34520 12767 34572 12776
rect 34520 12733 34529 12767
rect 34529 12733 34563 12767
rect 34563 12733 34572 12767
rect 34520 12724 34572 12733
rect 37004 12724 37056 12776
rect 37556 12835 37608 12844
rect 37556 12801 37590 12835
rect 37590 12801 37608 12835
rect 39764 12860 39816 12912
rect 37556 12792 37608 12801
rect 40592 12792 40644 12844
rect 42708 12792 42760 12844
rect 30196 12588 30248 12640
rect 30472 12588 30524 12640
rect 33600 12588 33652 12640
rect 40040 12724 40092 12776
rect 38568 12656 38620 12708
rect 39672 12588 39724 12640
rect 41972 12588 42024 12640
rect 44088 12588 44140 12640
rect 6424 12486 6476 12538
rect 6488 12486 6540 12538
rect 6552 12486 6604 12538
rect 6616 12486 6668 12538
rect 6680 12486 6732 12538
rect 17372 12486 17424 12538
rect 17436 12486 17488 12538
rect 17500 12486 17552 12538
rect 17564 12486 17616 12538
rect 17628 12486 17680 12538
rect 28320 12486 28372 12538
rect 28384 12486 28436 12538
rect 28448 12486 28500 12538
rect 28512 12486 28564 12538
rect 28576 12486 28628 12538
rect 39268 12486 39320 12538
rect 39332 12486 39384 12538
rect 39396 12486 39448 12538
rect 39460 12486 39512 12538
rect 39524 12486 39576 12538
rect 5448 12384 5500 12436
rect 12072 12384 12124 12436
rect 12256 12384 12308 12436
rect 8208 12316 8260 12368
rect 4436 12248 4488 12300
rect 9588 12248 9640 12300
rect 12348 12316 12400 12368
rect 12532 12291 12584 12300
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 13728 12316 13780 12368
rect 14648 12384 14700 12436
rect 15476 12384 15528 12436
rect 12532 12248 12584 12257
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 2688 12180 2740 12232
rect 6828 12180 6880 12232
rect 8852 12180 8904 12232
rect 8944 12180 8996 12232
rect 10784 12223 10836 12232
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 13084 12180 13136 12232
rect 13544 12180 13596 12232
rect 6552 12112 6604 12164
rect 10324 12112 10376 12164
rect 11520 12112 11572 12164
rect 13912 12180 13964 12232
rect 16488 12316 16540 12368
rect 17776 12316 17828 12368
rect 16028 12291 16080 12300
rect 16028 12257 16037 12291
rect 16037 12257 16071 12291
rect 16071 12257 16080 12291
rect 16028 12248 16080 12257
rect 20444 12316 20496 12368
rect 22100 12384 22152 12436
rect 23204 12384 23256 12436
rect 24216 12384 24268 12436
rect 24584 12427 24636 12436
rect 24584 12393 24593 12427
rect 24593 12393 24627 12427
rect 24627 12393 24636 12427
rect 24584 12384 24636 12393
rect 25228 12427 25280 12436
rect 25228 12393 25237 12427
rect 25237 12393 25271 12427
rect 25271 12393 25280 12427
rect 25228 12384 25280 12393
rect 25320 12384 25372 12436
rect 26332 12384 26384 12436
rect 27804 12427 27856 12436
rect 27804 12393 27813 12427
rect 27813 12393 27847 12427
rect 27847 12393 27856 12427
rect 27804 12384 27856 12393
rect 29092 12384 29144 12436
rect 29460 12384 29512 12436
rect 29920 12384 29972 12436
rect 30472 12384 30524 12436
rect 30564 12384 30616 12436
rect 33140 12384 33192 12436
rect 34336 12384 34388 12436
rect 22560 12316 22612 12368
rect 24676 12316 24728 12368
rect 26240 12316 26292 12368
rect 20352 12248 20404 12300
rect 20904 12291 20956 12300
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 15844 12180 15896 12232
rect 16764 12180 16816 12232
rect 16856 12223 16908 12232
rect 16856 12189 16865 12223
rect 16865 12189 16899 12223
rect 16899 12189 16908 12223
rect 17868 12223 17920 12232
rect 16856 12180 16908 12189
rect 17868 12189 17877 12223
rect 17877 12189 17911 12223
rect 17911 12189 17920 12223
rect 17868 12180 17920 12189
rect 18420 12180 18472 12232
rect 19156 12180 19208 12232
rect 20628 12180 20680 12232
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 22468 12248 22520 12300
rect 25228 12248 25280 12300
rect 26516 12248 26568 12300
rect 27436 12248 27488 12300
rect 23020 12180 23072 12232
rect 23388 12180 23440 12232
rect 2964 12044 3016 12096
rect 3884 12044 3936 12096
rect 7196 12087 7248 12096
rect 7196 12053 7205 12087
rect 7205 12053 7239 12087
rect 7239 12053 7248 12087
rect 7196 12044 7248 12053
rect 9220 12044 9272 12096
rect 9404 12087 9456 12096
rect 9404 12053 9413 12087
rect 9413 12053 9447 12087
rect 9447 12053 9456 12087
rect 9404 12044 9456 12053
rect 9864 12087 9916 12096
rect 9864 12053 9873 12087
rect 9873 12053 9907 12087
rect 9907 12053 9916 12087
rect 9864 12044 9916 12053
rect 10232 12044 10284 12096
rect 12348 12044 12400 12096
rect 12624 12044 12676 12096
rect 17224 12044 17276 12096
rect 17592 12044 17644 12096
rect 17960 12087 18012 12096
rect 17960 12053 17969 12087
rect 17969 12053 18003 12087
rect 18003 12053 18012 12087
rect 17960 12044 18012 12053
rect 18052 12044 18104 12096
rect 19800 12044 19852 12096
rect 21272 12112 21324 12164
rect 24032 12180 24084 12232
rect 24492 12112 24544 12164
rect 26424 12112 26476 12164
rect 27620 12180 27672 12232
rect 30748 12316 30800 12368
rect 31300 12248 31352 12300
rect 34244 12248 34296 12300
rect 37740 12384 37792 12436
rect 38016 12316 38068 12368
rect 39856 12316 39908 12368
rect 36544 12291 36596 12300
rect 36544 12257 36553 12291
rect 36553 12257 36587 12291
rect 36587 12257 36596 12291
rect 40500 12384 40552 12436
rect 42708 12384 42760 12436
rect 40408 12316 40460 12368
rect 36544 12248 36596 12257
rect 29092 12180 29144 12232
rect 30012 12223 30064 12232
rect 30012 12189 30021 12223
rect 30021 12189 30055 12223
rect 30055 12189 30064 12223
rect 30012 12180 30064 12189
rect 30288 12180 30340 12232
rect 33324 12180 33376 12232
rect 34152 12180 34204 12232
rect 37004 12223 37056 12232
rect 23480 12044 23532 12096
rect 24216 12044 24268 12096
rect 24768 12087 24820 12096
rect 24768 12053 24777 12087
rect 24777 12053 24811 12087
rect 24811 12053 24820 12087
rect 24768 12044 24820 12053
rect 25044 12044 25096 12096
rect 28632 12044 28684 12096
rect 29920 12087 29972 12096
rect 29920 12053 29929 12087
rect 29929 12053 29963 12087
rect 29963 12053 29972 12087
rect 29920 12044 29972 12053
rect 30196 12112 30248 12164
rect 30380 12112 30432 12164
rect 30656 12112 30708 12164
rect 33508 12112 33560 12164
rect 30748 12044 30800 12096
rect 31208 12044 31260 12096
rect 37004 12189 37013 12223
rect 37013 12189 37047 12223
rect 37047 12189 37056 12223
rect 37004 12180 37056 12189
rect 39028 12223 39080 12232
rect 39028 12189 39037 12223
rect 39037 12189 39071 12223
rect 39071 12189 39080 12223
rect 39028 12180 39080 12189
rect 40592 12248 40644 12300
rect 42616 12248 42668 12300
rect 39304 12223 39356 12232
rect 39304 12189 39313 12223
rect 39313 12189 39347 12223
rect 39347 12189 39356 12223
rect 39304 12180 39356 12189
rect 39672 12180 39724 12232
rect 37188 12044 37240 12096
rect 39856 12112 39908 12164
rect 40316 12112 40368 12164
rect 40776 12112 40828 12164
rect 41052 12112 41104 12164
rect 38292 12044 38344 12096
rect 39304 12044 39356 12096
rect 42432 12087 42484 12096
rect 42432 12053 42441 12087
rect 42441 12053 42475 12087
rect 42475 12053 42484 12087
rect 42432 12044 42484 12053
rect 11898 11942 11950 11994
rect 11962 11942 12014 11994
rect 12026 11942 12078 11994
rect 12090 11942 12142 11994
rect 12154 11942 12206 11994
rect 22846 11942 22898 11994
rect 22910 11942 22962 11994
rect 22974 11942 23026 11994
rect 23038 11942 23090 11994
rect 23102 11942 23154 11994
rect 33794 11942 33846 11994
rect 33858 11942 33910 11994
rect 33922 11942 33974 11994
rect 33986 11942 34038 11994
rect 34050 11942 34102 11994
rect 44742 11942 44794 11994
rect 44806 11942 44858 11994
rect 44870 11942 44922 11994
rect 44934 11942 44986 11994
rect 44998 11942 45050 11994
rect 2596 11840 2648 11892
rect 4620 11840 4672 11892
rect 5448 11883 5500 11892
rect 3700 11772 3752 11824
rect 5448 11849 5457 11883
rect 5457 11849 5491 11883
rect 5491 11849 5500 11883
rect 5448 11840 5500 11849
rect 7196 11840 7248 11892
rect 9864 11840 9916 11892
rect 17040 11883 17092 11892
rect 17040 11849 17049 11883
rect 17049 11849 17083 11883
rect 17083 11849 17092 11883
rect 17040 11840 17092 11849
rect 19156 11840 19208 11892
rect 19708 11840 19760 11892
rect 21088 11840 21140 11892
rect 21272 11840 21324 11892
rect 22744 11840 22796 11892
rect 9220 11815 9272 11824
rect 9220 11781 9229 11815
rect 9229 11781 9263 11815
rect 9263 11781 9272 11815
rect 9220 11772 9272 11781
rect 10600 11772 10652 11824
rect 12532 11772 12584 11824
rect 4252 11636 4304 11688
rect 4068 11568 4120 11620
rect 6092 11568 6144 11620
rect 6552 11611 6604 11620
rect 6552 11577 6561 11611
rect 6561 11577 6595 11611
rect 6595 11577 6604 11611
rect 6552 11568 6604 11577
rect 11704 11704 11756 11756
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 12164 11704 12216 11756
rect 18236 11772 18288 11824
rect 18604 11772 18656 11824
rect 8484 11636 8536 11688
rect 8944 11679 8996 11688
rect 8944 11645 8953 11679
rect 8953 11645 8987 11679
rect 8987 11645 8996 11679
rect 8944 11636 8996 11645
rect 10232 11636 10284 11688
rect 10508 11636 10560 11688
rect 7288 11500 7340 11552
rect 8024 11543 8076 11552
rect 8024 11509 8033 11543
rect 8033 11509 8067 11543
rect 8067 11509 8076 11543
rect 8024 11500 8076 11509
rect 8392 11500 8444 11552
rect 11704 11568 11756 11620
rect 12348 11636 12400 11688
rect 13452 11568 13504 11620
rect 15936 11704 15988 11756
rect 17224 11747 17276 11756
rect 17224 11713 17233 11747
rect 17233 11713 17267 11747
rect 17267 11713 17276 11747
rect 17224 11704 17276 11713
rect 15476 11679 15528 11688
rect 15200 11568 15252 11620
rect 15476 11645 15485 11679
rect 15485 11645 15519 11679
rect 15519 11645 15528 11679
rect 15476 11636 15528 11645
rect 15752 11636 15804 11688
rect 16672 11636 16724 11688
rect 17868 11679 17920 11688
rect 17868 11645 17877 11679
rect 17877 11645 17911 11679
rect 17911 11645 17920 11679
rect 17868 11636 17920 11645
rect 18144 11679 18196 11688
rect 18144 11645 18153 11679
rect 18153 11645 18187 11679
rect 18187 11645 18196 11679
rect 18144 11636 18196 11645
rect 18236 11636 18288 11688
rect 20352 11747 20404 11756
rect 20352 11713 20361 11747
rect 20361 11713 20395 11747
rect 20395 11713 20404 11747
rect 20352 11704 20404 11713
rect 20076 11636 20128 11688
rect 20996 11636 21048 11688
rect 22008 11704 22060 11756
rect 23480 11704 23532 11756
rect 23940 11772 23992 11824
rect 24216 11772 24268 11824
rect 26332 11840 26384 11892
rect 26792 11840 26844 11892
rect 27252 11840 27304 11892
rect 27988 11840 28040 11892
rect 28632 11840 28684 11892
rect 29920 11883 29972 11892
rect 29460 11772 29512 11824
rect 29920 11849 29929 11883
rect 29929 11849 29963 11883
rect 29963 11849 29972 11883
rect 29920 11840 29972 11849
rect 30656 11883 30708 11892
rect 30656 11849 30665 11883
rect 30665 11849 30699 11883
rect 30699 11849 30708 11883
rect 30656 11840 30708 11849
rect 33232 11883 33284 11892
rect 33232 11849 33241 11883
rect 33241 11849 33275 11883
rect 33275 11849 33284 11883
rect 33232 11840 33284 11849
rect 33508 11840 33560 11892
rect 34704 11883 34756 11892
rect 34704 11849 34713 11883
rect 34713 11849 34747 11883
rect 34747 11849 34756 11883
rect 34704 11840 34756 11849
rect 37556 11840 37608 11892
rect 39028 11840 39080 11892
rect 39948 11840 40000 11892
rect 41604 11840 41656 11892
rect 24492 11704 24544 11756
rect 24676 11747 24728 11756
rect 24676 11713 24685 11747
rect 24685 11713 24719 11747
rect 24719 11713 24728 11747
rect 24676 11704 24728 11713
rect 23940 11636 23992 11688
rect 12072 11500 12124 11552
rect 12716 11500 12768 11552
rect 14096 11500 14148 11552
rect 16672 11500 16724 11552
rect 26148 11636 26200 11688
rect 26424 11679 26476 11688
rect 26424 11645 26433 11679
rect 26433 11645 26467 11679
rect 26467 11645 26476 11679
rect 26424 11636 26476 11645
rect 26700 11704 26752 11756
rect 27252 11704 27304 11756
rect 27620 11747 27672 11756
rect 27620 11713 27629 11747
rect 27629 11713 27663 11747
rect 27663 11713 27672 11747
rect 27620 11704 27672 11713
rect 28816 11704 28868 11756
rect 20076 11500 20128 11552
rect 22008 11543 22060 11552
rect 22008 11509 22017 11543
rect 22017 11509 22051 11543
rect 22051 11509 22060 11543
rect 22008 11500 22060 11509
rect 23296 11543 23348 11552
rect 23296 11509 23305 11543
rect 23305 11509 23339 11543
rect 23339 11509 23348 11543
rect 23296 11500 23348 11509
rect 23480 11500 23532 11552
rect 24584 11500 24636 11552
rect 25964 11568 26016 11620
rect 27344 11568 27396 11620
rect 29736 11747 29788 11756
rect 29736 11713 29745 11747
rect 29745 11713 29779 11747
rect 29779 11713 29788 11747
rect 29736 11704 29788 11713
rect 30840 11679 30892 11688
rect 30840 11645 30849 11679
rect 30849 11645 30883 11679
rect 30883 11645 30892 11679
rect 30840 11636 30892 11645
rect 31208 11679 31260 11688
rect 30656 11568 30708 11620
rect 31208 11645 31217 11679
rect 31217 11645 31251 11679
rect 31251 11645 31260 11679
rect 31208 11636 31260 11645
rect 31300 11679 31352 11688
rect 31300 11645 31309 11679
rect 31309 11645 31343 11679
rect 31343 11645 31352 11679
rect 33232 11704 33284 11756
rect 33416 11747 33468 11756
rect 33416 11713 33425 11747
rect 33425 11713 33459 11747
rect 33459 11713 33468 11747
rect 33416 11704 33468 11713
rect 31300 11636 31352 11645
rect 32772 11636 32824 11688
rect 33140 11636 33192 11688
rect 34152 11704 34204 11756
rect 34612 11747 34664 11756
rect 34612 11713 34621 11747
rect 34621 11713 34655 11747
rect 34655 11713 34664 11747
rect 34612 11704 34664 11713
rect 36544 11747 36596 11756
rect 36544 11713 36553 11747
rect 36553 11713 36587 11747
rect 36587 11713 36596 11747
rect 36544 11704 36596 11713
rect 37648 11772 37700 11824
rect 37740 11747 37792 11756
rect 37740 11713 37749 11747
rect 37749 11713 37783 11747
rect 37783 11713 37792 11747
rect 37740 11704 37792 11713
rect 38292 11704 38344 11756
rect 38568 11772 38620 11824
rect 39304 11815 39356 11824
rect 39304 11781 39313 11815
rect 39313 11781 39347 11815
rect 39347 11781 39356 11815
rect 39304 11772 39356 11781
rect 40132 11772 40184 11824
rect 40500 11772 40552 11824
rect 41512 11772 41564 11824
rect 38476 11747 38528 11756
rect 38476 11713 38485 11747
rect 38485 11713 38519 11747
rect 38519 11713 38528 11747
rect 38936 11747 38988 11756
rect 38476 11704 38528 11713
rect 38936 11713 38945 11747
rect 38945 11713 38979 11747
rect 38979 11713 38988 11747
rect 38936 11704 38988 11713
rect 39028 11747 39080 11756
rect 39028 11713 39038 11747
rect 39038 11713 39072 11747
rect 39072 11713 39080 11747
rect 39028 11704 39080 11713
rect 38016 11636 38068 11688
rect 38108 11636 38160 11688
rect 39764 11704 39816 11756
rect 39948 11704 40000 11756
rect 40408 11747 40460 11756
rect 40408 11713 40417 11747
rect 40417 11713 40451 11747
rect 40451 11713 40460 11747
rect 40408 11704 40460 11713
rect 40592 11747 40644 11756
rect 40592 11713 40601 11747
rect 40601 11713 40635 11747
rect 40635 11713 40644 11747
rect 40592 11704 40644 11713
rect 40776 11704 40828 11756
rect 41972 11704 42024 11756
rect 42432 11679 42484 11688
rect 31944 11500 31996 11552
rect 37280 11500 37332 11552
rect 37556 11500 37608 11552
rect 38476 11500 38528 11552
rect 39028 11500 39080 11552
rect 40316 11568 40368 11620
rect 40500 11500 40552 11552
rect 42432 11645 42441 11679
rect 42441 11645 42475 11679
rect 42475 11645 42484 11679
rect 42432 11636 42484 11645
rect 42708 11679 42760 11688
rect 42708 11645 42717 11679
rect 42717 11645 42751 11679
rect 42751 11645 42760 11679
rect 42708 11636 42760 11645
rect 41328 11500 41380 11552
rect 6424 11398 6476 11450
rect 6488 11398 6540 11450
rect 6552 11398 6604 11450
rect 6616 11398 6668 11450
rect 6680 11398 6732 11450
rect 17372 11398 17424 11450
rect 17436 11398 17488 11450
rect 17500 11398 17552 11450
rect 17564 11398 17616 11450
rect 17628 11398 17680 11450
rect 28320 11398 28372 11450
rect 28384 11398 28436 11450
rect 28448 11398 28500 11450
rect 28512 11398 28564 11450
rect 28576 11398 28628 11450
rect 39268 11398 39320 11450
rect 39332 11398 39384 11450
rect 39396 11398 39448 11450
rect 39460 11398 39512 11450
rect 39524 11398 39576 11450
rect 2688 11296 2740 11348
rect 4160 11296 4212 11348
rect 8208 11339 8260 11348
rect 2964 11203 3016 11212
rect 2964 11169 2973 11203
rect 2973 11169 3007 11203
rect 3007 11169 3016 11203
rect 2964 11160 3016 11169
rect 4252 11160 4304 11212
rect 8208 11305 8217 11339
rect 8217 11305 8251 11339
rect 8251 11305 8260 11339
rect 8208 11296 8260 11305
rect 8852 11296 8904 11348
rect 10324 11339 10376 11348
rect 8484 11228 8536 11280
rect 10324 11305 10333 11339
rect 10333 11305 10367 11339
rect 10367 11305 10376 11339
rect 10324 11296 10376 11305
rect 10416 11296 10468 11348
rect 12624 11296 12676 11348
rect 12992 11296 13044 11348
rect 15936 11339 15988 11348
rect 12164 11228 12216 11280
rect 12440 11228 12492 11280
rect 15936 11305 15945 11339
rect 15945 11305 15979 11339
rect 15979 11305 15988 11339
rect 15936 11296 15988 11305
rect 18144 11296 18196 11348
rect 18604 11339 18656 11348
rect 18604 11305 18613 11339
rect 18613 11305 18647 11339
rect 18647 11305 18656 11339
rect 18604 11296 18656 11305
rect 16580 11228 16632 11280
rect 16856 11228 16908 11280
rect 20076 11296 20128 11348
rect 20352 11296 20404 11348
rect 23204 11296 23256 11348
rect 25964 11296 26016 11348
rect 26148 11339 26200 11348
rect 26148 11305 26157 11339
rect 26157 11305 26191 11339
rect 26191 11305 26200 11339
rect 26148 11296 26200 11305
rect 30656 11339 30708 11348
rect 3700 11092 3752 11144
rect 4620 11135 4672 11144
rect 4620 11101 4654 11135
rect 4654 11101 4672 11135
rect 4620 11092 4672 11101
rect 8300 11092 8352 11144
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8944 11135 8996 11144
rect 8392 11092 8444 11101
rect 8944 11101 8953 11135
rect 8953 11101 8987 11135
rect 8987 11101 8996 11135
rect 8944 11092 8996 11101
rect 11704 11160 11756 11212
rect 13452 11203 13504 11212
rect 13452 11169 13461 11203
rect 13461 11169 13495 11203
rect 13495 11169 13504 11203
rect 13452 11160 13504 11169
rect 14188 11203 14240 11212
rect 14188 11169 14197 11203
rect 14197 11169 14231 11203
rect 14231 11169 14240 11203
rect 14188 11160 14240 11169
rect 15752 11160 15804 11212
rect 17868 11160 17920 11212
rect 10508 11092 10560 11144
rect 12256 11092 12308 11144
rect 12532 11092 12584 11144
rect 14096 11092 14148 11144
rect 16672 11135 16724 11144
rect 5172 11024 5224 11076
rect 6828 11024 6880 11076
rect 9036 11024 9088 11076
rect 9588 11024 9640 11076
rect 10416 11024 10468 11076
rect 11244 11067 11296 11076
rect 11244 11033 11253 11067
rect 11253 11033 11287 11067
rect 11287 11033 11296 11067
rect 11244 11024 11296 11033
rect 14004 11024 14056 11076
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 19892 11092 19944 11144
rect 15476 11024 15528 11076
rect 18328 11024 18380 11076
rect 10232 10956 10284 11008
rect 12440 10956 12492 11008
rect 12624 10956 12676 11008
rect 15844 10956 15896 11008
rect 16028 10956 16080 11008
rect 16580 10956 16632 11008
rect 19340 10956 19392 11008
rect 19708 11024 19760 11076
rect 20444 11160 20496 11212
rect 22100 11160 22152 11212
rect 23204 11160 23256 11212
rect 23296 11160 23348 11212
rect 27436 11228 27488 11280
rect 29736 11228 29788 11280
rect 22376 11092 22428 11144
rect 23572 11092 23624 11144
rect 24768 11092 24820 11144
rect 25136 11092 25188 11144
rect 26516 11160 26568 11212
rect 22284 11024 22336 11076
rect 26240 11024 26292 11076
rect 26976 11092 27028 11144
rect 27620 11092 27672 11144
rect 30012 11228 30064 11280
rect 30012 11135 30064 11144
rect 30012 11101 30021 11135
rect 30021 11101 30055 11135
rect 30055 11101 30064 11135
rect 30012 11092 30064 11101
rect 30380 11024 30432 11076
rect 30656 11305 30665 11339
rect 30665 11305 30699 11339
rect 30699 11305 30708 11339
rect 30656 11296 30708 11305
rect 33416 11296 33468 11348
rect 30840 11228 30892 11280
rect 30656 11135 30708 11144
rect 30656 11101 30665 11135
rect 30665 11101 30699 11135
rect 30699 11101 30708 11135
rect 30656 11092 30708 11101
rect 30748 11135 30800 11144
rect 30748 11101 30757 11135
rect 30757 11101 30791 11135
rect 30791 11101 30800 11135
rect 30748 11092 30800 11101
rect 31944 11092 31996 11144
rect 32312 11135 32364 11144
rect 32312 11101 32321 11135
rect 32321 11101 32355 11135
rect 32355 11101 32364 11135
rect 32312 11092 32364 11101
rect 33692 11160 33744 11212
rect 34612 11160 34664 11212
rect 32588 11092 32640 11144
rect 34980 11135 35032 11144
rect 34980 11101 34989 11135
rect 34989 11101 35023 11135
rect 35023 11101 35032 11135
rect 34980 11092 35032 11101
rect 40592 11296 40644 11348
rect 41052 11339 41104 11348
rect 41052 11305 41061 11339
rect 41061 11305 41095 11339
rect 41095 11305 41104 11339
rect 41052 11296 41104 11305
rect 42064 11339 42116 11348
rect 42064 11305 42073 11339
rect 42073 11305 42107 11339
rect 42107 11305 42116 11339
rect 42064 11296 42116 11305
rect 37464 11228 37516 11280
rect 37004 11160 37056 11212
rect 37924 11203 37976 11212
rect 37924 11169 37933 11203
rect 37933 11169 37967 11203
rect 37967 11169 37976 11203
rect 37924 11160 37976 11169
rect 35624 11024 35676 11076
rect 37188 11067 37240 11076
rect 37188 11033 37197 11067
rect 37197 11033 37231 11067
rect 37231 11033 37240 11067
rect 37188 11024 37240 11033
rect 37556 11092 37608 11144
rect 19892 10956 19944 11008
rect 20628 10956 20680 11008
rect 22376 10956 22428 11008
rect 23664 10999 23716 11008
rect 23664 10965 23673 10999
rect 23673 10965 23707 10999
rect 23707 10965 23716 10999
rect 23664 10956 23716 10965
rect 24768 10999 24820 11008
rect 24768 10965 24777 10999
rect 24777 10965 24811 10999
rect 24811 10965 24820 10999
rect 24768 10956 24820 10965
rect 25228 10956 25280 11008
rect 27252 10956 27304 11008
rect 30196 10956 30248 11008
rect 36728 10999 36780 11008
rect 36728 10965 36737 10999
rect 36737 10965 36771 10999
rect 36771 10965 36780 10999
rect 36728 10956 36780 10965
rect 38568 11092 38620 11144
rect 38660 11092 38712 11144
rect 39948 11228 40000 11280
rect 41328 11160 41380 11212
rect 41512 11203 41564 11212
rect 41512 11169 41521 11203
rect 41521 11169 41555 11203
rect 41555 11169 41564 11203
rect 41512 11160 41564 11169
rect 42708 11160 42760 11212
rect 37740 11024 37792 11076
rect 37832 10956 37884 11008
rect 39764 11024 39816 11076
rect 40224 11135 40276 11144
rect 40224 11101 40233 11135
rect 40233 11101 40267 11135
rect 40267 11101 40276 11135
rect 40224 11092 40276 11101
rect 40408 11135 40460 11144
rect 40408 11101 40417 11135
rect 40417 11101 40451 11135
rect 40451 11101 40460 11135
rect 40408 11092 40460 11101
rect 40960 11092 41012 11144
rect 41420 11135 41472 11144
rect 41420 11101 41429 11135
rect 41429 11101 41463 11135
rect 41463 11101 41472 11135
rect 41420 11092 41472 11101
rect 41972 11135 42024 11144
rect 41972 11101 41981 11135
rect 41981 11101 42015 11135
rect 42015 11101 42024 11135
rect 41972 11092 42024 11101
rect 42432 11092 42484 11144
rect 41512 11024 41564 11076
rect 42524 11024 42576 11076
rect 40132 10956 40184 11008
rect 41052 10956 41104 11008
rect 42892 10956 42944 11008
rect 43536 10999 43588 11008
rect 43536 10965 43545 10999
rect 43545 10965 43579 10999
rect 43579 10965 43588 10999
rect 43536 10956 43588 10965
rect 11898 10854 11950 10906
rect 11962 10854 12014 10906
rect 12026 10854 12078 10906
rect 12090 10854 12142 10906
rect 12154 10854 12206 10906
rect 22846 10854 22898 10906
rect 22910 10854 22962 10906
rect 22974 10854 23026 10906
rect 23038 10854 23090 10906
rect 23102 10854 23154 10906
rect 33794 10854 33846 10906
rect 33858 10854 33910 10906
rect 33922 10854 33974 10906
rect 33986 10854 34038 10906
rect 34050 10854 34102 10906
rect 44742 10854 44794 10906
rect 44806 10854 44858 10906
rect 44870 10854 44922 10906
rect 44934 10854 44986 10906
rect 44998 10854 45050 10906
rect 3332 10752 3384 10804
rect 2780 10684 2832 10736
rect 6276 10752 6328 10804
rect 8024 10752 8076 10804
rect 4436 10684 4488 10736
rect 10600 10752 10652 10804
rect 10324 10684 10376 10736
rect 2872 10591 2924 10600
rect 2872 10557 2881 10591
rect 2881 10557 2915 10591
rect 2915 10557 2924 10591
rect 2872 10548 2924 10557
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 2228 10455 2280 10464
rect 2228 10421 2237 10455
rect 2237 10421 2271 10455
rect 2271 10421 2280 10455
rect 2228 10412 2280 10421
rect 3884 10616 3936 10668
rect 10692 10616 10744 10668
rect 14188 10752 14240 10804
rect 14280 10752 14332 10804
rect 14832 10795 14884 10804
rect 14832 10761 14841 10795
rect 14841 10761 14875 10795
rect 14875 10761 14884 10795
rect 14832 10752 14884 10761
rect 15476 10752 15528 10804
rect 15844 10752 15896 10804
rect 22008 10752 22060 10804
rect 22376 10752 22428 10804
rect 26240 10795 26292 10804
rect 26240 10761 26249 10795
rect 26249 10761 26283 10795
rect 26283 10761 26292 10795
rect 26240 10752 26292 10761
rect 32312 10752 32364 10804
rect 37004 10752 37056 10804
rect 13360 10727 13412 10736
rect 13360 10693 13369 10727
rect 13369 10693 13403 10727
rect 13403 10693 13412 10727
rect 13360 10684 13412 10693
rect 15016 10684 15068 10736
rect 15292 10659 15344 10668
rect 15292 10625 15301 10659
rect 15301 10625 15335 10659
rect 15335 10625 15344 10659
rect 15292 10616 15344 10625
rect 7288 10591 7340 10600
rect 7288 10557 7297 10591
rect 7297 10557 7331 10591
rect 7331 10557 7340 10591
rect 7288 10548 7340 10557
rect 9588 10548 9640 10600
rect 10416 10548 10468 10600
rect 4988 10480 5040 10532
rect 10232 10480 10284 10532
rect 14556 10548 14608 10600
rect 21916 10684 21968 10736
rect 20996 10659 21048 10668
rect 20996 10625 21005 10659
rect 21005 10625 21039 10659
rect 21039 10625 21048 10659
rect 20996 10616 21048 10625
rect 23020 10659 23072 10668
rect 23020 10625 23029 10659
rect 23029 10625 23063 10659
rect 23063 10625 23072 10659
rect 23020 10616 23072 10625
rect 24676 10684 24728 10736
rect 24768 10727 24820 10736
rect 24768 10693 24777 10727
rect 24777 10693 24811 10727
rect 24811 10693 24820 10727
rect 24768 10684 24820 10693
rect 25228 10684 25280 10736
rect 28724 10616 28776 10668
rect 28816 10616 28868 10668
rect 32588 10659 32640 10668
rect 32588 10625 32597 10659
rect 32597 10625 32631 10659
rect 32631 10625 32640 10659
rect 32588 10616 32640 10625
rect 18512 10548 18564 10600
rect 22284 10591 22336 10600
rect 22284 10557 22293 10591
rect 22293 10557 22327 10591
rect 22327 10557 22336 10591
rect 22284 10548 22336 10557
rect 22468 10591 22520 10600
rect 22468 10557 22477 10591
rect 22477 10557 22511 10591
rect 22511 10557 22520 10591
rect 22468 10548 22520 10557
rect 30288 10591 30340 10600
rect 30288 10557 30297 10591
rect 30297 10557 30331 10591
rect 30331 10557 30340 10591
rect 30288 10548 30340 10557
rect 35808 10616 35860 10668
rect 35992 10659 36044 10668
rect 35992 10625 36001 10659
rect 36001 10625 36035 10659
rect 36035 10625 36044 10659
rect 35992 10616 36044 10625
rect 39672 10752 39724 10804
rect 41420 10752 41472 10804
rect 38292 10727 38344 10736
rect 38292 10693 38301 10727
rect 38301 10693 38335 10727
rect 38335 10693 38344 10727
rect 38292 10684 38344 10693
rect 42892 10727 42944 10736
rect 42892 10693 42901 10727
rect 42901 10693 42935 10727
rect 42935 10693 42944 10727
rect 42892 10684 42944 10693
rect 5080 10412 5132 10464
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 8208 10412 8260 10464
rect 8944 10412 8996 10464
rect 9220 10412 9272 10464
rect 21732 10480 21784 10532
rect 21916 10480 21968 10532
rect 15476 10412 15528 10464
rect 15568 10412 15620 10464
rect 17776 10455 17828 10464
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 17776 10412 17828 10421
rect 22468 10412 22520 10464
rect 23204 10412 23256 10464
rect 25780 10480 25832 10532
rect 34980 10548 35032 10600
rect 36544 10548 36596 10600
rect 37464 10591 37516 10600
rect 37464 10557 37473 10591
rect 37473 10557 37507 10591
rect 37507 10557 37516 10591
rect 37464 10548 37516 10557
rect 37648 10591 37700 10600
rect 37648 10557 37657 10591
rect 37657 10557 37691 10591
rect 37691 10557 37700 10591
rect 37648 10548 37700 10557
rect 34060 10480 34112 10532
rect 37280 10480 37332 10532
rect 37372 10523 37424 10532
rect 37372 10489 37381 10523
rect 37381 10489 37415 10523
rect 37415 10489 37424 10523
rect 39120 10616 39172 10668
rect 40500 10616 40552 10668
rect 41604 10659 41656 10668
rect 38476 10548 38528 10600
rect 41052 10591 41104 10600
rect 37372 10480 37424 10489
rect 40500 10480 40552 10532
rect 41052 10557 41061 10591
rect 41061 10557 41095 10591
rect 41095 10557 41104 10591
rect 41052 10548 41104 10557
rect 41236 10480 41288 10532
rect 41604 10625 41613 10659
rect 41613 10625 41647 10659
rect 41647 10625 41656 10659
rect 41604 10616 41656 10625
rect 42800 10659 42852 10668
rect 42800 10625 42809 10659
rect 42809 10625 42843 10659
rect 42843 10625 42852 10659
rect 42800 10616 42852 10625
rect 43536 10616 43588 10668
rect 44180 10659 44232 10668
rect 44180 10625 44189 10659
rect 44189 10625 44223 10659
rect 44223 10625 44232 10659
rect 44180 10616 44232 10625
rect 43352 10548 43404 10600
rect 32496 10412 32548 10464
rect 32772 10412 32824 10464
rect 40592 10455 40644 10464
rect 40592 10421 40601 10455
rect 40601 10421 40635 10455
rect 40635 10421 40644 10455
rect 40592 10412 40644 10421
rect 40776 10412 40828 10464
rect 42708 10412 42760 10464
rect 6424 10310 6476 10362
rect 6488 10310 6540 10362
rect 6552 10310 6604 10362
rect 6616 10310 6668 10362
rect 6680 10310 6732 10362
rect 17372 10310 17424 10362
rect 17436 10310 17488 10362
rect 17500 10310 17552 10362
rect 17564 10310 17616 10362
rect 17628 10310 17680 10362
rect 28320 10310 28372 10362
rect 28384 10310 28436 10362
rect 28448 10310 28500 10362
rect 28512 10310 28564 10362
rect 28576 10310 28628 10362
rect 39268 10310 39320 10362
rect 39332 10310 39384 10362
rect 39396 10310 39448 10362
rect 39460 10310 39512 10362
rect 39524 10310 39576 10362
rect 2872 10208 2924 10260
rect 4988 10208 5040 10260
rect 5080 10208 5132 10260
rect 9036 10208 9088 10260
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 12348 10208 12400 10260
rect 10692 10140 10744 10192
rect 12440 10140 12492 10192
rect 8300 10072 8352 10124
rect 9496 10072 9548 10124
rect 12348 10072 12400 10124
rect 13084 10208 13136 10260
rect 14556 10208 14608 10260
rect 15016 10251 15068 10260
rect 15016 10217 15025 10251
rect 15025 10217 15059 10251
rect 15059 10217 15068 10251
rect 15016 10208 15068 10217
rect 19708 10251 19760 10260
rect 19708 10217 19717 10251
rect 19717 10217 19751 10251
rect 19751 10217 19760 10251
rect 19708 10208 19760 10217
rect 15752 10115 15804 10124
rect 3240 10004 3292 10056
rect 4436 10004 4488 10056
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 9404 10004 9456 10056
rect 11336 10004 11388 10056
rect 2228 9936 2280 9988
rect 6828 9936 6880 9988
rect 8484 9936 8536 9988
rect 10416 9936 10468 9988
rect 15752 10081 15761 10115
rect 15761 10081 15795 10115
rect 15795 10081 15804 10115
rect 15752 10072 15804 10081
rect 22284 10208 22336 10260
rect 23020 10208 23072 10260
rect 25228 10208 25280 10260
rect 27252 10208 27304 10260
rect 26976 10140 27028 10192
rect 33232 10208 33284 10260
rect 35624 10251 35676 10260
rect 35624 10217 35633 10251
rect 35633 10217 35667 10251
rect 35667 10217 35676 10251
rect 35624 10208 35676 10217
rect 35808 10208 35860 10260
rect 20628 10115 20680 10124
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 7380 9911 7432 9920
rect 7380 9877 7389 9911
rect 7389 9877 7423 9911
rect 7423 9877 7432 9911
rect 7380 9868 7432 9877
rect 12256 9868 12308 9920
rect 12440 9868 12492 9920
rect 12992 9868 13044 9920
rect 13636 9868 13688 9920
rect 18328 10004 18380 10056
rect 20628 10081 20637 10115
rect 20637 10081 20671 10115
rect 20671 10081 20680 10115
rect 20628 10072 20680 10081
rect 21732 10072 21784 10124
rect 19892 10047 19944 10056
rect 19892 10013 19901 10047
rect 19901 10013 19935 10047
rect 19935 10013 19944 10047
rect 19892 10004 19944 10013
rect 21180 10004 21232 10056
rect 22008 10004 22060 10056
rect 25228 10004 25280 10056
rect 25412 10047 25464 10056
rect 25412 10013 25421 10047
rect 25421 10013 25455 10047
rect 25455 10013 25464 10047
rect 25412 10004 25464 10013
rect 26700 10047 26752 10056
rect 26700 10013 26709 10047
rect 26709 10013 26743 10047
rect 26743 10013 26752 10047
rect 26700 10004 26752 10013
rect 26976 10047 27028 10056
rect 26976 10013 26985 10047
rect 26985 10013 27019 10047
rect 27019 10013 27028 10047
rect 26976 10004 27028 10013
rect 27528 10004 27580 10056
rect 28816 10072 28868 10124
rect 30288 10072 30340 10124
rect 34152 10072 34204 10124
rect 16028 9979 16080 9988
rect 16028 9945 16037 9979
rect 16037 9945 16071 9979
rect 16071 9945 16080 9979
rect 16028 9936 16080 9945
rect 17776 9936 17828 9988
rect 25136 9936 25188 9988
rect 27620 9936 27672 9988
rect 34520 10004 34572 10056
rect 34796 10004 34848 10056
rect 36176 10047 36228 10056
rect 36176 10013 36185 10047
rect 36185 10013 36219 10047
rect 36219 10013 36228 10047
rect 36176 10004 36228 10013
rect 37556 10140 37608 10192
rect 39672 10208 39724 10260
rect 40132 10208 40184 10260
rect 40316 10251 40368 10260
rect 40316 10217 40325 10251
rect 40325 10217 40359 10251
rect 40359 10217 40368 10251
rect 40316 10208 40368 10217
rect 40500 10251 40552 10260
rect 40500 10217 40509 10251
rect 40509 10217 40543 10251
rect 40543 10217 40552 10251
rect 40500 10208 40552 10217
rect 40592 10208 40644 10260
rect 37924 10115 37976 10124
rect 37924 10081 37933 10115
rect 37933 10081 37967 10115
rect 37967 10081 37976 10115
rect 37924 10072 37976 10081
rect 41972 10072 42024 10124
rect 38476 10004 38528 10056
rect 40132 10047 40184 10056
rect 40132 10013 40141 10047
rect 40141 10013 40175 10047
rect 40175 10013 40184 10047
rect 40132 10004 40184 10013
rect 40316 10047 40368 10056
rect 40316 10013 40325 10047
rect 40325 10013 40359 10047
rect 40359 10013 40368 10047
rect 40316 10004 40368 10013
rect 40684 10004 40736 10056
rect 41144 10047 41196 10056
rect 41144 10013 41151 10047
rect 41151 10013 41196 10047
rect 41144 10004 41196 10013
rect 15292 9868 15344 9920
rect 16672 9868 16724 9920
rect 18328 9868 18380 9920
rect 18512 9868 18564 9920
rect 18696 9868 18748 9920
rect 22100 9868 22152 9920
rect 24952 9868 25004 9920
rect 26332 9868 26384 9920
rect 27436 9868 27488 9920
rect 28448 9868 28500 9920
rect 29920 9936 29972 9988
rect 30380 9936 30432 9988
rect 30012 9868 30064 9920
rect 32496 9936 32548 9988
rect 36544 9936 36596 9988
rect 37648 9936 37700 9988
rect 38844 9936 38896 9988
rect 41328 10047 41380 10056
rect 41328 10013 41337 10047
rect 41337 10013 41371 10047
rect 41371 10013 41380 10047
rect 41328 10004 41380 10013
rect 41512 10004 41564 10056
rect 42064 10004 42116 10056
rect 42800 10208 42852 10260
rect 42340 10047 42392 10056
rect 42340 10013 42349 10047
rect 42349 10013 42383 10047
rect 42383 10013 42392 10047
rect 42340 10004 42392 10013
rect 43444 10004 43496 10056
rect 41972 9936 42024 9988
rect 35072 9911 35124 9920
rect 35072 9877 35081 9911
rect 35081 9877 35115 9911
rect 35115 9877 35124 9911
rect 35072 9868 35124 9877
rect 39028 9868 39080 9920
rect 40868 9868 40920 9920
rect 42156 9868 42208 9920
rect 43628 9868 43680 9920
rect 11898 9766 11950 9818
rect 11962 9766 12014 9818
rect 12026 9766 12078 9818
rect 12090 9766 12142 9818
rect 12154 9766 12206 9818
rect 22846 9766 22898 9818
rect 22910 9766 22962 9818
rect 22974 9766 23026 9818
rect 23038 9766 23090 9818
rect 23102 9766 23154 9818
rect 33794 9766 33846 9818
rect 33858 9766 33910 9818
rect 33922 9766 33974 9818
rect 33986 9766 34038 9818
rect 34050 9766 34102 9818
rect 44742 9766 44794 9818
rect 44806 9766 44858 9818
rect 44870 9766 44922 9818
rect 44934 9766 44986 9818
rect 44998 9766 45050 9818
rect 3516 9596 3568 9648
rect 4896 9596 4948 9648
rect 12256 9664 12308 9716
rect 3424 9528 3476 9580
rect 3240 9435 3292 9444
rect 3240 9401 3249 9435
rect 3249 9401 3283 9435
rect 3283 9401 3292 9435
rect 3240 9392 3292 9401
rect 2780 9324 2832 9376
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 11060 9596 11112 9648
rect 12440 9596 12492 9648
rect 12900 9596 12952 9648
rect 15752 9664 15804 9716
rect 19892 9664 19944 9716
rect 25136 9707 25188 9716
rect 25136 9673 25145 9707
rect 25145 9673 25179 9707
rect 25179 9673 25188 9707
rect 25136 9664 25188 9673
rect 25228 9664 25280 9716
rect 27528 9664 27580 9716
rect 30012 9664 30064 9716
rect 6828 9528 6880 9537
rect 8208 9528 8260 9580
rect 9496 9571 9548 9580
rect 9496 9537 9505 9571
rect 9505 9537 9539 9571
rect 9539 9537 9548 9571
rect 9496 9528 9548 9537
rect 3700 9503 3752 9512
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 6920 9503 6972 9512
rect 3700 9460 3752 9469
rect 6920 9469 6929 9503
rect 6929 9469 6963 9503
rect 6963 9469 6972 9503
rect 12348 9528 12400 9580
rect 12992 9571 13044 9580
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 13544 9528 13596 9580
rect 16672 9571 16724 9580
rect 16672 9537 16681 9571
rect 16681 9537 16715 9571
rect 16715 9537 16724 9571
rect 16672 9528 16724 9537
rect 18052 9596 18104 9648
rect 18512 9596 18564 9648
rect 19340 9596 19392 9648
rect 20628 9596 20680 9648
rect 23664 9639 23716 9648
rect 23664 9605 23673 9639
rect 23673 9605 23707 9639
rect 23707 9605 23716 9639
rect 23664 9596 23716 9605
rect 24952 9596 25004 9648
rect 28448 9596 28500 9648
rect 19432 9528 19484 9580
rect 25412 9528 25464 9580
rect 30380 9528 30432 9580
rect 31576 9596 31628 9648
rect 34888 9664 34940 9716
rect 35072 9664 35124 9716
rect 31116 9528 31168 9580
rect 32680 9571 32732 9580
rect 32680 9537 32689 9571
rect 32689 9537 32723 9571
rect 32723 9537 32732 9571
rect 32680 9528 32732 9537
rect 32772 9571 32824 9580
rect 32772 9537 32781 9571
rect 32781 9537 32815 9571
rect 32815 9537 32824 9571
rect 32772 9528 32824 9537
rect 33232 9528 33284 9580
rect 33416 9528 33468 9580
rect 35808 9571 35860 9580
rect 6920 9460 6972 9469
rect 15844 9503 15896 9512
rect 15844 9469 15853 9503
rect 15853 9469 15887 9503
rect 15887 9469 15896 9503
rect 15844 9460 15896 9469
rect 15936 9503 15988 9512
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 15936 9460 15988 9469
rect 16396 9460 16448 9512
rect 17040 9460 17092 9512
rect 3976 9324 4028 9376
rect 5540 9367 5592 9376
rect 5540 9333 5549 9367
rect 5549 9333 5583 9367
rect 5583 9333 5592 9367
rect 5540 9324 5592 9333
rect 5724 9324 5776 9376
rect 8208 9367 8260 9376
rect 8208 9333 8217 9367
rect 8217 9333 8251 9367
rect 8251 9333 8260 9367
rect 8208 9324 8260 9333
rect 9312 9324 9364 9376
rect 17132 9392 17184 9444
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 21732 9460 21784 9512
rect 22008 9460 22060 9512
rect 23388 9503 23440 9512
rect 21180 9392 21232 9444
rect 23388 9469 23397 9503
rect 23397 9469 23431 9503
rect 23431 9469 23440 9503
rect 23388 9460 23440 9469
rect 26240 9460 26292 9512
rect 11336 9324 11388 9376
rect 11520 9367 11572 9376
rect 11520 9333 11529 9367
rect 11529 9333 11563 9367
rect 11563 9333 11572 9367
rect 11520 9324 11572 9333
rect 14648 9324 14700 9376
rect 16488 9324 16540 9376
rect 16672 9324 16724 9376
rect 19708 9324 19760 9376
rect 21272 9324 21324 9376
rect 27804 9460 27856 9512
rect 29644 9503 29696 9512
rect 29644 9469 29653 9503
rect 29653 9469 29687 9503
rect 29687 9469 29696 9503
rect 29644 9460 29696 9469
rect 29828 9324 29880 9376
rect 33140 9460 33192 9512
rect 34244 9460 34296 9512
rect 34520 9460 34572 9512
rect 35808 9537 35817 9571
rect 35817 9537 35851 9571
rect 35851 9537 35860 9571
rect 35808 9528 35860 9537
rect 35900 9571 35952 9580
rect 35900 9537 35909 9571
rect 35909 9537 35943 9571
rect 35943 9537 35952 9571
rect 38660 9639 38712 9648
rect 38660 9605 38669 9639
rect 38669 9605 38703 9639
rect 38703 9605 38712 9639
rect 38660 9596 38712 9605
rect 39120 9664 39172 9716
rect 40776 9664 40828 9716
rect 41236 9707 41288 9716
rect 41236 9673 41245 9707
rect 41245 9673 41279 9707
rect 41279 9673 41288 9707
rect 41236 9664 41288 9673
rect 39672 9596 39724 9648
rect 35900 9528 35952 9537
rect 36544 9571 36596 9580
rect 36544 9537 36553 9571
rect 36553 9537 36587 9571
rect 36587 9537 36596 9571
rect 36544 9528 36596 9537
rect 38568 9571 38620 9580
rect 38568 9537 38577 9571
rect 38577 9537 38611 9571
rect 38611 9537 38620 9571
rect 38568 9528 38620 9537
rect 38752 9528 38804 9580
rect 33600 9392 33652 9444
rect 38936 9460 38988 9512
rect 39856 9460 39908 9512
rect 40132 9528 40184 9580
rect 42340 9664 42392 9716
rect 40960 9571 41012 9580
rect 40960 9537 40969 9571
rect 40969 9537 41003 9571
rect 41003 9537 41012 9571
rect 40960 9528 41012 9537
rect 41328 9528 41380 9580
rect 43352 9596 43404 9648
rect 42616 9571 42668 9580
rect 42616 9537 42625 9571
rect 42625 9537 42659 9571
rect 42659 9537 42668 9571
rect 42616 9528 42668 9537
rect 42708 9571 42760 9580
rect 42708 9537 42717 9571
rect 42717 9537 42751 9571
rect 42751 9537 42760 9571
rect 42708 9528 42760 9537
rect 43444 9571 43496 9580
rect 42064 9460 42116 9512
rect 42524 9460 42576 9512
rect 35808 9392 35860 9444
rect 38476 9392 38528 9444
rect 40224 9392 40276 9444
rect 43444 9537 43453 9571
rect 43453 9537 43487 9571
rect 43487 9537 43496 9571
rect 43444 9528 43496 9537
rect 43628 9571 43680 9580
rect 43628 9537 43637 9571
rect 43637 9537 43671 9571
rect 43671 9537 43680 9571
rect 43628 9528 43680 9537
rect 43352 9392 43404 9444
rect 34428 9324 34480 9376
rect 34704 9367 34756 9376
rect 34704 9333 34713 9367
rect 34713 9333 34747 9367
rect 34747 9333 34756 9367
rect 34704 9324 34756 9333
rect 34796 9324 34848 9376
rect 40132 9324 40184 9376
rect 40868 9324 40920 9376
rect 41512 9324 41564 9376
rect 41696 9367 41748 9376
rect 41696 9333 41705 9367
rect 41705 9333 41739 9367
rect 41739 9333 41748 9367
rect 41696 9324 41748 9333
rect 6424 9222 6476 9274
rect 6488 9222 6540 9274
rect 6552 9222 6604 9274
rect 6616 9222 6668 9274
rect 6680 9222 6732 9274
rect 17372 9222 17424 9274
rect 17436 9222 17488 9274
rect 17500 9222 17552 9274
rect 17564 9222 17616 9274
rect 17628 9222 17680 9274
rect 28320 9222 28372 9274
rect 28384 9222 28436 9274
rect 28448 9222 28500 9274
rect 28512 9222 28564 9274
rect 28576 9222 28628 9274
rect 39268 9222 39320 9274
rect 39332 9222 39384 9274
rect 39396 9222 39448 9274
rect 39460 9222 39512 9274
rect 39524 9222 39576 9274
rect 3424 9120 3476 9172
rect 5724 9120 5776 9172
rect 6828 9120 6880 9172
rect 12440 9120 12492 9172
rect 12992 9120 13044 9172
rect 27804 9163 27856 9172
rect 4344 9052 4396 9104
rect 6276 9095 6328 9104
rect 6276 9061 6285 9095
rect 6285 9061 6319 9095
rect 6319 9061 6328 9095
rect 6276 9052 6328 9061
rect 8208 9052 8260 9104
rect 17040 9095 17092 9104
rect 17040 9061 17049 9095
rect 17049 9061 17083 9095
rect 17083 9061 17092 9095
rect 17040 9052 17092 9061
rect 21180 9095 21232 9104
rect 21180 9061 21189 9095
rect 21189 9061 21223 9095
rect 21223 9061 21232 9095
rect 21180 9052 21232 9061
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 4160 8916 4212 8968
rect 2780 8848 2832 8900
rect 3056 8780 3108 8832
rect 5080 8916 5132 8968
rect 6920 8984 6972 9036
rect 7288 8984 7340 9036
rect 10508 8984 10560 9036
rect 14648 9027 14700 9036
rect 14648 8993 14657 9027
rect 14657 8993 14691 9027
rect 14691 8993 14700 9027
rect 14648 8984 14700 8993
rect 14740 8984 14792 9036
rect 19708 9027 19760 9036
rect 19708 8993 19717 9027
rect 19717 8993 19751 9027
rect 19751 8993 19760 9027
rect 19708 8984 19760 8993
rect 20720 8984 20772 9036
rect 27804 9129 27813 9163
rect 27813 9129 27847 9163
rect 27847 9129 27856 9163
rect 27804 9120 27856 9129
rect 30380 9163 30432 9172
rect 30380 9129 30389 9163
rect 30389 9129 30423 9163
rect 30423 9129 30432 9163
rect 30380 9120 30432 9129
rect 32772 9120 32824 9172
rect 35072 9163 35124 9172
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 7840 8959 7892 8968
rect 7840 8925 7849 8959
rect 7849 8925 7883 8959
rect 7883 8925 7892 8959
rect 7840 8916 7892 8925
rect 7472 8848 7524 8900
rect 9680 8916 9732 8968
rect 11704 8916 11756 8968
rect 13084 8916 13136 8968
rect 16672 8916 16724 8968
rect 18052 8916 18104 8968
rect 19248 8916 19300 8968
rect 28724 8984 28776 9036
rect 24584 8959 24636 8968
rect 10416 8848 10468 8900
rect 10876 8891 10928 8900
rect 10876 8857 10910 8891
rect 10910 8857 10928 8891
rect 10876 8848 10928 8857
rect 15292 8848 15344 8900
rect 15568 8891 15620 8900
rect 15568 8857 15577 8891
rect 15577 8857 15611 8891
rect 15611 8857 15620 8891
rect 15568 8848 15620 8857
rect 8760 8780 8812 8832
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 13268 8823 13320 8832
rect 13268 8789 13277 8823
rect 13277 8789 13311 8823
rect 13311 8789 13320 8823
rect 13268 8780 13320 8789
rect 15476 8780 15528 8832
rect 22100 8891 22152 8900
rect 22100 8857 22109 8891
rect 22109 8857 22143 8891
rect 22143 8857 22152 8891
rect 22100 8848 22152 8857
rect 22744 8780 22796 8832
rect 24584 8925 24593 8959
rect 24593 8925 24627 8959
rect 24627 8925 24636 8959
rect 24584 8916 24636 8925
rect 24492 8848 24544 8900
rect 27436 8916 27488 8968
rect 27620 8916 27672 8968
rect 28448 8916 28500 8968
rect 26240 8848 26292 8900
rect 26332 8891 26384 8900
rect 26332 8857 26341 8891
rect 26341 8857 26375 8891
rect 26375 8857 26384 8891
rect 29828 8916 29880 8968
rect 26332 8848 26384 8857
rect 29552 8848 29604 8900
rect 31576 9052 31628 9104
rect 31668 9052 31720 9104
rect 31944 8984 31996 9036
rect 32312 8984 32364 9036
rect 35072 9129 35081 9163
rect 35081 9129 35115 9163
rect 35115 9129 35124 9163
rect 35072 9120 35124 9129
rect 38200 9163 38252 9172
rect 38200 9129 38209 9163
rect 38209 9129 38243 9163
rect 38243 9129 38252 9163
rect 38200 9120 38252 9129
rect 38844 9163 38896 9172
rect 38844 9129 38853 9163
rect 38853 9129 38887 9163
rect 38887 9129 38896 9163
rect 38844 9120 38896 9129
rect 40132 9120 40184 9172
rect 43352 9120 43404 9172
rect 34888 9052 34940 9104
rect 34980 8984 35032 9036
rect 35900 8984 35952 9036
rect 39120 9052 39172 9104
rect 39856 9052 39908 9104
rect 42156 9095 42208 9104
rect 39580 8984 39632 9036
rect 30748 8959 30800 8968
rect 30748 8925 30757 8959
rect 30757 8925 30791 8959
rect 30791 8925 30800 8959
rect 30748 8916 30800 8925
rect 31484 8916 31536 8968
rect 31576 8959 31628 8968
rect 31576 8925 31585 8959
rect 31585 8925 31619 8959
rect 31619 8925 31628 8959
rect 31576 8916 31628 8925
rect 34704 8916 34756 8968
rect 34888 8959 34940 8968
rect 34888 8925 34897 8959
rect 34897 8925 34931 8959
rect 34931 8925 34940 8959
rect 34888 8916 34940 8925
rect 33692 8848 33744 8900
rect 34428 8848 34480 8900
rect 38568 8916 38620 8968
rect 39028 8959 39080 8968
rect 39028 8925 39037 8959
rect 39037 8925 39071 8959
rect 39071 8925 39080 8959
rect 39028 8916 39080 8925
rect 39672 8916 39724 8968
rect 40040 8959 40092 8968
rect 40040 8925 40049 8959
rect 40049 8925 40083 8959
rect 40083 8925 40092 8959
rect 40040 8916 40092 8925
rect 25044 8780 25096 8832
rect 25228 8823 25280 8832
rect 25228 8789 25237 8823
rect 25237 8789 25271 8823
rect 25271 8789 25280 8823
rect 25228 8780 25280 8789
rect 26700 8780 26752 8832
rect 27620 8780 27672 8832
rect 28908 8823 28960 8832
rect 28908 8789 28917 8823
rect 28917 8789 28951 8823
rect 28951 8789 28960 8823
rect 28908 8780 28960 8789
rect 29000 8780 29052 8832
rect 31668 8780 31720 8832
rect 32680 8780 32732 8832
rect 34520 8780 34572 8832
rect 34704 8823 34756 8832
rect 34704 8789 34713 8823
rect 34713 8789 34747 8823
rect 34747 8789 34756 8823
rect 34704 8780 34756 8789
rect 38660 8848 38712 8900
rect 39212 8780 39264 8832
rect 39304 8780 39356 8832
rect 40224 8848 40276 8900
rect 40500 8916 40552 8968
rect 40776 8848 40828 8900
rect 41512 8916 41564 8968
rect 42156 9061 42165 9095
rect 42165 9061 42199 9095
rect 42199 9061 42208 9095
rect 42156 9052 42208 9061
rect 42616 8959 42668 8968
rect 42616 8925 42625 8959
rect 42625 8925 42659 8959
rect 42659 8925 42668 8959
rect 42616 8916 42668 8925
rect 42800 8780 42852 8832
rect 11898 8678 11950 8730
rect 11962 8678 12014 8730
rect 12026 8678 12078 8730
rect 12090 8678 12142 8730
rect 12154 8678 12206 8730
rect 22846 8678 22898 8730
rect 22910 8678 22962 8730
rect 22974 8678 23026 8730
rect 23038 8678 23090 8730
rect 23102 8678 23154 8730
rect 33794 8678 33846 8730
rect 33858 8678 33910 8730
rect 33922 8678 33974 8730
rect 33986 8678 34038 8730
rect 34050 8678 34102 8730
rect 44742 8678 44794 8730
rect 44806 8678 44858 8730
rect 44870 8678 44922 8730
rect 44934 8678 44986 8730
rect 44998 8678 45050 8730
rect 3056 8619 3108 8628
rect 3056 8585 3065 8619
rect 3065 8585 3099 8619
rect 3099 8585 3108 8619
rect 3056 8576 3108 8585
rect 3148 8576 3200 8628
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 7656 8576 7708 8628
rect 9864 8576 9916 8628
rect 10600 8619 10652 8628
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 13084 8619 13136 8628
rect 13084 8585 13093 8619
rect 13093 8585 13127 8619
rect 13127 8585 13136 8619
rect 13084 8576 13136 8585
rect 13544 8619 13596 8628
rect 13544 8585 13553 8619
rect 13553 8585 13587 8619
rect 13587 8585 13596 8619
rect 13544 8576 13596 8585
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 3148 8440 3200 8492
rect 3240 8440 3292 8492
rect 4344 8440 4396 8492
rect 5356 8440 5408 8492
rect 6828 8440 6880 8492
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 9312 8440 9364 8492
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 11796 8440 11848 8492
rect 14740 8483 14792 8492
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 14740 8440 14792 8449
rect 15292 8440 15344 8492
rect 15568 8440 15620 8492
rect 15844 8576 15896 8628
rect 19432 8619 19484 8628
rect 19432 8585 19441 8619
rect 19441 8585 19475 8619
rect 19475 8585 19484 8619
rect 19432 8576 19484 8585
rect 16488 8508 16540 8560
rect 25596 8576 25648 8628
rect 22376 8508 22428 8560
rect 17960 8440 18012 8492
rect 21088 8440 21140 8492
rect 21272 8483 21324 8492
rect 21272 8449 21281 8483
rect 21281 8449 21315 8483
rect 21315 8449 21324 8483
rect 21272 8440 21324 8449
rect 23204 8440 23256 8492
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 4988 8372 5040 8424
rect 7472 8372 7524 8424
rect 14188 8415 14240 8424
rect 14188 8381 14197 8415
rect 14197 8381 14231 8415
rect 14231 8381 14240 8415
rect 14188 8372 14240 8381
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 20352 8415 20404 8424
rect 20352 8381 20361 8415
rect 20361 8381 20395 8415
rect 20395 8381 20404 8415
rect 20352 8372 20404 8381
rect 20444 8372 20496 8424
rect 21824 8415 21876 8424
rect 21824 8381 21833 8415
rect 21833 8381 21867 8415
rect 21867 8381 21876 8415
rect 21824 8372 21876 8381
rect 27712 8508 27764 8560
rect 28448 8551 28500 8560
rect 28448 8517 28457 8551
rect 28457 8517 28491 8551
rect 28491 8517 28500 8551
rect 28448 8508 28500 8517
rect 28908 8508 28960 8560
rect 5816 8347 5868 8356
rect 5816 8313 5825 8347
rect 5825 8313 5859 8347
rect 5859 8313 5868 8347
rect 5816 8304 5868 8313
rect 6828 8304 6880 8356
rect 8576 8279 8628 8288
rect 8576 8245 8585 8279
rect 8585 8245 8619 8279
rect 8619 8245 8628 8279
rect 8576 8236 8628 8245
rect 10784 8236 10836 8288
rect 13360 8236 13412 8288
rect 13452 8236 13504 8288
rect 19892 8279 19944 8288
rect 19892 8245 19901 8279
rect 19901 8245 19935 8279
rect 19935 8245 19944 8279
rect 19892 8236 19944 8245
rect 25044 8440 25096 8492
rect 27344 8483 27396 8492
rect 24492 8415 24544 8424
rect 24492 8381 24501 8415
rect 24501 8381 24535 8415
rect 24535 8381 24544 8415
rect 24492 8372 24544 8381
rect 20444 8236 20496 8288
rect 27344 8449 27353 8483
rect 27353 8449 27387 8483
rect 27387 8449 27396 8483
rect 27344 8440 27396 8449
rect 29000 8483 29052 8492
rect 25596 8372 25648 8424
rect 29000 8449 29009 8483
rect 29009 8449 29043 8483
rect 29043 8449 29052 8483
rect 29000 8440 29052 8449
rect 29552 8440 29604 8492
rect 29828 8440 29880 8492
rect 30012 8483 30064 8492
rect 30012 8449 30021 8483
rect 30021 8449 30055 8483
rect 30055 8449 30064 8483
rect 30012 8440 30064 8449
rect 33692 8576 33744 8628
rect 34796 8576 34848 8628
rect 34888 8576 34940 8628
rect 38936 8576 38988 8628
rect 40500 8576 40552 8628
rect 32128 8440 32180 8492
rect 32404 8483 32456 8492
rect 32404 8449 32413 8483
rect 32413 8449 32447 8483
rect 32447 8449 32456 8483
rect 32404 8440 32456 8449
rect 33048 8440 33100 8492
rect 34704 8440 34756 8492
rect 37372 8483 37424 8492
rect 37372 8449 37381 8483
rect 37381 8449 37415 8483
rect 37415 8449 37424 8483
rect 37372 8440 37424 8449
rect 38200 8440 38252 8492
rect 27528 8415 27580 8424
rect 27528 8381 27537 8415
rect 27537 8381 27571 8415
rect 27571 8381 27580 8415
rect 27528 8372 27580 8381
rect 28816 8372 28868 8424
rect 38476 8440 38528 8492
rect 38936 8440 38988 8492
rect 39856 8508 39908 8560
rect 42800 8551 42852 8560
rect 39304 8483 39356 8492
rect 39304 8449 39338 8483
rect 39338 8449 39356 8483
rect 39304 8440 39356 8449
rect 39580 8440 39632 8492
rect 42800 8517 42809 8551
rect 42809 8517 42843 8551
rect 42843 8517 42852 8551
rect 42800 8508 42852 8517
rect 41236 8440 41288 8492
rect 43260 8483 43312 8492
rect 43260 8449 43269 8483
rect 43269 8449 43303 8483
rect 43303 8449 43312 8483
rect 43260 8440 43312 8449
rect 44180 8483 44232 8492
rect 44180 8449 44189 8483
rect 44189 8449 44223 8483
rect 44223 8449 44232 8483
rect 44180 8440 44232 8449
rect 31484 8304 31536 8356
rect 32496 8304 32548 8356
rect 33508 8304 33560 8356
rect 26976 8279 27028 8288
rect 26976 8245 26985 8279
rect 26985 8245 27019 8279
rect 27019 8245 27028 8279
rect 26976 8236 27028 8245
rect 30288 8279 30340 8288
rect 30288 8245 30297 8279
rect 30297 8245 30331 8279
rect 30331 8245 30340 8279
rect 30288 8236 30340 8245
rect 32864 8236 32916 8288
rect 34980 8347 35032 8356
rect 34980 8313 34989 8347
rect 34989 8313 35023 8347
rect 35023 8313 35032 8347
rect 34980 8304 35032 8313
rect 38752 8304 38804 8356
rect 34612 8236 34664 8288
rect 40408 8372 40460 8424
rect 41144 8415 41196 8424
rect 41144 8381 41153 8415
rect 41153 8381 41187 8415
rect 41187 8381 41196 8415
rect 41144 8372 41196 8381
rect 41512 8372 41564 8424
rect 42524 8372 42576 8424
rect 42616 8304 42668 8356
rect 6424 8134 6476 8186
rect 6488 8134 6540 8186
rect 6552 8134 6604 8186
rect 6616 8134 6668 8186
rect 6680 8134 6732 8186
rect 17372 8134 17424 8186
rect 17436 8134 17488 8186
rect 17500 8134 17552 8186
rect 17564 8134 17616 8186
rect 17628 8134 17680 8186
rect 28320 8134 28372 8186
rect 28384 8134 28436 8186
rect 28448 8134 28500 8186
rect 28512 8134 28564 8186
rect 28576 8134 28628 8186
rect 39268 8134 39320 8186
rect 39332 8134 39384 8186
rect 39396 8134 39448 8186
rect 39460 8134 39512 8186
rect 39524 8134 39576 8186
rect 5356 8075 5408 8084
rect 5356 8041 5365 8075
rect 5365 8041 5399 8075
rect 5399 8041 5408 8075
rect 5356 8032 5408 8041
rect 7840 8075 7892 8084
rect 7840 8041 7849 8075
rect 7849 8041 7883 8075
rect 7883 8041 7892 8075
rect 7840 8032 7892 8041
rect 10876 8032 10928 8084
rect 13360 8032 13412 8084
rect 15568 8075 15620 8084
rect 15568 8041 15577 8075
rect 15577 8041 15611 8075
rect 15611 8041 15620 8075
rect 15568 8032 15620 8041
rect 15936 8032 15988 8084
rect 18696 8032 18748 8084
rect 19892 8032 19944 8084
rect 21088 8075 21140 8084
rect 21088 8041 21097 8075
rect 21097 8041 21131 8075
rect 21131 8041 21140 8075
rect 21088 8032 21140 8041
rect 16028 8007 16080 8016
rect 16028 7973 16037 8007
rect 16037 7973 16071 8007
rect 16071 7973 16080 8007
rect 16028 7964 16080 7973
rect 16488 7964 16540 8016
rect 11704 7896 11756 7948
rect 17500 7896 17552 7948
rect 4068 7828 4120 7880
rect 7012 7828 7064 7880
rect 9680 7828 9732 7880
rect 11520 7828 11572 7880
rect 13360 7828 13412 7880
rect 14740 7828 14792 7880
rect 15384 7828 15436 7880
rect 16672 7828 16724 7880
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 19248 7871 19300 7880
rect 19248 7837 19257 7871
rect 19257 7837 19291 7871
rect 19291 7837 19300 7871
rect 19248 7828 19300 7837
rect 22376 7896 22428 7948
rect 22284 7828 22336 7880
rect 23388 8032 23440 8084
rect 24584 8032 24636 8084
rect 32864 8032 32916 8084
rect 40040 8032 40092 8084
rect 41236 8075 41288 8084
rect 41236 8041 41245 8075
rect 41245 8041 41279 8075
rect 41279 8041 41288 8075
rect 41236 8032 41288 8041
rect 42708 8032 42760 8084
rect 33232 7964 33284 8016
rect 26240 7896 26292 7948
rect 27712 7896 27764 7948
rect 28816 7939 28868 7948
rect 28816 7905 28825 7939
rect 28825 7905 28859 7939
rect 28859 7905 28868 7939
rect 28816 7896 28868 7905
rect 33508 7896 33560 7948
rect 24492 7828 24544 7880
rect 25228 7828 25280 7880
rect 29736 7871 29788 7880
rect 29736 7837 29745 7871
rect 29745 7837 29779 7871
rect 29779 7837 29788 7871
rect 29736 7828 29788 7837
rect 30288 7828 30340 7880
rect 32220 7828 32272 7880
rect 5540 7760 5592 7812
rect 6276 7760 6328 7812
rect 8576 7760 8628 7812
rect 11060 7760 11112 7812
rect 11704 7692 11756 7744
rect 13268 7735 13320 7744
rect 13268 7701 13277 7735
rect 13277 7701 13311 7735
rect 13311 7701 13320 7735
rect 22652 7760 22704 7812
rect 13268 7692 13320 7701
rect 19340 7692 19392 7744
rect 26148 7692 26200 7744
rect 26332 7760 26384 7812
rect 32312 7760 32364 7812
rect 33692 7828 33744 7880
rect 34612 7828 34664 7880
rect 38936 7896 38988 7948
rect 39856 7939 39908 7948
rect 39120 7871 39172 7880
rect 32496 7760 32548 7812
rect 39120 7837 39129 7871
rect 39129 7837 39163 7871
rect 39163 7837 39172 7871
rect 39120 7828 39172 7837
rect 39856 7905 39865 7939
rect 39865 7905 39899 7939
rect 39899 7905 39908 7939
rect 39856 7896 39908 7905
rect 41144 7896 41196 7948
rect 39396 7828 39448 7880
rect 41880 7871 41932 7880
rect 41880 7837 41889 7871
rect 41889 7837 41923 7871
rect 41923 7837 41932 7871
rect 41880 7828 41932 7837
rect 42616 7828 42668 7880
rect 44180 7871 44232 7880
rect 44180 7837 44189 7871
rect 44189 7837 44223 7871
rect 44223 7837 44232 7871
rect 44180 7828 44232 7837
rect 39856 7760 39908 7812
rect 28264 7735 28316 7744
rect 28264 7701 28273 7735
rect 28273 7701 28307 7735
rect 28307 7701 28316 7735
rect 28264 7692 28316 7701
rect 28816 7692 28868 7744
rect 30012 7692 30064 7744
rect 32128 7692 32180 7744
rect 34704 7735 34756 7744
rect 34704 7701 34713 7735
rect 34713 7701 34747 7735
rect 34747 7701 34756 7735
rect 34704 7692 34756 7701
rect 40408 7692 40460 7744
rect 41144 7692 41196 7744
rect 11898 7590 11950 7642
rect 11962 7590 12014 7642
rect 12026 7590 12078 7642
rect 12090 7590 12142 7642
rect 12154 7590 12206 7642
rect 22846 7590 22898 7642
rect 22910 7590 22962 7642
rect 22974 7590 23026 7642
rect 23038 7590 23090 7642
rect 23102 7590 23154 7642
rect 33794 7590 33846 7642
rect 33858 7590 33910 7642
rect 33922 7590 33974 7642
rect 33986 7590 34038 7642
rect 34050 7590 34102 7642
rect 44742 7590 44794 7642
rect 44806 7590 44858 7642
rect 44870 7590 44922 7642
rect 44934 7590 44986 7642
rect 44998 7590 45050 7642
rect 3516 7488 3568 7540
rect 5172 7488 5224 7540
rect 12808 7488 12860 7540
rect 15384 7488 15436 7540
rect 15476 7488 15528 7540
rect 19340 7488 19392 7540
rect 20352 7488 20404 7540
rect 22652 7531 22704 7540
rect 7380 7420 7432 7472
rect 9496 7463 9548 7472
rect 9496 7429 9505 7463
rect 9505 7429 9539 7463
rect 9539 7429 9548 7463
rect 9496 7420 9548 7429
rect 10784 7420 10836 7472
rect 11704 7420 11756 7472
rect 19248 7420 19300 7472
rect 13360 7395 13412 7404
rect 13360 7361 13369 7395
rect 13369 7361 13403 7395
rect 13403 7361 13412 7395
rect 13360 7352 13412 7361
rect 14096 7352 14148 7404
rect 18328 7395 18380 7404
rect 18328 7361 18362 7395
rect 18362 7361 18380 7395
rect 21824 7420 21876 7472
rect 22652 7497 22661 7531
rect 22661 7497 22695 7531
rect 22695 7497 22704 7531
rect 22652 7488 22704 7497
rect 22744 7488 22796 7540
rect 26148 7531 26200 7540
rect 26148 7497 26157 7531
rect 26157 7497 26191 7531
rect 26191 7497 26200 7531
rect 26148 7488 26200 7497
rect 27344 7488 27396 7540
rect 28816 7488 28868 7540
rect 29644 7488 29696 7540
rect 32588 7488 32640 7540
rect 34704 7488 34756 7540
rect 39856 7531 39908 7540
rect 39856 7497 39865 7531
rect 39865 7497 39899 7531
rect 39899 7497 39908 7531
rect 39856 7488 39908 7497
rect 40776 7531 40828 7540
rect 40776 7497 40785 7531
rect 40785 7497 40819 7531
rect 40819 7497 40828 7531
rect 40776 7488 40828 7497
rect 18328 7352 18380 7361
rect 20168 7395 20220 7404
rect 20168 7361 20202 7395
rect 20202 7361 20220 7395
rect 20168 7352 20220 7361
rect 23296 7352 23348 7404
rect 28264 7420 28316 7472
rect 24032 7395 24084 7404
rect 24032 7361 24041 7395
rect 24041 7361 24075 7395
rect 24075 7361 24084 7395
rect 24032 7352 24084 7361
rect 26976 7352 27028 7404
rect 30012 7420 30064 7472
rect 32312 7420 32364 7472
rect 33416 7420 33468 7472
rect 35808 7420 35860 7472
rect 28724 7352 28776 7404
rect 30380 7352 30432 7404
rect 32128 7395 32180 7404
rect 12348 7327 12400 7336
rect 12348 7293 12357 7327
rect 12357 7293 12391 7327
rect 12391 7293 12400 7327
rect 12348 7284 12400 7293
rect 15660 7327 15712 7336
rect 15660 7293 15669 7327
rect 15669 7293 15703 7327
rect 15703 7293 15712 7327
rect 15660 7284 15712 7293
rect 17500 7327 17552 7336
rect 16672 7216 16724 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 11244 7148 11296 7200
rect 11704 7191 11756 7200
rect 11704 7157 11713 7191
rect 11713 7157 11747 7191
rect 11747 7157 11756 7191
rect 11704 7148 11756 7157
rect 16856 7191 16908 7200
rect 16856 7157 16865 7191
rect 16865 7157 16899 7191
rect 16899 7157 16908 7191
rect 16856 7148 16908 7157
rect 17500 7293 17509 7327
rect 17509 7293 17543 7327
rect 17543 7293 17552 7327
rect 17500 7284 17552 7293
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 21364 7216 21416 7268
rect 26056 7284 26108 7336
rect 27712 7327 27764 7336
rect 27712 7293 27721 7327
rect 27721 7293 27755 7327
rect 27755 7293 27764 7327
rect 27712 7284 27764 7293
rect 29920 7284 29972 7336
rect 32128 7361 32137 7395
rect 32137 7361 32171 7395
rect 32171 7361 32180 7395
rect 32128 7352 32180 7361
rect 32220 7352 32272 7404
rect 32680 7352 32732 7404
rect 33048 7395 33100 7404
rect 33048 7361 33057 7395
rect 33057 7361 33091 7395
rect 33091 7361 33100 7395
rect 33048 7352 33100 7361
rect 39396 7395 39448 7404
rect 39396 7361 39405 7395
rect 39405 7361 39439 7395
rect 39439 7361 39448 7395
rect 39396 7352 39448 7361
rect 39948 7352 40000 7404
rect 40316 7395 40368 7404
rect 31300 7284 31352 7336
rect 35348 7284 35400 7336
rect 40316 7361 40325 7395
rect 40325 7361 40359 7395
rect 40359 7361 40368 7395
rect 40316 7352 40368 7361
rect 40960 7395 41012 7404
rect 40960 7361 40969 7395
rect 40969 7361 41003 7395
rect 41003 7361 41012 7395
rect 40960 7352 41012 7361
rect 41144 7395 41196 7404
rect 41144 7361 41153 7395
rect 41153 7361 41187 7395
rect 41187 7361 41196 7395
rect 41144 7352 41196 7361
rect 41512 7352 41564 7404
rect 40408 7284 40460 7336
rect 43904 7284 43956 7336
rect 26148 7216 26200 7268
rect 18696 7148 18748 7200
rect 20812 7148 20864 7200
rect 22376 7148 22428 7200
rect 25780 7148 25832 7200
rect 31024 7191 31076 7200
rect 31024 7157 31033 7191
rect 31033 7157 31067 7191
rect 31067 7157 31076 7191
rect 31024 7148 31076 7157
rect 32772 7148 32824 7200
rect 34796 7191 34848 7200
rect 34796 7157 34805 7191
rect 34805 7157 34839 7191
rect 34839 7157 34848 7191
rect 34796 7148 34848 7157
rect 41880 7148 41932 7200
rect 6424 7046 6476 7098
rect 6488 7046 6540 7098
rect 6552 7046 6604 7098
rect 6616 7046 6668 7098
rect 6680 7046 6732 7098
rect 17372 7046 17424 7098
rect 17436 7046 17488 7098
rect 17500 7046 17552 7098
rect 17564 7046 17616 7098
rect 17628 7046 17680 7098
rect 28320 7046 28372 7098
rect 28384 7046 28436 7098
rect 28448 7046 28500 7098
rect 28512 7046 28564 7098
rect 28576 7046 28628 7098
rect 39268 7046 39320 7098
rect 39332 7046 39384 7098
rect 39396 7046 39448 7098
rect 39460 7046 39512 7098
rect 39524 7046 39576 7098
rect 7012 6851 7064 6860
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 5816 6740 5868 6792
rect 15660 6944 15712 6996
rect 18328 6944 18380 6996
rect 18696 6944 18748 6996
rect 23296 6987 23348 6996
rect 12348 6876 12400 6928
rect 20260 6876 20312 6928
rect 23296 6953 23305 6987
rect 23305 6953 23339 6987
rect 23339 6953 23348 6987
rect 23296 6944 23348 6953
rect 26056 6944 26108 6996
rect 27712 6944 27764 6996
rect 28816 6944 28868 6996
rect 32588 6944 32640 6996
rect 40960 6944 41012 6996
rect 6000 6672 6052 6724
rect 8208 6672 8260 6724
rect 9680 6740 9732 6792
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 10784 6783 10836 6792
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 14740 6740 14792 6792
rect 16856 6808 16908 6860
rect 16948 6808 17000 6860
rect 31116 6876 31168 6928
rect 21364 6851 21416 6860
rect 21364 6817 21373 6851
rect 21373 6817 21407 6851
rect 21407 6817 21416 6851
rect 21364 6808 21416 6817
rect 26240 6808 26292 6860
rect 26976 6851 27028 6860
rect 26976 6817 26985 6851
rect 26985 6817 27019 6851
rect 27019 6817 27028 6851
rect 26976 6808 27028 6817
rect 29736 6808 29788 6860
rect 31300 6808 31352 6860
rect 8944 6715 8996 6724
rect 8944 6681 8953 6715
rect 8953 6681 8987 6715
rect 8987 6681 8996 6715
rect 8944 6672 8996 6681
rect 9036 6672 9088 6724
rect 10324 6672 10376 6724
rect 15752 6740 15804 6792
rect 20812 6740 20864 6792
rect 25780 6783 25832 6792
rect 25780 6749 25789 6783
rect 25789 6749 25823 6783
rect 25823 6749 25832 6783
rect 25780 6740 25832 6749
rect 26148 6740 26200 6792
rect 32680 6851 32732 6860
rect 32680 6817 32689 6851
rect 32689 6817 32723 6851
rect 32723 6817 32732 6851
rect 32680 6808 32732 6817
rect 39948 6808 40000 6860
rect 33232 6740 33284 6792
rect 40132 6740 40184 6792
rect 9128 6604 9180 6656
rect 12256 6604 12308 6656
rect 14280 6604 14332 6656
rect 20720 6647 20772 6656
rect 20720 6613 20729 6647
rect 20729 6613 20763 6647
rect 20763 6613 20772 6647
rect 20720 6604 20772 6613
rect 21088 6647 21140 6656
rect 21088 6613 21097 6647
rect 21097 6613 21131 6647
rect 21131 6613 21140 6647
rect 21088 6604 21140 6613
rect 22284 6672 22336 6724
rect 27344 6672 27396 6724
rect 22376 6604 22428 6656
rect 26240 6604 26292 6656
rect 26424 6604 26476 6656
rect 29092 6604 29144 6656
rect 30472 6604 30524 6656
rect 32036 6672 32088 6724
rect 11898 6502 11950 6554
rect 11962 6502 12014 6554
rect 12026 6502 12078 6554
rect 12090 6502 12142 6554
rect 12154 6502 12206 6554
rect 22846 6502 22898 6554
rect 22910 6502 22962 6554
rect 22974 6502 23026 6554
rect 23038 6502 23090 6554
rect 23102 6502 23154 6554
rect 33794 6502 33846 6554
rect 33858 6502 33910 6554
rect 33922 6502 33974 6554
rect 33986 6502 34038 6554
rect 34050 6502 34102 6554
rect 44742 6502 44794 6554
rect 44806 6502 44858 6554
rect 44870 6502 44922 6554
rect 44934 6502 44986 6554
rect 44998 6502 45050 6554
rect 8208 6443 8260 6452
rect 8208 6409 8217 6443
rect 8217 6409 8251 6443
rect 8251 6409 8260 6443
rect 8208 6400 8260 6409
rect 10324 6400 10376 6452
rect 11796 6400 11848 6452
rect 17960 6443 18012 6452
rect 7012 6332 7064 6384
rect 6000 6196 6052 6248
rect 9036 6264 9088 6316
rect 10784 6332 10836 6384
rect 11612 6332 11664 6384
rect 8944 6128 8996 6180
rect 11336 6264 11388 6316
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 11152 6196 11204 6248
rect 15200 6332 15252 6384
rect 14648 6264 14700 6316
rect 17960 6409 17969 6443
rect 17969 6409 18003 6443
rect 18003 6409 18012 6443
rect 17960 6400 18012 6409
rect 21180 6400 21232 6452
rect 18328 6264 18380 6316
rect 20720 6264 20772 6316
rect 21824 6307 21876 6316
rect 21824 6273 21833 6307
rect 21833 6273 21867 6307
rect 21867 6273 21876 6307
rect 21824 6264 21876 6273
rect 29828 6400 29880 6452
rect 31852 6400 31904 6452
rect 10692 6060 10744 6112
rect 10784 6060 10836 6112
rect 11336 6060 11388 6112
rect 11796 6060 11848 6112
rect 13176 6060 13228 6112
rect 16764 6128 16816 6180
rect 21640 6196 21692 6248
rect 23296 6196 23348 6248
rect 19892 6128 19944 6180
rect 21364 6128 21416 6180
rect 24032 6264 24084 6316
rect 26424 6264 26476 6316
rect 26976 6307 27028 6316
rect 26976 6273 26985 6307
rect 26985 6273 27019 6307
rect 27019 6273 27028 6307
rect 26976 6264 27028 6273
rect 30472 6264 30524 6316
rect 31300 6307 31352 6316
rect 31300 6273 31309 6307
rect 31309 6273 31343 6307
rect 31343 6273 31352 6307
rect 31300 6264 31352 6273
rect 26884 6196 26936 6248
rect 29920 6196 29972 6248
rect 31576 6332 31628 6384
rect 35808 6400 35860 6452
rect 32128 6307 32180 6316
rect 32128 6273 32137 6307
rect 32137 6273 32171 6307
rect 32171 6273 32180 6307
rect 32128 6264 32180 6273
rect 32588 6264 32640 6316
rect 32680 6264 32732 6316
rect 34520 6264 34572 6316
rect 35716 6264 35768 6316
rect 34704 6196 34756 6248
rect 15568 6060 15620 6112
rect 16856 6103 16908 6112
rect 16856 6069 16865 6103
rect 16865 6069 16899 6103
rect 16899 6069 16908 6103
rect 16856 6060 16908 6069
rect 21088 6060 21140 6112
rect 22928 6060 22980 6112
rect 24400 6060 24452 6112
rect 30012 6128 30064 6180
rect 29000 6060 29052 6112
rect 29092 6060 29144 6112
rect 31116 6060 31168 6112
rect 33600 6060 33652 6112
rect 6424 5958 6476 6010
rect 6488 5958 6540 6010
rect 6552 5958 6604 6010
rect 6616 5958 6668 6010
rect 6680 5958 6732 6010
rect 17372 5958 17424 6010
rect 17436 5958 17488 6010
rect 17500 5958 17552 6010
rect 17564 5958 17616 6010
rect 17628 5958 17680 6010
rect 28320 5958 28372 6010
rect 28384 5958 28436 6010
rect 28448 5958 28500 6010
rect 28512 5958 28564 6010
rect 28576 5958 28628 6010
rect 39268 5958 39320 6010
rect 39332 5958 39384 6010
rect 39396 5958 39448 6010
rect 39460 5958 39512 6010
rect 39524 5958 39576 6010
rect 10048 5856 10100 5908
rect 11612 5856 11664 5908
rect 11796 5856 11848 5908
rect 12624 5856 12676 5908
rect 15752 5899 15804 5908
rect 15752 5865 15761 5899
rect 15761 5865 15795 5899
rect 15795 5865 15804 5899
rect 15752 5856 15804 5865
rect 18328 5899 18380 5908
rect 18328 5865 18337 5899
rect 18337 5865 18371 5899
rect 18371 5865 18380 5899
rect 18328 5856 18380 5865
rect 23480 5856 23532 5908
rect 11060 5788 11112 5840
rect 11336 5788 11388 5840
rect 8944 5720 8996 5772
rect 16764 5788 16816 5840
rect 16948 5788 17000 5840
rect 7012 5652 7064 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9128 5652 9180 5661
rect 8208 5584 8260 5636
rect 12992 5652 13044 5704
rect 13176 5695 13228 5704
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 11796 5584 11848 5636
rect 13452 5720 13504 5772
rect 26792 5856 26844 5908
rect 26884 5899 26936 5908
rect 26884 5865 26893 5899
rect 26893 5865 26927 5899
rect 26927 5865 26936 5899
rect 26884 5856 26936 5865
rect 30932 5856 30984 5908
rect 31116 5856 31168 5908
rect 34520 5856 34572 5908
rect 34704 5899 34756 5908
rect 34704 5865 34713 5899
rect 34713 5865 34747 5899
rect 34747 5865 34756 5899
rect 34704 5856 34756 5865
rect 35348 5899 35400 5908
rect 35348 5865 35357 5899
rect 35357 5865 35391 5899
rect 35391 5865 35400 5899
rect 35348 5856 35400 5865
rect 20536 5720 20588 5772
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 22928 5720 22980 5729
rect 15568 5695 15620 5704
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 17500 5652 17552 5704
rect 18052 5652 18104 5704
rect 14556 5627 14608 5636
rect 8944 5559 8996 5568
rect 8944 5525 8953 5559
rect 8953 5525 8987 5559
rect 8987 5525 8996 5559
rect 8944 5516 8996 5525
rect 12716 5516 12768 5568
rect 14556 5593 14565 5627
rect 14565 5593 14599 5627
rect 14599 5593 14608 5627
rect 14556 5584 14608 5593
rect 16856 5584 16908 5636
rect 21732 5652 21784 5704
rect 28356 5788 28408 5840
rect 29000 5788 29052 5840
rect 29644 5788 29696 5840
rect 31024 5788 31076 5840
rect 24400 5695 24452 5704
rect 24400 5661 24409 5695
rect 24409 5661 24443 5695
rect 24443 5661 24452 5695
rect 24400 5652 24452 5661
rect 24676 5695 24728 5704
rect 24676 5661 24685 5695
rect 24685 5661 24719 5695
rect 24719 5661 24728 5695
rect 24676 5652 24728 5661
rect 26424 5695 26476 5704
rect 26424 5661 26433 5695
rect 26433 5661 26467 5695
rect 26467 5661 26476 5695
rect 26424 5652 26476 5661
rect 27620 5652 27672 5704
rect 27804 5695 27856 5704
rect 27804 5661 27813 5695
rect 27813 5661 27847 5695
rect 27847 5661 27856 5695
rect 27804 5652 27856 5661
rect 28356 5652 28408 5704
rect 29000 5652 29052 5704
rect 29828 5695 29880 5704
rect 29828 5661 29837 5695
rect 29837 5661 29871 5695
rect 29871 5661 29880 5695
rect 29828 5652 29880 5661
rect 21180 5516 21232 5568
rect 24032 5516 24084 5568
rect 24308 5516 24360 5568
rect 28172 5516 28224 5568
rect 28540 5516 28592 5568
rect 28632 5559 28684 5568
rect 28632 5525 28641 5559
rect 28641 5525 28675 5559
rect 28675 5525 28684 5559
rect 29644 5584 29696 5636
rect 30012 5695 30064 5704
rect 30012 5661 30021 5695
rect 30021 5661 30055 5695
rect 30055 5661 30064 5695
rect 30012 5652 30064 5661
rect 30380 5652 30432 5704
rect 32680 5720 32732 5772
rect 32128 5652 32180 5704
rect 33692 5720 33744 5772
rect 30748 5584 30800 5636
rect 31576 5584 31628 5636
rect 33140 5584 33192 5636
rect 35624 5652 35676 5704
rect 43904 5695 43956 5704
rect 43904 5661 43913 5695
rect 43913 5661 43947 5695
rect 43947 5661 43956 5695
rect 43904 5652 43956 5661
rect 28632 5516 28684 5525
rect 31392 5516 31444 5568
rect 33508 5559 33560 5568
rect 33508 5525 33517 5559
rect 33517 5525 33551 5559
rect 33551 5525 33560 5559
rect 33508 5516 33560 5525
rect 35440 5516 35492 5568
rect 44088 5559 44140 5568
rect 44088 5525 44097 5559
rect 44097 5525 44131 5559
rect 44131 5525 44140 5559
rect 44088 5516 44140 5525
rect 11898 5414 11950 5466
rect 11962 5414 12014 5466
rect 12026 5414 12078 5466
rect 12090 5414 12142 5466
rect 12154 5414 12206 5466
rect 22846 5414 22898 5466
rect 22910 5414 22962 5466
rect 22974 5414 23026 5466
rect 23038 5414 23090 5466
rect 23102 5414 23154 5466
rect 33794 5414 33846 5466
rect 33858 5414 33910 5466
rect 33922 5414 33974 5466
rect 33986 5414 34038 5466
rect 34050 5414 34102 5466
rect 44742 5414 44794 5466
rect 44806 5414 44858 5466
rect 44870 5414 44922 5466
rect 44934 5414 44986 5466
rect 44998 5414 45050 5466
rect 10692 5312 10744 5364
rect 11796 5355 11848 5364
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 12256 5355 12308 5364
rect 12256 5321 12265 5355
rect 12265 5321 12299 5355
rect 12299 5321 12308 5355
rect 12256 5312 12308 5321
rect 13636 5312 13688 5364
rect 8944 5244 8996 5296
rect 7012 5176 7064 5228
rect 11336 5244 11388 5296
rect 12992 5287 13044 5296
rect 12992 5253 13001 5287
rect 13001 5253 13035 5287
rect 13035 5253 13044 5287
rect 12992 5244 13044 5253
rect 10784 5219 10836 5228
rect 10784 5185 10793 5219
rect 10793 5185 10827 5219
rect 10827 5185 10836 5219
rect 10784 5176 10836 5185
rect 16028 5244 16080 5296
rect 17776 5244 17828 5296
rect 19340 5312 19392 5364
rect 19800 5312 19852 5364
rect 14832 5176 14884 5228
rect 17224 5176 17276 5228
rect 17500 5176 17552 5228
rect 20444 5219 20496 5228
rect 20444 5185 20453 5219
rect 20453 5185 20487 5219
rect 20487 5185 20496 5219
rect 20444 5176 20496 5185
rect 20720 5219 20772 5228
rect 20720 5185 20729 5219
rect 20729 5185 20763 5219
rect 20763 5185 20772 5219
rect 20720 5176 20772 5185
rect 23112 5219 23164 5228
rect 23112 5185 23121 5219
rect 23121 5185 23155 5219
rect 23155 5185 23164 5219
rect 23112 5176 23164 5185
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 6276 5108 6328 5160
rect 9864 5108 9916 5160
rect 12348 5151 12400 5160
rect 11152 5040 11204 5092
rect 12348 5117 12357 5151
rect 12357 5117 12391 5151
rect 12391 5117 12400 5151
rect 12348 5108 12400 5117
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 15752 5108 15804 5160
rect 19892 5151 19944 5160
rect 19892 5117 19901 5151
rect 19901 5117 19935 5151
rect 19935 5117 19944 5151
rect 19892 5108 19944 5117
rect 20536 5151 20588 5160
rect 20536 5117 20545 5151
rect 20545 5117 20579 5151
rect 20579 5117 20588 5151
rect 20536 5108 20588 5117
rect 22284 5108 22336 5160
rect 13452 5040 13504 5092
rect 21640 5040 21692 5092
rect 23480 5151 23532 5160
rect 23480 5117 23489 5151
rect 23489 5117 23523 5151
rect 23523 5117 23532 5151
rect 23480 5108 23532 5117
rect 27528 5244 27580 5296
rect 28448 5287 28500 5296
rect 28448 5253 28457 5287
rect 28457 5253 28491 5287
rect 28491 5253 28500 5287
rect 28448 5244 28500 5253
rect 28540 5244 28592 5296
rect 30472 5244 30524 5296
rect 23848 5176 23900 5228
rect 25044 5219 25096 5228
rect 25044 5185 25053 5219
rect 25053 5185 25087 5219
rect 25087 5185 25096 5219
rect 25044 5176 25096 5185
rect 25136 5219 25188 5228
rect 25136 5185 25145 5219
rect 25145 5185 25179 5219
rect 25179 5185 25188 5219
rect 25320 5219 25372 5228
rect 25136 5176 25188 5185
rect 25320 5185 25329 5219
rect 25329 5185 25363 5219
rect 25363 5185 25372 5219
rect 25320 5176 25372 5185
rect 25504 5219 25556 5228
rect 25504 5185 25513 5219
rect 25513 5185 25547 5219
rect 25547 5185 25556 5219
rect 25504 5176 25556 5185
rect 27344 5176 27396 5228
rect 24860 5108 24912 5160
rect 28448 5108 28500 5160
rect 29276 5151 29328 5160
rect 29276 5117 29285 5151
rect 29285 5117 29319 5151
rect 29319 5117 29328 5151
rect 29276 5108 29328 5117
rect 29368 5108 29420 5160
rect 29828 5176 29880 5228
rect 30932 5287 30984 5296
rect 30932 5253 30941 5287
rect 30941 5253 30975 5287
rect 30975 5253 30984 5287
rect 30932 5244 30984 5253
rect 31760 5244 31812 5296
rect 31944 5244 31996 5296
rect 30748 5219 30800 5228
rect 30748 5185 30757 5219
rect 30757 5185 30791 5219
rect 30791 5185 30800 5219
rect 30748 5176 30800 5185
rect 29920 5108 29972 5160
rect 32128 5219 32180 5228
rect 32128 5185 32137 5219
rect 32137 5185 32171 5219
rect 32171 5185 32180 5219
rect 32128 5176 32180 5185
rect 32680 5176 32732 5228
rect 35716 5219 35768 5228
rect 35716 5185 35725 5219
rect 35725 5185 35759 5219
rect 35759 5185 35768 5219
rect 35716 5176 35768 5185
rect 35440 5108 35492 5160
rect 24676 5040 24728 5092
rect 27620 5040 27672 5092
rect 30932 5040 30984 5092
rect 33324 5040 33376 5092
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 15016 4972 15068 5024
rect 18052 4972 18104 5024
rect 19432 4972 19484 5024
rect 22744 4972 22796 5024
rect 23572 4972 23624 5024
rect 24400 4972 24452 5024
rect 28172 4972 28224 5024
rect 31944 4972 31996 5024
rect 32588 4972 32640 5024
rect 42800 5015 42852 5024
rect 42800 4981 42809 5015
rect 42809 4981 42843 5015
rect 42843 4981 42852 5015
rect 42800 4972 42852 4981
rect 6424 4870 6476 4922
rect 6488 4870 6540 4922
rect 6552 4870 6604 4922
rect 6616 4870 6668 4922
rect 6680 4870 6732 4922
rect 17372 4870 17424 4922
rect 17436 4870 17488 4922
rect 17500 4870 17552 4922
rect 17564 4870 17616 4922
rect 17628 4870 17680 4922
rect 28320 4870 28372 4922
rect 28384 4870 28436 4922
rect 28448 4870 28500 4922
rect 28512 4870 28564 4922
rect 28576 4870 28628 4922
rect 39268 4870 39320 4922
rect 39332 4870 39384 4922
rect 39396 4870 39448 4922
rect 39460 4870 39512 4922
rect 39524 4870 39576 4922
rect 11704 4768 11756 4820
rect 12348 4768 12400 4820
rect 14096 4811 14148 4820
rect 14096 4777 14105 4811
rect 14105 4777 14139 4811
rect 14139 4777 14148 4811
rect 14096 4768 14148 4777
rect 17776 4768 17828 4820
rect 20444 4768 20496 4820
rect 24400 4768 24452 4820
rect 24860 4811 24912 4820
rect 24860 4777 24869 4811
rect 24869 4777 24903 4811
rect 24903 4777 24912 4811
rect 24860 4768 24912 4777
rect 25044 4811 25096 4820
rect 25044 4777 25053 4811
rect 25053 4777 25087 4811
rect 25087 4777 25096 4811
rect 25044 4768 25096 4777
rect 25136 4768 25188 4820
rect 26148 4768 26200 4820
rect 26884 4768 26936 4820
rect 29092 4768 29144 4820
rect 29460 4768 29512 4820
rect 32772 4811 32824 4820
rect 11796 4700 11848 4752
rect 20720 4700 20772 4752
rect 29276 4700 29328 4752
rect 32772 4777 32781 4811
rect 32781 4777 32815 4811
rect 32815 4777 32824 4811
rect 32772 4768 32824 4777
rect 33140 4768 33192 4820
rect 33232 4768 33284 4820
rect 35624 4768 35676 4820
rect 9128 4632 9180 4684
rect 11428 4564 11480 4616
rect 11612 4632 11664 4684
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 19340 4675 19392 4684
rect 12716 4564 12768 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 15016 4607 15068 4616
rect 15016 4573 15050 4607
rect 15050 4573 15068 4607
rect 15016 4564 15068 4573
rect 18052 4564 18104 4616
rect 6276 4496 6328 4548
rect 11152 4428 11204 4480
rect 11704 4428 11756 4480
rect 12440 4539 12492 4548
rect 12440 4505 12474 4539
rect 12474 4505 12492 4539
rect 19340 4641 19349 4675
rect 19349 4641 19383 4675
rect 19383 4641 19392 4675
rect 19340 4632 19392 4641
rect 22192 4632 22244 4684
rect 23112 4632 23164 4684
rect 29552 4675 29604 4684
rect 12440 4496 12492 4505
rect 15108 4428 15160 4480
rect 18144 4428 18196 4480
rect 20628 4564 20680 4616
rect 23204 4564 23256 4616
rect 26056 4564 26108 4616
rect 26608 4539 26660 4548
rect 26608 4505 26617 4539
rect 26617 4505 26651 4539
rect 26651 4505 26660 4539
rect 26608 4496 26660 4505
rect 27620 4539 27672 4548
rect 27252 4428 27304 4480
rect 27620 4505 27629 4539
rect 27629 4505 27663 4539
rect 27663 4505 27672 4539
rect 27620 4496 27672 4505
rect 29552 4641 29561 4675
rect 29561 4641 29595 4675
rect 29595 4641 29604 4675
rect 29552 4632 29604 4641
rect 29460 4564 29512 4616
rect 30932 4564 30984 4616
rect 29828 4539 29880 4548
rect 29184 4428 29236 4480
rect 29828 4505 29837 4539
rect 29837 4505 29871 4539
rect 29871 4505 29880 4539
rect 29828 4496 29880 4505
rect 31944 4539 31996 4548
rect 31944 4505 31969 4539
rect 31969 4505 31996 4539
rect 33692 4700 33744 4752
rect 31944 4496 31996 4505
rect 30012 4428 30064 4480
rect 31392 4428 31444 4480
rect 33324 4564 33376 4616
rect 34796 4564 34848 4616
rect 42800 4564 42852 4616
rect 33416 4539 33468 4548
rect 33416 4505 33425 4539
rect 33425 4505 33459 4539
rect 33459 4505 33468 4539
rect 33416 4496 33468 4505
rect 33600 4539 33652 4548
rect 33600 4505 33625 4539
rect 33625 4505 33652 4539
rect 33600 4496 33652 4505
rect 33508 4428 33560 4480
rect 44088 4471 44140 4480
rect 44088 4437 44097 4471
rect 44097 4437 44131 4471
rect 44131 4437 44140 4471
rect 44088 4428 44140 4437
rect 11898 4326 11950 4378
rect 11962 4326 12014 4378
rect 12026 4326 12078 4378
rect 12090 4326 12142 4378
rect 12154 4326 12206 4378
rect 22846 4326 22898 4378
rect 22910 4326 22962 4378
rect 22974 4326 23026 4378
rect 23038 4326 23090 4378
rect 23102 4326 23154 4378
rect 33794 4326 33846 4378
rect 33858 4326 33910 4378
rect 33922 4326 33974 4378
rect 33986 4326 34038 4378
rect 34050 4326 34102 4378
rect 44742 4326 44794 4378
rect 44806 4326 44858 4378
rect 44870 4326 44922 4378
rect 44934 4326 44986 4378
rect 44998 4326 45050 4378
rect 14832 4224 14884 4276
rect 15108 4267 15160 4276
rect 15108 4233 15117 4267
rect 15117 4233 15151 4267
rect 15151 4233 15160 4267
rect 15108 4224 15160 4233
rect 15200 4267 15252 4276
rect 15200 4233 15209 4267
rect 15209 4233 15243 4267
rect 15243 4233 15252 4267
rect 15200 4224 15252 4233
rect 25320 4224 25372 4276
rect 26148 4267 26200 4276
rect 26148 4233 26157 4267
rect 26157 4233 26191 4267
rect 26191 4233 26200 4267
rect 26148 4224 26200 4233
rect 29092 4224 29144 4276
rect 30564 4224 30616 4276
rect 11796 4156 11848 4208
rect 11612 4088 11664 4140
rect 12716 4088 12768 4140
rect 17224 4088 17276 4140
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 14556 4020 14608 4072
rect 18144 4063 18196 4072
rect 18144 4029 18153 4063
rect 18153 4029 18187 4063
rect 18187 4029 18196 4063
rect 18144 4020 18196 4029
rect 19432 4020 19484 4072
rect 22284 4156 22336 4208
rect 24400 4156 24452 4208
rect 24860 4156 24912 4208
rect 24308 4131 24360 4140
rect 24308 4097 24317 4131
rect 24317 4097 24351 4131
rect 24351 4097 24360 4131
rect 24308 4088 24360 4097
rect 12532 3884 12584 3936
rect 16764 3884 16816 3936
rect 17776 3884 17828 3936
rect 19248 3884 19300 3936
rect 23388 4020 23440 4072
rect 25044 4088 25096 4140
rect 26056 4131 26108 4140
rect 24768 4020 24820 4072
rect 26056 4097 26065 4131
rect 26065 4097 26099 4131
rect 26099 4097 26108 4131
rect 26056 4088 26108 4097
rect 27620 4156 27672 4208
rect 28080 4156 28132 4208
rect 31760 4156 31812 4208
rect 26976 4088 27028 4140
rect 29460 4088 29512 4140
rect 30012 4131 30064 4140
rect 30012 4097 30021 4131
rect 30021 4097 30055 4131
rect 30055 4097 30064 4131
rect 30012 4088 30064 4097
rect 31300 4088 31352 4140
rect 33416 4224 33468 4276
rect 32680 4156 32732 4208
rect 32864 4156 32916 4208
rect 27528 4063 27580 4072
rect 27528 4029 27537 4063
rect 27537 4029 27571 4063
rect 27571 4029 27580 4063
rect 27528 4020 27580 4029
rect 27620 4020 27672 4072
rect 29368 4020 29420 4072
rect 22192 3884 22244 3936
rect 22744 3884 22796 3936
rect 23848 3927 23900 3936
rect 23848 3893 23857 3927
rect 23857 3893 23891 3927
rect 23891 3893 23900 3927
rect 23848 3884 23900 3893
rect 25504 3952 25556 4004
rect 25044 3927 25096 3936
rect 25044 3893 25053 3927
rect 25053 3893 25087 3927
rect 25087 3893 25096 3927
rect 25044 3884 25096 3893
rect 29092 3884 29144 3936
rect 31300 3884 31352 3936
rect 43904 3884 43956 3936
rect 6424 3782 6476 3834
rect 6488 3782 6540 3834
rect 6552 3782 6604 3834
rect 6616 3782 6668 3834
rect 6680 3782 6732 3834
rect 17372 3782 17424 3834
rect 17436 3782 17488 3834
rect 17500 3782 17552 3834
rect 17564 3782 17616 3834
rect 17628 3782 17680 3834
rect 28320 3782 28372 3834
rect 28384 3782 28436 3834
rect 28448 3782 28500 3834
rect 28512 3782 28564 3834
rect 28576 3782 28628 3834
rect 39268 3782 39320 3834
rect 39332 3782 39384 3834
rect 39396 3782 39448 3834
rect 39460 3782 39512 3834
rect 39524 3782 39576 3834
rect 12440 3680 12492 3732
rect 18236 3680 18288 3732
rect 23572 3723 23624 3732
rect 11428 3612 11480 3664
rect 23572 3689 23581 3723
rect 23581 3689 23615 3723
rect 23615 3689 23624 3723
rect 23572 3680 23624 3689
rect 23756 3723 23808 3732
rect 23756 3689 23765 3723
rect 23765 3689 23799 3723
rect 23799 3689 23808 3723
rect 23756 3680 23808 3689
rect 24400 3680 24452 3732
rect 27528 3680 27580 3732
rect 28080 3723 28132 3732
rect 28080 3689 28089 3723
rect 28089 3689 28123 3723
rect 28123 3689 28132 3723
rect 28080 3680 28132 3689
rect 29828 3680 29880 3732
rect 30932 3680 30984 3732
rect 33232 3680 33284 3732
rect 23848 3612 23900 3664
rect 24768 3612 24820 3664
rect 12624 3587 12676 3596
rect 12624 3553 12633 3587
rect 12633 3553 12667 3587
rect 12667 3553 12676 3587
rect 12624 3544 12676 3553
rect 12716 3587 12768 3596
rect 12716 3553 12725 3587
rect 12725 3553 12759 3587
rect 12759 3553 12768 3587
rect 16764 3587 16816 3596
rect 12716 3544 12768 3553
rect 16764 3553 16773 3587
rect 16773 3553 16807 3587
rect 16807 3553 16816 3587
rect 16764 3544 16816 3553
rect 19248 3587 19300 3596
rect 19248 3553 19257 3587
rect 19257 3553 19291 3587
rect 19291 3553 19300 3587
rect 19248 3544 19300 3553
rect 22100 3544 22152 3596
rect 1584 3519 1636 3528
rect 1584 3485 1593 3519
rect 1593 3485 1627 3519
rect 1627 3485 1636 3519
rect 1584 3476 1636 3485
rect 11152 3476 11204 3528
rect 12532 3519 12584 3528
rect 12532 3485 12541 3519
rect 12541 3485 12575 3519
rect 12575 3485 12584 3519
rect 12532 3476 12584 3485
rect 12992 3476 13044 3528
rect 15752 3519 15804 3528
rect 15752 3485 15761 3519
rect 15761 3485 15795 3519
rect 15795 3485 15804 3519
rect 15752 3476 15804 3485
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 21732 3476 21784 3528
rect 17132 3408 17184 3460
rect 20168 3408 20220 3460
rect 18144 3340 18196 3392
rect 22744 3476 22796 3528
rect 25044 3408 25096 3460
rect 27252 3476 27304 3528
rect 27988 3519 28040 3528
rect 27988 3485 27997 3519
rect 27997 3485 28031 3519
rect 28031 3485 28040 3519
rect 27988 3476 28040 3485
rect 29092 3476 29144 3528
rect 29184 3476 29236 3528
rect 26608 3340 26660 3392
rect 29368 3340 29420 3392
rect 30564 3544 30616 3596
rect 30932 3519 30984 3528
rect 30932 3485 30941 3519
rect 30941 3485 30975 3519
rect 30975 3485 30984 3519
rect 30932 3476 30984 3485
rect 31760 3519 31812 3528
rect 31760 3485 31769 3519
rect 31769 3485 31803 3519
rect 31803 3485 31812 3519
rect 31760 3476 31812 3485
rect 32588 3476 32640 3528
rect 44180 3519 44232 3528
rect 44180 3485 44189 3519
rect 44189 3485 44223 3519
rect 44223 3485 44232 3519
rect 44180 3476 44232 3485
rect 33508 3340 33560 3392
rect 11898 3238 11950 3290
rect 11962 3238 12014 3290
rect 12026 3238 12078 3290
rect 12090 3238 12142 3290
rect 12154 3238 12206 3290
rect 22846 3238 22898 3290
rect 22910 3238 22962 3290
rect 22974 3238 23026 3290
rect 23038 3238 23090 3290
rect 23102 3238 23154 3290
rect 33794 3238 33846 3290
rect 33858 3238 33910 3290
rect 33922 3238 33974 3290
rect 33986 3238 34038 3290
rect 34050 3238 34102 3290
rect 44742 3238 44794 3290
rect 44806 3238 44858 3290
rect 44870 3238 44922 3290
rect 44934 3238 44986 3290
rect 44998 3238 45050 3290
rect 17132 3136 17184 3188
rect 19616 3136 19668 3188
rect 20168 3179 20220 3188
rect 20168 3145 20177 3179
rect 20177 3145 20211 3179
rect 20211 3145 20220 3179
rect 20168 3136 20220 3145
rect 23204 3136 23256 3188
rect 23388 3136 23440 3188
rect 32864 3136 32916 3188
rect 34152 3136 34204 3188
rect 43260 3179 43312 3188
rect 43260 3145 43269 3179
rect 43269 3145 43303 3179
rect 43303 3145 43312 3179
rect 43260 3136 43312 3145
rect 43444 3136 43496 3188
rect 6828 3000 6880 3052
rect 11244 3000 11296 3052
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 22468 3000 22520 3052
rect 22744 3000 22796 3052
rect 23756 3043 23808 3052
rect 23756 3009 23765 3043
rect 23765 3009 23799 3043
rect 23799 3009 23808 3043
rect 23756 3000 23808 3009
rect 27988 3000 28040 3052
rect 30932 3000 30984 3052
rect 43812 3000 43864 3052
rect 45100 2932 45152 2984
rect 17776 2864 17828 2916
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 6276 2796 6328 2848
rect 14464 2796 14516 2848
rect 22652 2796 22704 2848
rect 35532 2796 35584 2848
rect 6424 2694 6476 2746
rect 6488 2694 6540 2746
rect 6552 2694 6604 2746
rect 6616 2694 6668 2746
rect 6680 2694 6732 2746
rect 17372 2694 17424 2746
rect 17436 2694 17488 2746
rect 17500 2694 17552 2746
rect 17564 2694 17616 2746
rect 17628 2694 17680 2746
rect 28320 2694 28372 2746
rect 28384 2694 28436 2746
rect 28448 2694 28500 2746
rect 28512 2694 28564 2746
rect 28576 2694 28628 2746
rect 39268 2694 39320 2746
rect 39332 2694 39384 2746
rect 39396 2694 39448 2746
rect 39460 2694 39512 2746
rect 39524 2694 39576 2746
rect 12992 2635 13044 2644
rect 12992 2601 13001 2635
rect 13001 2601 13035 2635
rect 13035 2601 13044 2635
rect 12992 2592 13044 2601
rect 35992 2592 36044 2644
rect 37372 2592 37424 2644
rect 15108 2524 15160 2576
rect 20 2456 72 2508
rect 17776 2499 17828 2508
rect 17776 2465 17785 2499
rect 17785 2465 17819 2499
rect 17819 2465 17828 2499
rect 17776 2456 17828 2465
rect 1308 2388 1360 2440
rect 3240 2388 3292 2440
rect 4528 2388 4580 2440
rect 6276 2388 6328 2440
rect 7748 2388 7800 2440
rect 9680 2388 9732 2440
rect 10968 2388 11020 2440
rect 12900 2388 12952 2440
rect 14464 2431 14516 2440
rect 14464 2397 14473 2431
rect 14473 2397 14507 2431
rect 14507 2397 14516 2431
rect 14464 2388 14516 2397
rect 16120 2388 16172 2440
rect 17408 2388 17460 2440
rect 19340 2388 19392 2440
rect 20628 2388 20680 2440
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 23848 2388 23900 2440
rect 25780 2388 25832 2440
rect 27068 2388 27120 2440
rect 29000 2388 29052 2440
rect 30288 2388 30340 2440
rect 35532 2431 35584 2440
rect 35532 2397 35541 2431
rect 35541 2397 35575 2431
rect 35575 2397 35584 2431
rect 35532 2388 35584 2397
rect 36728 2388 36780 2440
rect 38660 2388 38712 2440
rect 39948 2388 40000 2440
rect 43904 2431 43956 2440
rect 43904 2397 43913 2431
rect 43913 2397 43947 2431
rect 43947 2397 43956 2431
rect 43904 2388 43956 2397
rect 19708 2320 19760 2372
rect 6460 2252 6512 2304
rect 9680 2252 9732 2304
rect 14188 2252 14240 2304
rect 22560 2252 22612 2304
rect 27436 2252 27488 2304
rect 32220 2320 32272 2372
rect 41880 2320 41932 2372
rect 32312 2252 32364 2304
rect 35440 2252 35492 2304
rect 44088 2295 44140 2304
rect 44088 2261 44097 2295
rect 44097 2261 44131 2295
rect 44131 2261 44140 2295
rect 44088 2252 44140 2261
rect 11898 2150 11950 2202
rect 11962 2150 12014 2202
rect 12026 2150 12078 2202
rect 12090 2150 12142 2202
rect 12154 2150 12206 2202
rect 22846 2150 22898 2202
rect 22910 2150 22962 2202
rect 22974 2150 23026 2202
rect 23038 2150 23090 2202
rect 23102 2150 23154 2202
rect 33794 2150 33846 2202
rect 33858 2150 33910 2202
rect 33922 2150 33974 2202
rect 33986 2150 34038 2202
rect 34050 2150 34102 2202
rect 44742 2150 44794 2202
rect 44806 2150 44858 2202
rect 44870 2150 44922 2202
rect 44934 2150 44986 2202
rect 44998 2150 45050 2202
<< metal2 >>
rect -10 19200 102 20000
rect 1278 19200 1390 20000
rect 3210 19200 3322 20000
rect 4498 19200 4610 20000
rect 6430 19200 6542 20000
rect 7718 19200 7830 20000
rect 9650 19200 9762 20000
rect 10938 19200 11050 20000
rect 12870 19200 12982 20000
rect 14158 19200 14270 20000
rect 16090 19200 16202 20000
rect 17378 19200 17490 20000
rect 19310 19200 19422 20000
rect 20598 19200 20710 20000
rect 22530 19200 22642 20000
rect 23818 19200 23930 20000
rect 25750 19200 25862 20000
rect 27682 19200 27794 20000
rect 28970 19200 29082 20000
rect 30902 19200 31014 20000
rect 32190 19200 32302 20000
rect 34122 19200 34234 20000
rect 35410 19200 35522 20000
rect 37342 19200 37454 20000
rect 38630 19200 38742 20000
rect 40562 19200 40674 20000
rect 41850 19200 41962 20000
rect 43782 19200 43894 20000
rect 45070 19200 45182 20000
rect 32 16590 60 19200
rect 1320 17270 1348 19200
rect 3252 17270 3280 19200
rect 3974 18456 4030 18465
rect 3974 18391 4030 18400
rect 1308 17264 1360 17270
rect 1308 17206 1360 17212
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2240 17105 2268 17138
rect 2226 17096 2282 17105
rect 2226 17031 2282 17040
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 20 16584 72 16590
rect 20 16526 72 16532
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1596 15065 1624 15302
rect 1582 15056 1638 15065
rect 1582 14991 1638 15000
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1596 13705 1624 13806
rect 3068 13734 3096 16934
rect 3988 16794 4016 18391
rect 4540 17202 4568 19200
rect 6472 17202 6500 19200
rect 7760 17202 7788 19200
rect 9692 17202 9720 19200
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 9680 17196 9732 17202
rect 10980 17184 11008 19200
rect 11898 17436 12206 17445
rect 11898 17434 11904 17436
rect 11960 17434 11984 17436
rect 12040 17434 12064 17436
rect 12120 17434 12144 17436
rect 12200 17434 12206 17436
rect 11960 17382 11962 17434
rect 12142 17382 12144 17434
rect 11898 17380 11904 17382
rect 11960 17380 11984 17382
rect 12040 17380 12064 17382
rect 12120 17380 12144 17382
rect 12200 17380 12206 17382
rect 11898 17371 12206 17380
rect 12912 17202 12940 19200
rect 14200 17202 14228 19200
rect 16132 17202 16160 19200
rect 17420 17338 17448 19200
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 19352 17202 19380 19200
rect 20640 17354 20668 19200
rect 20640 17338 20760 17354
rect 20640 17332 20772 17338
rect 20640 17326 20720 17332
rect 20720 17274 20772 17280
rect 22572 17202 22600 19200
rect 22846 17436 23154 17445
rect 22846 17434 22852 17436
rect 22908 17434 22932 17436
rect 22988 17434 23012 17436
rect 23068 17434 23092 17436
rect 23148 17434 23154 17436
rect 22908 17382 22910 17434
rect 23090 17382 23092 17434
rect 22846 17380 22852 17382
rect 22908 17380 22932 17382
rect 22988 17380 23012 17382
rect 23068 17380 23092 17382
rect 23148 17380 23154 17382
rect 22846 17371 23154 17380
rect 23860 17202 23888 19200
rect 25792 17202 25820 19200
rect 27724 17202 27752 19200
rect 29012 17202 29040 19200
rect 30944 17202 30972 19200
rect 32232 17202 32260 19200
rect 33794 17436 34102 17445
rect 33794 17434 33800 17436
rect 33856 17434 33880 17436
rect 33936 17434 33960 17436
rect 34016 17434 34040 17436
rect 34096 17434 34102 17436
rect 33856 17382 33858 17434
rect 34038 17382 34040 17434
rect 33794 17380 33800 17382
rect 33856 17380 33880 17382
rect 33936 17380 33960 17382
rect 34016 17380 34040 17382
rect 34096 17380 34102 17382
rect 33794 17371 34102 17380
rect 34164 17202 34192 19200
rect 35452 17202 35480 19200
rect 37280 17332 37332 17338
rect 37280 17274 37332 17280
rect 11060 17196 11112 17202
rect 10980 17156 11060 17184
rect 9680 17138 9732 17144
rect 11060 17138 11112 17144
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 25780 17196 25832 17202
rect 25780 17138 25832 17144
rect 27712 17196 27764 17202
rect 27712 17138 27764 17144
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 30932 17196 30984 17202
rect 30932 17138 30984 17144
rect 32220 17196 32272 17202
rect 32220 17138 32272 17144
rect 34152 17196 34204 17202
rect 34152 17138 34204 17144
rect 35440 17196 35492 17202
rect 35440 17138 35492 17144
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3160 14074 3188 15438
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3056 13728 3108 13734
rect 1582 13696 1638 13705
rect 3056 13670 3108 13676
rect 1582 13631 1638 13640
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2608 11898 2636 12174
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2700 11354 2728 12174
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2792 10742 2820 12582
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2976 11218 3004 12038
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 3344 10810 3372 13874
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3712 11150 3740 11766
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 1596 10305 1624 10406
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 2240 9994 2268 10406
rect 2884 10266 2912 10542
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 3252 9450 3280 9998
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 8906 2820 9318
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 8634 3096 8774
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3160 8498 3188 8570
rect 3252 8498 3280 9386
rect 3436 9178 3464 9522
rect 3528 9466 3556 9590
rect 3712 9518 3740 11086
rect 3896 10674 3924 12038
rect 4066 11656 4122 11665
rect 4066 11591 4068 11600
rect 4120 11591 4122 11600
rect 4068 11562 4120 11568
rect 4172 11354 4200 17002
rect 4908 16794 4936 17070
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 6424 16892 6732 16901
rect 6424 16890 6430 16892
rect 6486 16890 6510 16892
rect 6566 16890 6590 16892
rect 6646 16890 6670 16892
rect 6726 16890 6732 16892
rect 6486 16838 6488 16890
rect 6668 16838 6670 16890
rect 6424 16836 6430 16838
rect 6486 16836 6510 16838
rect 6566 16836 6590 16838
rect 6646 16836 6670 16838
rect 6726 16836 6732 16838
rect 6424 16827 6732 16836
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 6424 15804 6732 15813
rect 6424 15802 6430 15804
rect 6486 15802 6510 15804
rect 6566 15802 6590 15804
rect 6646 15802 6670 15804
rect 6726 15802 6732 15804
rect 6486 15750 6488 15802
rect 6668 15750 6670 15802
rect 6424 15748 6430 15750
rect 6486 15748 6510 15750
rect 6566 15748 6590 15750
rect 6646 15748 6670 15750
rect 6726 15748 6732 15750
rect 6424 15739 6732 15748
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 6424 14716 6732 14725
rect 6424 14714 6430 14716
rect 6486 14714 6510 14716
rect 6566 14714 6590 14716
rect 6646 14714 6670 14716
rect 6726 14714 6732 14716
rect 6486 14662 6488 14714
rect 6668 14662 6670 14714
rect 6424 14660 6430 14662
rect 6486 14660 6510 14662
rect 6566 14660 6590 14662
rect 6646 14660 6670 14662
rect 6726 14660 6732 14662
rect 6424 14651 6732 14660
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 7392 14006 7420 14214
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 4448 13326 4476 13942
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4448 12850 4476 13262
rect 5368 12918 5396 13670
rect 6424 13628 6732 13637
rect 6424 13626 6430 13628
rect 6486 13626 6510 13628
rect 6566 13626 6590 13628
rect 6646 13626 6670 13628
rect 6726 13626 6732 13628
rect 6486 13574 6488 13626
rect 6668 13574 6670 13626
rect 6424 13572 6430 13574
rect 6486 13572 6510 13574
rect 6566 13572 6590 13574
rect 6646 13572 6670 13574
rect 6726 13572 6732 13574
rect 6424 13563 6732 13572
rect 7116 13326 7144 13806
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 8036 13258 8064 14214
rect 8404 14074 8432 14554
rect 8772 14346 8800 14826
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8404 13530 8432 14010
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 4448 12306 4476 12786
rect 8404 12782 8432 13466
rect 8588 12918 8616 14214
rect 8772 13734 8800 14282
rect 8956 13938 8984 14758
rect 9140 14346 9168 14826
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 9128 14340 9180 14346
rect 9128 14282 9180 14288
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8680 13394 8708 13670
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8772 12850 8800 13670
rect 8956 13462 8984 13874
rect 9232 13802 9260 14486
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9508 13530 9536 14418
rect 9600 14006 9628 14894
rect 9588 14000 9640 14006
rect 9588 13942 9640 13948
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4264 11218 4292 11630
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4448 10742 4476 12242
rect 5460 11898 5488 12378
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 4632 11150 4660 11834
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 4436 10736 4488 10742
rect 4436 10678 4488 10684
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 4448 10062 4476 10678
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5000 10266 5028 10474
rect 5184 10470 5212 11018
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5092 10266 5120 10406
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4436 10056 4488 10062
rect 4436 9998 4488 10004
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 3700 9512 3752 9518
rect 3528 9460 3700 9466
rect 3528 9454 3752 9460
rect 3528 9438 3740 9454
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 1596 8265 1624 8434
rect 3528 8430 3556 9438
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3988 8974 4016 9318
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 3528 7546 3556 8366
rect 4172 7970 4200 8910
rect 4356 8498 4384 9046
rect 4908 8634 4936 9590
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 5000 8430 5028 10202
rect 5092 8974 5120 10202
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4080 7942 4200 7970
rect 4080 7886 4108 7942
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 5184 7546 5212 10406
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5368 8090 5396 8434
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5552 7818 5580 9318
rect 5736 9178 5764 9318
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6905 1624 7142
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 5828 6798 5856 8298
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 6012 6730 6040 12582
rect 6424 12540 6732 12549
rect 6424 12538 6430 12540
rect 6486 12538 6510 12540
rect 6566 12538 6590 12540
rect 6646 12538 6670 12540
rect 6726 12538 6732 12540
rect 6486 12486 6488 12538
rect 6668 12486 6670 12538
rect 6424 12484 6430 12486
rect 6486 12484 6510 12486
rect 6566 12484 6590 12486
rect 6646 12484 6670 12486
rect 6726 12484 6732 12486
rect 6424 12475 6732 12484
rect 8864 12434 8892 13262
rect 9048 12918 9076 13466
rect 9600 13258 9628 13942
rect 9692 13870 9720 16934
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9784 13734 9812 14350
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 8864 12406 8984 12434
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6564 11626 6592 12106
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6104 10062 6132 11562
rect 6424 11452 6732 11461
rect 6424 11450 6430 11452
rect 6486 11450 6510 11452
rect 6566 11450 6590 11452
rect 6646 11450 6670 11452
rect 6726 11450 6732 11452
rect 6486 11398 6488 11450
rect 6668 11398 6670 11450
rect 6424 11396 6430 11398
rect 6486 11396 6510 11398
rect 6566 11396 6590 11398
rect 6646 11396 6670 11398
rect 6726 11396 6732 11398
rect 6424 11387 6732 11396
rect 6840 11082 6868 12174
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7208 11898 7236 12038
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6288 9110 6316 10746
rect 7300 10606 7328 11494
rect 8036 10810 8064 11494
rect 8220 11354 8248 12310
rect 8956 12238 8984 12406
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8404 11150 8432 11494
rect 8496 11286 8524 11630
rect 8864 11354 8892 12174
rect 8956 11694 8984 12174
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9232 11830 9260 12038
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 6424 10364 6732 10373
rect 6424 10362 6430 10364
rect 6486 10362 6510 10364
rect 6566 10362 6590 10364
rect 6646 10362 6670 10364
rect 6726 10362 6732 10364
rect 6486 10310 6488 10362
rect 6668 10310 6670 10362
rect 6424 10308 6430 10310
rect 6486 10308 6510 10310
rect 6566 10308 6590 10310
rect 6646 10308 6670 10310
rect 6726 10308 6732 10310
rect 6424 10299 6732 10308
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6840 9586 6868 9930
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6748 9466 6776 9522
rect 6920 9512 6972 9518
rect 6748 9438 6868 9466
rect 6920 9454 6972 9460
rect 6424 9276 6732 9285
rect 6424 9274 6430 9276
rect 6486 9274 6510 9276
rect 6566 9274 6590 9276
rect 6646 9274 6670 9276
rect 6726 9274 6732 9276
rect 6486 9222 6488 9274
rect 6668 9222 6670 9274
rect 6424 9220 6430 9222
rect 6486 9220 6510 9222
rect 6566 9220 6590 9222
rect 6646 9220 6670 9222
rect 6726 9220 6732 9222
rect 6424 9211 6732 9220
rect 6840 9178 6868 9438
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 6840 8498 6868 9114
rect 6932 9042 6960 9454
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7300 8498 7328 8978
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6424 8188 6732 8197
rect 6424 8186 6430 8188
rect 6486 8186 6510 8188
rect 6566 8186 6590 8188
rect 6646 8186 6670 8188
rect 6726 8186 6732 8188
rect 6486 8134 6488 8186
rect 6668 8134 6670 8186
rect 6424 8132 6430 8134
rect 6486 8132 6510 8134
rect 6566 8132 6590 8134
rect 6646 8132 6670 8134
rect 6726 8132 6732 8134
rect 6424 8123 6732 8132
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6000 6724 6052 6730
rect 6000 6666 6052 6672
rect 6012 6254 6040 6666
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6288 5166 6316 7754
rect 6424 7100 6732 7109
rect 6424 7098 6430 7100
rect 6486 7098 6510 7100
rect 6566 7098 6590 7100
rect 6646 7098 6670 7100
rect 6726 7098 6732 7100
rect 6486 7046 6488 7098
rect 6668 7046 6670 7098
rect 6424 7044 6430 7046
rect 6486 7044 6510 7046
rect 6566 7044 6590 7046
rect 6646 7044 6670 7046
rect 6726 7044 6732 7046
rect 6424 7035 6732 7044
rect 6424 6012 6732 6021
rect 6424 6010 6430 6012
rect 6486 6010 6510 6012
rect 6566 6010 6590 6012
rect 6646 6010 6670 6012
rect 6726 6010 6732 6012
rect 6486 5958 6488 6010
rect 6668 5958 6670 6010
rect 6424 5956 6430 5958
rect 6486 5956 6510 5958
rect 6566 5956 6590 5958
rect 6646 5956 6670 5958
rect 6726 5956 6732 5958
rect 6424 5947 6732 5956
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 1412 4865 1440 5102
rect 1398 4856 1454 4865
rect 1398 4791 1454 4800
rect 6288 4554 6316 5102
rect 6424 4924 6732 4933
rect 6424 4922 6430 4924
rect 6486 4922 6510 4924
rect 6566 4922 6590 4924
rect 6646 4922 6670 4924
rect 6726 4922 6732 4924
rect 6486 4870 6488 4922
rect 6668 4870 6670 4922
rect 6424 4868 6430 4870
rect 6486 4868 6510 4870
rect 6566 4868 6590 4870
rect 6646 4868 6670 4870
rect 6726 4868 6732 4870
rect 6424 4859 6732 4868
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6424 3836 6732 3845
rect 6424 3834 6430 3836
rect 6486 3834 6510 3836
rect 6566 3834 6590 3836
rect 6646 3834 6670 3836
rect 6726 3834 6732 3836
rect 6486 3782 6488 3834
rect 6668 3782 6670 3834
rect 6424 3780 6430 3782
rect 6486 3780 6510 3782
rect 6566 3780 6590 3782
rect 6646 3780 6670 3782
rect 6726 3780 6732 3782
rect 6424 3771 6732 3780
rect 1584 3528 1636 3534
rect 1582 3496 1584 3505
rect 1636 3496 1638 3505
rect 1582 3431 1638 3440
rect 6840 3058 6868 8298
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7024 6866 7052 7822
rect 7392 7478 7420 9862
rect 8220 9586 8248 10406
rect 8312 10130 8340 11086
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8496 9994 8524 11222
rect 8956 11150 8984 11630
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8956 10470 8984 11086
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 9048 10266 9076 11018
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 9110 8248 9318
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7472 8900 7524 8906
rect 7472 8842 7524 8848
rect 7484 8430 7512 8842
rect 7668 8634 7696 8910
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7852 8090 7880 8910
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8498 8800 8774
rect 9232 8498 9260 10406
rect 9416 10062 9444 12038
rect 9600 11082 9628 12242
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 9876 11898 9904 12038
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 10244 11694 10272 12038
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10336 11354 10364 12106
rect 10520 11694 10548 12786
rect 10612 11830 10640 13126
rect 10704 12850 10732 16662
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 11164 13326 11192 13738
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9600 10606 9628 11018
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 10244 10538 10272 10950
rect 10336 10742 10364 11290
rect 10428 11082 10456 11290
rect 10520 11150 10548 11630
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10704 10962 10732 12786
rect 10796 12238 10824 13194
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10520 10934 10732 10962
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9508 9586 9536 10066
rect 10428 9994 10456 10542
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9324 8498 9352 9318
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 8588 7818 8616 8230
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 9508 7478 9536 9522
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9692 7886 9720 8910
rect 10428 8906 10456 9930
rect 10520 9042 10548 10934
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10612 8634 10640 10746
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10704 10198 10732 10610
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10888 9058 10916 12582
rect 11532 12170 11560 13126
rect 11520 12164 11572 12170
rect 11520 12106 11572 12112
rect 11716 11762 11744 16730
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 11898 16348 12206 16357
rect 11898 16346 11904 16348
rect 11960 16346 11984 16348
rect 12040 16346 12064 16348
rect 12120 16346 12144 16348
rect 12200 16346 12206 16348
rect 11960 16294 11962 16346
rect 12142 16294 12144 16346
rect 11898 16292 11904 16294
rect 11960 16292 11984 16294
rect 12040 16292 12064 16294
rect 12120 16292 12144 16294
rect 12200 16292 12206 16294
rect 11898 16283 12206 16292
rect 11898 15260 12206 15269
rect 11898 15258 11904 15260
rect 11960 15258 11984 15260
rect 12040 15258 12064 15260
rect 12120 15258 12144 15260
rect 12200 15258 12206 15260
rect 11960 15206 11962 15258
rect 12142 15206 12144 15258
rect 11898 15204 11904 15206
rect 11960 15204 11984 15206
rect 12040 15204 12064 15206
rect 12120 15204 12144 15206
rect 12200 15204 12206 15206
rect 11898 15195 12206 15204
rect 12256 15020 12308 15026
rect 12900 15020 12952 15026
rect 12256 14962 12308 14968
rect 12728 14980 12900 15008
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11808 13410 11836 14758
rect 11898 14172 12206 14181
rect 11898 14170 11904 14172
rect 11960 14170 11984 14172
rect 12040 14170 12064 14172
rect 12120 14170 12144 14172
rect 12200 14170 12206 14172
rect 11960 14118 11962 14170
rect 12142 14118 12144 14170
rect 11898 14116 11904 14118
rect 11960 14116 11984 14118
rect 12040 14116 12064 14118
rect 12120 14116 12144 14118
rect 12200 14116 12206 14118
rect 11898 14107 12206 14116
rect 12268 14074 12296 14962
rect 12728 14482 12756 14980
rect 12900 14962 12952 14968
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12360 13734 12388 14214
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 11808 13382 11928 13410
rect 11900 13326 11928 13382
rect 12544 13326 12572 14418
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12636 13938 12664 14282
rect 12728 14074 12756 14418
rect 13096 14414 13124 14962
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13280 14414 13308 14758
rect 13556 14414 13584 14758
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12820 13938 12848 14214
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12912 13190 12940 14350
rect 13096 14074 13124 14350
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 13004 13462 13032 14010
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 11898 13084 12206 13093
rect 11898 13082 11904 13084
rect 11960 13082 11984 13084
rect 12040 13082 12064 13084
rect 12120 13082 12144 13084
rect 12200 13082 12206 13084
rect 11960 13030 11962 13082
rect 12142 13030 12144 13082
rect 11898 13028 11904 13030
rect 11960 13028 11984 13030
rect 12040 13028 12064 13030
rect 12120 13028 12144 13030
rect 12200 13028 12206 13030
rect 11898 13019 12206 13028
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12072 12436 12124 12442
rect 12176 12434 12204 12582
rect 12256 12436 12308 12442
rect 12176 12406 12256 12434
rect 12072 12378 12124 12384
rect 12256 12378 12308 12384
rect 12084 12209 12112 12378
rect 12070 12200 12126 12209
rect 12070 12135 12126 12144
rect 11898 11996 12206 12005
rect 11898 11994 11904 11996
rect 11960 11994 11984 11996
rect 12040 11994 12064 11996
rect 12120 11994 12144 11996
rect 12200 11994 12206 11996
rect 11960 11942 11962 11994
rect 12142 11942 12144 11994
rect 11898 11940 11904 11942
rect 11960 11940 11984 11942
rect 12040 11940 12064 11942
rect 12120 11940 12144 11942
rect 12200 11940 12206 11942
rect 11898 11931 12206 11940
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 11704 11620 11756 11626
rect 11704 11562 11756 11568
rect 11716 11218 11744 11562
rect 12084 11558 12112 11698
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12176 11286 12204 11698
rect 12164 11280 12216 11286
rect 12164 11222 12216 11228
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 12268 11150 12296 12378
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12360 12102 12388 12310
rect 12544 12306 12572 12854
rect 14476 12850 14504 13330
rect 15028 13190 15056 14010
rect 15488 14006 15516 14350
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15580 14006 15608 14282
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12544 11830 12572 12242
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11072 9654 11100 10202
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10796 9030 10916 9058
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7024 6390 7052 6802
rect 9876 6798 9904 8570
rect 10796 8294 10824 9030
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 7478 10824 8230
rect 10888 8090 10916 8842
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10784 7472 10836 7478
rect 10784 7414 10836 7420
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 8220 6458 8248 6666
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 7024 5710 7052 6326
rect 8956 6186 8984 6666
rect 9048 6322 9076 6666
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8956 5778 8984 6122
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 9140 5710 9168 6598
rect 7012 5704 7064 5710
rect 9128 5704 9180 5710
rect 7012 5646 7064 5652
rect 8206 5672 8262 5681
rect 7024 5234 7052 5646
rect 9128 5646 9180 5652
rect 8206 5607 8208 5616
rect 8260 5607 8262 5616
rect 8208 5578 8260 5584
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 5302 8984 5510
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9140 4690 9168 4966
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 20 2508 72 2514
rect 20 2450 72 2456
rect 32 800 60 2450
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 1320 800 1348 2382
rect 1596 1465 1624 2790
rect 6288 2446 6316 2790
rect 6424 2748 6732 2757
rect 6424 2746 6430 2748
rect 6486 2746 6510 2748
rect 6566 2746 6590 2748
rect 6646 2746 6670 2748
rect 6726 2746 6732 2748
rect 6486 2694 6488 2746
rect 6668 2694 6670 2746
rect 6424 2692 6430 2694
rect 6486 2692 6510 2694
rect 6566 2692 6590 2694
rect 6646 2692 6670 2694
rect 6726 2692 6732 2694
rect 6424 2683 6732 2692
rect 9692 2446 9720 6734
rect 9876 5166 9904 6734
rect 10060 5914 10088 6734
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10336 6458 10364 6666
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10796 6390 10824 6734
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10704 5370 10732 6054
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10796 5234 10824 6054
rect 11072 5846 11100 7754
rect 11256 7290 11284 11018
rect 11898 10908 12206 10917
rect 11898 10906 11904 10908
rect 11960 10906 11984 10908
rect 12040 10906 12064 10908
rect 12120 10906 12144 10908
rect 12200 10906 12206 10908
rect 11960 10854 11962 10906
rect 12142 10854 12144 10906
rect 11898 10852 11904 10854
rect 11960 10852 11984 10854
rect 12040 10852 12064 10854
rect 12120 10852 12144 10854
rect 12200 10852 12206 10854
rect 11898 10843 12206 10852
rect 12360 10266 12388 11630
rect 12636 11354 12664 12038
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12452 11014 12480 11222
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12440 10192 12492 10198
rect 12440 10134 12492 10140
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11348 9382 11376 9998
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 11898 9820 12206 9829
rect 11898 9818 11904 9820
rect 11960 9818 11984 9820
rect 12040 9818 12064 9820
rect 12120 9818 12144 9820
rect 12200 9818 12206 9820
rect 11960 9766 11962 9818
rect 12142 9766 12144 9818
rect 11898 9764 11904 9766
rect 11960 9764 11984 9766
rect 12040 9764 12064 9766
rect 12120 9764 12144 9766
rect 12200 9764 12206 9766
rect 11898 9755 12206 9764
rect 12268 9722 12296 9862
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12360 9586 12388 10066
rect 12452 9926 12480 10134
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11532 7886 11560 9318
rect 12452 9178 12480 9590
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11716 8498 11744 8910
rect 11898 8732 12206 8741
rect 11898 8730 11904 8732
rect 11960 8730 11984 8732
rect 12040 8730 12064 8732
rect 12120 8730 12144 8732
rect 12200 8730 12206 8732
rect 11960 8678 11962 8730
rect 12142 8678 12144 8730
rect 11898 8676 11904 8678
rect 11960 8676 11984 8678
rect 12040 8676 12064 8678
rect 12120 8676 12144 8678
rect 12200 8676 12206 8678
rect 11898 8667 12206 8676
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11716 7954 11744 8434
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11716 7478 11744 7686
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11256 7262 11376 7290
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 11164 5098 11192 6190
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 3534 11192 4422
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11256 3058 11284 7142
rect 11348 6322 11376 7262
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11348 6118 11376 6258
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11624 5914 11652 6326
rect 11716 6322 11744 7142
rect 11808 6458 11836 8434
rect 11898 7644 12206 7653
rect 11898 7642 11904 7644
rect 11960 7642 11984 7644
rect 12040 7642 12064 7644
rect 12120 7642 12144 7644
rect 12200 7642 12206 7644
rect 11960 7590 11962 7642
rect 12142 7590 12144 7642
rect 11898 7588 11904 7590
rect 11960 7588 11984 7590
rect 12040 7588 12064 7590
rect 12120 7588 12144 7590
rect 12200 7588 12206 7590
rect 11898 7579 12206 7588
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12360 6934 12388 7278
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 11898 6556 12206 6565
rect 11898 6554 11904 6556
rect 11960 6554 11984 6556
rect 12040 6554 12064 6556
rect 12120 6554 12144 6556
rect 12200 6554 12206 6556
rect 11960 6502 11962 6554
rect 12142 6502 12144 6554
rect 11898 6500 11904 6502
rect 11960 6500 11984 6502
rect 12040 6500 12064 6502
rect 12120 6500 12144 6502
rect 12200 6500 12206 6502
rect 11898 6491 12206 6500
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11808 5914 11836 6054
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11348 5302 11376 5782
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11624 4690 11652 5850
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11808 5370 11836 5578
rect 11898 5468 12206 5477
rect 11898 5466 11904 5468
rect 11960 5466 11984 5468
rect 12040 5466 12064 5468
rect 12120 5466 12144 5468
rect 12200 5466 12206 5468
rect 11960 5414 11962 5466
rect 12142 5414 12144 5466
rect 11898 5412 11904 5414
rect 11960 5412 11984 5414
rect 12040 5412 12064 5414
rect 12120 5412 12144 5414
rect 12200 5412 12206 5414
rect 11898 5403 12206 5412
rect 12268 5370 12296 6598
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12360 5166 12388 6870
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11440 3670 11468 4558
rect 11624 4146 11652 4626
rect 11716 4486 11744 4762
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 12360 4706 12388 4762
rect 12544 4706 12572 11086
rect 12636 11014 12664 11290
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11808 4214 11836 4694
rect 12360 4678 12572 4706
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 11898 4380 12206 4389
rect 11898 4378 11904 4380
rect 11960 4378 11984 4380
rect 12040 4378 12064 4380
rect 12120 4378 12144 4380
rect 12200 4378 12206 4380
rect 11960 4326 11962 4378
rect 12142 4326 12144 4378
rect 11898 4324 11904 4326
rect 11960 4324 11984 4326
rect 12040 4324 12064 4326
rect 12120 4324 12144 4326
rect 12200 4324 12206 4326
rect 11898 4315 12206 4324
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 12452 3738 12480 4490
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 12544 3534 12572 3878
rect 12636 3602 12664 5850
rect 12728 5681 12756 11494
rect 13004 11354 13032 12786
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13096 10266 13124 12174
rect 13372 10742 13400 12582
rect 13728 12368 13780 12374
rect 13556 12328 13728 12356
rect 13556 12238 13584 12328
rect 13728 12310 13780 12316
rect 13924 12238 13952 12786
rect 14660 12442 14688 12786
rect 15028 12764 15056 13126
rect 15304 12918 15332 13262
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15292 12776 15344 12782
rect 15028 12736 15292 12764
rect 15292 12718 15344 12724
rect 15488 12442 15516 13262
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 13450 11792 13506 11801
rect 13450 11727 13506 11736
rect 13464 11626 13492 11727
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 13464 11218 13492 11562
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 14108 11150 14136 11494
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 14016 10690 14044 11018
rect 14200 10810 14228 11154
rect 14844 10810 14872 12174
rect 15474 11792 15530 11801
rect 15474 11727 15530 11736
rect 15488 11694 15516 11727
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14292 10690 14320 10746
rect 14016 10662 14320 10690
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14568 10266 14596 10542
rect 15028 10266 15056 10678
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 12900 10056 12952 10062
rect 14280 10056 14332 10062
rect 12900 9998 12952 10004
rect 14278 10024 14280 10033
rect 14332 10024 14334 10033
rect 12912 9654 12940 9998
rect 14278 9959 14334 9968
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 13004 9586 13032 9862
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13004 9178 13032 9522
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12820 7546 12848 8774
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 13004 5710 13032 9114
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13096 8634 13124 8910
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13280 7750 13308 8774
rect 13556 8634 13584 9522
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13372 8090 13400 8230
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13372 7410 13400 7822
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13464 6866 13492 8230
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13188 5710 13216 6054
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 12992 5704 13044 5710
rect 12714 5672 12770 5681
rect 12992 5646 13044 5652
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 12714 5607 12770 5616
rect 12728 5574 12756 5607
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 13004 5302 13032 5646
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 13464 5098 13492 5714
rect 13648 5370 13676 9862
rect 14292 9674 14320 9959
rect 14200 9646 14320 9674
rect 14200 8430 14228 9646
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14660 9042 14688 9318
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14752 8498 14780 8978
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14752 7886 14780 8434
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 14108 4826 14136 7346
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14292 4622 14320 6598
rect 14648 6316 14700 6322
rect 14752 6304 14780 6734
rect 15212 6390 15240 11562
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15488 10810 15516 11018
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15304 9926 15332 10610
rect 15672 10554 15700 16526
rect 16776 16454 16804 17138
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 32588 17128 32640 17134
rect 32588 17070 32640 17076
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16868 16794 16896 16934
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16868 15722 16896 16730
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 16776 15694 16896 15722
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15764 14346 15792 14758
rect 15752 14340 15804 14346
rect 15752 14282 15804 14288
rect 16132 14074 16160 14962
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15856 12238 15884 12582
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15948 11762 15976 12854
rect 16040 12306 16068 13398
rect 16316 13326 16344 13806
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16212 13252 16264 13258
rect 16212 13194 16264 13200
rect 16224 12850 16252 13194
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16316 12782 16344 13262
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15764 11218 15792 11630
rect 15948 11354 15976 11698
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15488 10526 15700 10554
rect 15488 10470 15516 10526
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15580 8906 15608 10406
rect 15764 10130 15792 11154
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 15856 10810 15884 10950
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15764 9722 15792 10066
rect 16040 9994 16068 10950
rect 16028 9988 16080 9994
rect 16028 9930 16080 9936
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 16408 9518 16436 13738
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16500 12374 16528 13126
rect 16684 12850 16712 14350
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 16684 11694 16712 12786
rect 16776 12238 16804 15694
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16868 13938 16896 14214
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16868 12238 16896 13670
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16592 11014 16620 11222
rect 16684 11150 16712 11494
rect 16868 11286 16896 12174
rect 17052 11898 17080 12718
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16684 9586 16712 9862
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15304 8498 15332 8842
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15396 7546 15424 7822
rect 15488 7546 15516 8774
rect 15856 8634 15884 9454
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15580 8090 15608 8434
rect 15948 8090 15976 9454
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16500 8566 16528 9318
rect 16684 8974 16712 9318
rect 17052 9110 17080 9454
rect 17144 9450 17172 16526
rect 17236 12434 17264 17070
rect 17372 16892 17680 16901
rect 17372 16890 17378 16892
rect 17434 16890 17458 16892
rect 17514 16890 17538 16892
rect 17594 16890 17618 16892
rect 17674 16890 17680 16892
rect 17434 16838 17436 16890
rect 17616 16838 17618 16890
rect 17372 16836 17378 16838
rect 17434 16836 17458 16838
rect 17514 16836 17538 16838
rect 17594 16836 17618 16838
rect 17674 16836 17680 16838
rect 17372 16827 17680 16836
rect 17972 16454 18000 17070
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 22846 16348 23154 16357
rect 22846 16346 22852 16348
rect 22908 16346 22932 16348
rect 22988 16346 23012 16348
rect 23068 16346 23092 16348
rect 23148 16346 23154 16348
rect 22908 16294 22910 16346
rect 23090 16294 23092 16346
rect 22846 16292 22852 16294
rect 22908 16292 22932 16294
rect 22988 16292 23012 16294
rect 23068 16292 23092 16294
rect 23148 16292 23154 16294
rect 22846 16283 23154 16292
rect 17372 15804 17680 15813
rect 17372 15802 17378 15804
rect 17434 15802 17458 15804
rect 17514 15802 17538 15804
rect 17594 15802 17618 15804
rect 17674 15802 17680 15804
rect 17434 15750 17436 15802
rect 17616 15750 17618 15802
rect 17372 15748 17378 15750
rect 17434 15748 17458 15750
rect 17514 15748 17538 15750
rect 17594 15748 17618 15750
rect 17674 15748 17680 15750
rect 17372 15739 17680 15748
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 18064 15094 18092 15302
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 18616 14890 18644 15438
rect 19168 15366 19196 15438
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19432 15428 19484 15434
rect 19432 15370 19484 15376
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19168 15162 19196 15302
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 18604 14884 18656 14890
rect 18604 14826 18656 14832
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 17372 14716 17680 14725
rect 17372 14714 17378 14716
rect 17434 14714 17458 14716
rect 17514 14714 17538 14716
rect 17594 14714 17618 14716
rect 17674 14714 17680 14716
rect 17434 14662 17436 14714
rect 17616 14662 17618 14714
rect 17372 14660 17378 14662
rect 17434 14660 17458 14662
rect 17514 14660 17538 14662
rect 17594 14660 17618 14662
rect 17674 14660 17680 14662
rect 17372 14651 17680 14660
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17604 14074 17632 14282
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 18432 13734 18460 14758
rect 18616 14278 18644 14826
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18708 14006 18736 15098
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18800 14278 18828 14962
rect 19168 14550 19196 15098
rect 19260 15094 19288 15370
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19156 14544 19208 14550
rect 19156 14486 19208 14492
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 17372 13628 17680 13637
rect 17372 13626 17378 13628
rect 17434 13626 17458 13628
rect 17514 13626 17538 13628
rect 17594 13626 17618 13628
rect 17674 13626 17680 13628
rect 17434 13574 17436 13626
rect 17616 13574 17618 13626
rect 17372 13572 17378 13574
rect 17434 13572 17458 13574
rect 17514 13572 17538 13574
rect 17594 13572 17618 13574
rect 17674 13572 17680 13574
rect 17372 13563 17680 13572
rect 18524 13462 18552 13942
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18616 13734 18644 13874
rect 18604 13728 18656 13734
rect 18604 13670 18656 13676
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18800 13394 18828 14214
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 19168 13326 19196 14486
rect 19260 14414 19288 15030
rect 19444 14958 19472 15370
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19352 13938 19380 14758
rect 19444 14498 19472 14894
rect 19536 14618 19564 15302
rect 22846 15260 23154 15269
rect 22846 15258 22852 15260
rect 22908 15258 22932 15260
rect 22988 15258 23012 15260
rect 23068 15258 23092 15260
rect 23148 15258 23154 15260
rect 22908 15206 22910 15258
rect 23090 15206 23092 15258
rect 22846 15204 22852 15206
rect 22908 15204 22932 15206
rect 22988 15204 23012 15206
rect 23068 15204 23092 15206
rect 23148 15204 23154 15206
rect 22846 15195 23154 15204
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19444 14470 19656 14498
rect 19812 14482 19840 14962
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19444 13462 19472 14470
rect 19628 14414 19656 14470
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 19800 14340 19852 14346
rect 19800 14282 19852 14288
rect 19812 14074 19840 14282
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19996 13734 20024 14214
rect 20180 14074 20208 14350
rect 20548 14346 20576 14758
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 21284 13938 21312 14214
rect 21376 14006 21404 14214
rect 22846 14172 23154 14181
rect 22846 14170 22852 14172
rect 22908 14170 22932 14172
rect 22988 14170 23012 14172
rect 23068 14170 23092 14172
rect 23148 14170 23154 14172
rect 22908 14118 22910 14170
rect 23090 14118 23092 14170
rect 22846 14116 22852 14118
rect 22908 14116 22932 14118
rect 22988 14116 23012 14118
rect 23068 14116 23092 14118
rect 23148 14116 23154 14118
rect 22846 14107 23154 14116
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19432 13456 19484 13462
rect 19352 13416 19432 13444
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 17776 12912 17828 12918
rect 17776 12854 17828 12860
rect 17372 12540 17680 12549
rect 17372 12538 17378 12540
rect 17434 12538 17458 12540
rect 17514 12538 17538 12540
rect 17594 12538 17618 12540
rect 17674 12538 17680 12540
rect 17434 12486 17436 12538
rect 17616 12486 17618 12538
rect 17372 12484 17378 12486
rect 17434 12484 17458 12486
rect 17514 12484 17538 12486
rect 17594 12484 17618 12486
rect 17674 12484 17680 12486
rect 17372 12475 17680 12484
rect 17236 12406 17632 12434
rect 17604 12102 17632 12406
rect 17788 12374 17816 12854
rect 17880 12850 17908 13262
rect 19352 13258 19380 13416
rect 19432 13398 19484 13404
rect 20260 13456 20312 13462
rect 20260 13398 20312 13404
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17880 12238 17908 12786
rect 18432 12238 18460 13194
rect 20272 12782 20300 13398
rect 20640 13394 20668 13806
rect 22204 13518 22784 13546
rect 20996 13456 21048 13462
rect 20996 13398 21048 13404
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 17868 12232 17920 12238
rect 18420 12232 18472 12238
rect 17868 12174 17920 12180
rect 18326 12200 18382 12209
rect 18420 12174 18472 12180
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 18326 12135 18382 12144
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17236 11762 17264 12038
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17372 11452 17680 11461
rect 17372 11450 17378 11452
rect 17434 11450 17458 11452
rect 17514 11450 17538 11452
rect 17594 11450 17618 11452
rect 17674 11450 17680 11452
rect 17434 11398 17436 11450
rect 17616 11398 17618 11450
rect 17372 11396 17378 11398
rect 17434 11396 17458 11398
rect 17514 11396 17538 11398
rect 17594 11396 17618 11398
rect 17674 11396 17680 11398
rect 17372 11387 17680 11396
rect 17880 11218 17908 11630
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17372 10364 17680 10373
rect 17372 10362 17378 10364
rect 17434 10362 17458 10364
rect 17514 10362 17538 10364
rect 17594 10362 17618 10364
rect 17674 10362 17680 10364
rect 17434 10310 17436 10362
rect 17616 10310 17618 10362
rect 17372 10308 17378 10310
rect 17434 10308 17458 10310
rect 17514 10308 17538 10310
rect 17594 10308 17618 10310
rect 17674 10308 17680 10310
rect 17372 10299 17680 10308
rect 17788 9994 17816 10406
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17132 9444 17184 9450
rect 17132 9386 17184 9392
rect 17372 9276 17680 9285
rect 17372 9274 17378 9276
rect 17434 9274 17458 9276
rect 17514 9274 17538 9276
rect 17594 9274 17618 9276
rect 17674 9274 17680 9276
rect 17434 9222 17436 9274
rect 17616 9222 17618 9274
rect 17372 9220 17378 9222
rect 17434 9220 17458 9222
rect 17514 9220 17538 9222
rect 17594 9220 17618 9222
rect 17674 9220 17680 9222
rect 17372 9211 17680 9220
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 16500 8022 16528 8502
rect 17972 8498 18000 12038
rect 18064 11150 18092 12038
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18248 11694 18276 11766
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18156 11354 18184 11630
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18340 11082 18368 12135
rect 19168 11898 19196 12174
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 18604 11824 18656 11830
rect 18604 11766 18656 11772
rect 19246 11792 19302 11801
rect 18616 11354 18644 11766
rect 19720 11778 19748 11834
rect 19302 11750 19748 11778
rect 19246 11727 19302 11736
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18524 10606 18552 11086
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18694 10024 18750 10033
rect 18340 9926 18368 9998
rect 18694 9959 18750 9968
rect 18708 9926 18736 9959
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 18524 9654 18552 9862
rect 19352 9654 19380 10950
rect 19720 10266 19748 11018
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18512 9648 18564 9654
rect 18512 9590 18564 9596
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 18064 8974 18092 9590
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17372 8188 17680 8197
rect 17372 8186 17378 8188
rect 17434 8186 17458 8188
rect 17514 8186 17538 8188
rect 17594 8186 17618 8188
rect 17674 8186 17680 8188
rect 17434 8134 17436 8186
rect 17616 8134 17618 8186
rect 17372 8132 17378 8134
rect 17434 8132 17458 8134
rect 17514 8132 17538 8134
rect 17594 8132 17618 8134
rect 17674 8132 17680 8134
rect 17372 8123 17680 8132
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15672 7002 15700 7278
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 14700 6276 14780 6304
rect 14648 6258 14700 6264
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 12728 4146 12756 4558
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12728 3602 12756 4082
rect 14568 4078 14596 5578
rect 14752 5166 14780 6276
rect 15212 5658 15240 6326
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5710 15608 6054
rect 15764 5914 15792 6734
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15120 5630 15240 5658
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14752 4690 14780 5102
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14844 4282 14872 5170
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 15028 4622 15056 4966
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 15120 4570 15148 5630
rect 16040 5302 16068 7958
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16684 7274 16712 7822
rect 17512 7342 17540 7890
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16868 6866 16896 7142
rect 17372 7100 17680 7109
rect 17372 7098 17378 7100
rect 17434 7098 17458 7100
rect 17514 7098 17538 7100
rect 17594 7098 17618 7100
rect 17674 7098 17680 7100
rect 17434 7046 17436 7098
rect 17616 7046 17618 7098
rect 17372 7044 17378 7046
rect 17434 7044 17458 7046
rect 17514 7044 17538 7046
rect 17594 7044 17618 7046
rect 17674 7044 17680 7046
rect 17372 7035 17680 7044
rect 16856 6860 16908 6866
rect 16856 6802 16908 6808
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16776 5846 16804 6122
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16764 5840 16816 5846
rect 16764 5782 16816 5788
rect 16868 5642 16896 6054
rect 16960 5846 16988 6802
rect 17972 6458 18000 8434
rect 18064 8430 18092 8910
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 18064 7342 18092 8366
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18708 7886 18736 8026
rect 19260 7886 19288 8910
rect 19444 8634 19472 9522
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19720 9042 19748 9318
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19260 7478 19288 7822
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 7546 19380 7686
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17372 6012 17680 6021
rect 17372 6010 17378 6012
rect 17434 6010 17458 6012
rect 17514 6010 17538 6012
rect 17594 6010 17618 6012
rect 17674 6010 17680 6012
rect 17434 5958 17436 6010
rect 17616 5958 17618 6010
rect 17372 5956 17378 5958
rect 17434 5956 17458 5958
rect 17514 5956 17538 5958
rect 17594 5956 17618 5958
rect 17674 5956 17680 5958
rect 17372 5947 17680 5956
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 18064 5710 18092 7278
rect 18340 7002 18368 7346
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18708 7002 18736 7142
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18340 5914 18368 6258
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 17512 5234 17540 5646
rect 19812 5370 19840 12038
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 20088 11558 20116 11630
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20088 11354 20116 11494
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19904 11014 19932 11086
rect 19892 11008 19944 11014
rect 19892 10950 19944 10956
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19904 9722 19932 9998
rect 19892 9716 19944 9722
rect 19892 9658 19944 9664
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 19904 8090 19932 8230
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 20272 7426 20300 12718
rect 20444 12368 20496 12374
rect 20444 12310 20496 12316
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20364 11762 20392 12242
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20364 11354 20392 11698
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20456 11218 20484 12310
rect 20640 12238 20668 13330
rect 21008 12782 21036 13398
rect 22204 13394 22232 13518
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22284 13388 22336 13394
rect 22284 13330 22336 13336
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20916 12306 20944 12582
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20640 11014 20668 12174
rect 21100 11898 21128 12718
rect 21376 12714 21404 13262
rect 22296 12986 22324 13330
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22388 12986 22416 13126
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 22480 12866 22508 13518
rect 22756 13462 22784 13518
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22744 13252 22796 13258
rect 22744 13194 22796 13200
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22388 12838 22508 12866
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 22112 12442 22140 12718
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21284 11898 21312 12106
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20640 10130 20668 10950
rect 21008 10674 21036 11630
rect 22020 11558 22048 11698
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 21916 10736 21968 10742
rect 22020 10713 22048 10746
rect 21916 10678 21968 10684
rect 22006 10704 22062 10713
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 21008 10146 21036 10610
rect 21928 10538 21956 10678
rect 22006 10639 22062 10648
rect 21732 10532 21784 10538
rect 21732 10474 21784 10480
rect 21916 10532 21968 10538
rect 21916 10474 21968 10480
rect 20628 10124 20680 10130
rect 21008 10118 21220 10146
rect 21744 10130 21772 10474
rect 20628 10066 20680 10072
rect 21192 10062 21220 10118
rect 21732 10124 21784 10130
rect 21732 10066 21784 10072
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20640 9518 20668 9590
rect 22020 9518 22048 9998
rect 22112 9926 22140 11154
rect 22296 11082 22324 12582
rect 22388 11150 22416 12838
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22480 12306 22508 12718
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 22388 10810 22416 10950
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22284 10600 22336 10606
rect 22468 10600 22520 10606
rect 22284 10542 22336 10548
rect 22388 10560 22468 10588
rect 22296 10266 22324 10542
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 20640 9058 20668 9454
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 21192 9110 21220 9386
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21180 9104 21232 9110
rect 20640 9042 20760 9058
rect 21180 9046 21232 9052
rect 20640 9036 20772 9042
rect 20640 9030 20720 9036
rect 20720 8978 20772 8984
rect 21284 8498 21312 9318
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20364 7546 20392 8366
rect 20456 8294 20484 8366
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20456 7857 20484 8230
rect 21100 8090 21128 8434
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 20442 7848 20498 7857
rect 20442 7783 20498 7792
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20180 7410 20300 7426
rect 20168 7404 20300 7410
rect 20220 7398 20300 7404
rect 20168 7346 20220 7352
rect 20272 6934 20300 7398
rect 21364 7268 21416 7274
rect 21364 7210 21416 7216
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20260 6928 20312 6934
rect 20260 6870 20312 6876
rect 20824 6798 20852 7142
rect 21376 6866 21404 7210
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 20732 6322 20760 6598
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 19892 6180 19944 6186
rect 19892 6122 19944 6128
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19800 5364 19852 5370
rect 19800 5306 19852 5312
rect 17776 5296 17828 5302
rect 17776 5238 17828 5244
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15120 4542 15240 4570
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15120 4282 15148 4422
rect 15212 4282 15240 4542
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 15212 4162 15240 4218
rect 15120 4134 15240 4162
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 11898 3292 12206 3301
rect 11898 3290 11904 3292
rect 11960 3290 11984 3292
rect 12040 3290 12064 3292
rect 12120 3290 12144 3292
rect 12200 3290 12206 3292
rect 11960 3238 11962 3290
rect 12142 3238 12144 3290
rect 11898 3236 11904 3238
rect 11960 3236 11984 3238
rect 12040 3236 12064 3238
rect 12120 3236 12144 3238
rect 12200 3236 12206 3238
rect 11898 3227 12206 3236
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 13004 2650 13032 3470
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 14476 2446 14504 2790
rect 15120 2582 15148 4134
rect 15764 3534 15792 5102
rect 17236 4146 17264 5170
rect 17372 4924 17680 4933
rect 17372 4922 17378 4924
rect 17434 4922 17458 4924
rect 17514 4922 17538 4924
rect 17594 4922 17618 4924
rect 17674 4922 17680 4924
rect 17434 4870 17436 4922
rect 17616 4870 17618 4922
rect 17372 4868 17378 4870
rect 17434 4868 17458 4870
rect 17514 4868 17538 4870
rect 17594 4868 17618 4870
rect 17674 4868 17680 4870
rect 17372 4859 17680 4868
rect 17788 4826 17816 5238
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 18064 4622 18092 4966
rect 19352 4690 19380 5306
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 18156 4078 18184 4422
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 16776 3602 16804 3878
rect 17372 3836 17680 3845
rect 17372 3834 17378 3836
rect 17434 3834 17458 3836
rect 17514 3834 17538 3836
rect 17594 3834 17618 3836
rect 17674 3834 17680 3836
rect 17434 3782 17436 3834
rect 17616 3782 17618 3834
rect 17372 3780 17378 3782
rect 17434 3780 17458 3782
rect 17514 3780 17538 3782
rect 17594 3780 17618 3782
rect 17674 3780 17680 3782
rect 17372 3771 17680 3780
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 17144 3194 17172 3402
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17788 3058 17816 3878
rect 18248 3738 18276 4082
rect 19444 4078 19472 4966
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 19260 3602 19288 3878
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 18156 3058 18184 3334
rect 19628 3194 19656 3470
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 17776 2916 17828 2922
rect 17776 2858 17828 2864
rect 17372 2748 17680 2757
rect 17372 2746 17378 2748
rect 17434 2746 17458 2748
rect 17514 2746 17538 2748
rect 17594 2746 17618 2748
rect 17674 2746 17680 2748
rect 17434 2694 17436 2746
rect 17616 2694 17618 2746
rect 17372 2692 17378 2694
rect 17434 2692 17458 2694
rect 17514 2692 17538 2694
rect 17594 2692 17618 2694
rect 17674 2692 17680 2694
rect 17372 2683 17680 2692
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 17788 2514 17816 2858
rect 19812 2774 19840 5306
rect 19904 5166 19932 6122
rect 21100 6118 21128 6598
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 19892 5160 19944 5166
rect 19892 5102 19944 5108
rect 20456 4826 20484 5170
rect 20548 5166 20576 5714
rect 20626 5672 20682 5681
rect 20626 5607 20682 5616
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20640 4622 20668 5607
rect 21192 5574 21220 6394
rect 21376 6186 21404 6802
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 21364 6180 21416 6186
rect 21364 6122 21416 6128
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20732 4758 20760 5170
rect 21652 5098 21680 6190
rect 21744 5710 21772 9454
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21836 7478 21864 8366
rect 21824 7472 21876 7478
rect 21824 7414 21876 7420
rect 21836 6322 21864 7414
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 21640 5092 21692 5098
rect 21640 5034 21692 5040
rect 20720 4752 20772 4758
rect 20720 4694 20772 4700
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 21744 3534 21772 5646
rect 22112 4298 22140 8842
rect 22388 8566 22416 10560
rect 22572 10588 22600 12310
rect 22520 10560 22600 10588
rect 22468 10542 22520 10548
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22376 8560 22428 8566
rect 22376 8502 22428 8508
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22284 7880 22336 7886
rect 22284 7822 22336 7828
rect 22296 6730 22324 7822
rect 22388 7449 22416 7890
rect 22374 7440 22430 7449
rect 22374 7375 22430 7384
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22284 6724 22336 6730
rect 22284 6666 22336 6672
rect 22296 6610 22324 6666
rect 22388 6662 22416 7142
rect 22204 6582 22324 6610
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22204 4690 22232 6582
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 22020 4270 22140 4298
rect 22020 4026 22048 4270
rect 22020 3998 22140 4026
rect 22112 3602 22140 3998
rect 22204 3942 22232 4626
rect 22296 4214 22324 5102
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 20168 3460 20220 3466
rect 20168 3402 20220 3408
rect 20180 3194 20208 3402
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 22480 3058 22508 10406
rect 22664 7818 22692 13126
rect 22756 11898 22784 13194
rect 22846 13084 23154 13093
rect 22846 13082 22852 13084
rect 22908 13082 22932 13084
rect 22988 13082 23012 13084
rect 23068 13082 23092 13084
rect 23148 13082 23154 13084
rect 22908 13030 22910 13082
rect 23090 13030 23092 13082
rect 22846 13028 22852 13030
rect 22908 13028 22932 13030
rect 22988 13028 23012 13030
rect 23068 13028 23092 13030
rect 23148 13028 23154 13030
rect 22846 13019 23154 13028
rect 23020 12708 23072 12714
rect 23020 12650 23072 12656
rect 23032 12238 23060 12650
rect 23216 12442 23244 13806
rect 23308 13326 23336 14894
rect 23388 14884 23440 14890
rect 23388 14826 23440 14832
rect 23400 14074 23428 14826
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23308 12986 23336 13126
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23400 12850 23428 13874
rect 23480 13728 23532 13734
rect 23480 13670 23532 13676
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23492 12782 23520 13670
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23388 12708 23440 12714
rect 23388 12650 23440 12656
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 23400 12238 23428 12650
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 22846 11996 23154 12005
rect 22846 11994 22852 11996
rect 22908 11994 22932 11996
rect 22988 11994 23012 11996
rect 23068 11994 23092 11996
rect 23148 11994 23154 11996
rect 22908 11942 22910 11994
rect 23090 11942 23092 11994
rect 22846 11940 22852 11942
rect 22908 11940 22932 11942
rect 22988 11940 23012 11942
rect 23068 11940 23092 11942
rect 23148 11940 23154 11942
rect 22846 11931 23154 11940
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 23492 11762 23520 12038
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23492 11558 23520 11698
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23216 11218 23244 11290
rect 23308 11218 23336 11494
rect 23204 11212 23256 11218
rect 23204 11154 23256 11160
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23584 11150 23612 16934
rect 28320 16892 28628 16901
rect 28320 16890 28326 16892
rect 28382 16890 28406 16892
rect 28462 16890 28486 16892
rect 28542 16890 28566 16892
rect 28622 16890 28628 16892
rect 28382 16838 28384 16890
rect 28564 16838 28566 16890
rect 28320 16836 28326 16838
rect 28382 16836 28406 16838
rect 28462 16836 28486 16838
rect 28542 16836 28566 16838
rect 28622 16836 28628 16838
rect 28320 16827 28628 16836
rect 28320 15804 28628 15813
rect 28320 15802 28326 15804
rect 28382 15802 28406 15804
rect 28462 15802 28486 15804
rect 28542 15802 28566 15804
rect 28622 15802 28628 15804
rect 28382 15750 28384 15802
rect 28564 15750 28566 15802
rect 28320 15748 28326 15750
rect 28382 15748 28406 15750
rect 28462 15748 28486 15750
rect 28542 15748 28566 15750
rect 28622 15748 28628 15750
rect 28320 15739 28628 15748
rect 28320 14716 28628 14725
rect 28320 14714 28326 14716
rect 28382 14714 28406 14716
rect 28462 14714 28486 14716
rect 28542 14714 28566 14716
rect 28622 14714 28628 14716
rect 28382 14662 28384 14714
rect 28564 14662 28566 14714
rect 28320 14660 28326 14662
rect 28382 14660 28406 14662
rect 28462 14660 28486 14662
rect 28542 14660 28566 14662
rect 28622 14660 28628 14662
rect 28320 14651 28628 14660
rect 23940 14612 23992 14618
rect 23940 14554 23992 14560
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23860 12986 23888 14214
rect 23952 13870 23980 14554
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 24228 13326 24256 13874
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 24044 12238 24072 12922
rect 24216 12844 24268 12850
rect 24216 12786 24268 12792
rect 24228 12442 24256 12786
rect 24584 12708 24636 12714
rect 24584 12650 24636 12656
rect 24596 12442 24624 12650
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24584 12436 24636 12442
rect 24584 12378 24636 12384
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 24228 12102 24256 12378
rect 24492 12164 24544 12170
rect 24492 12106 24544 12112
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 24228 11830 24256 12038
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 24216 11824 24268 11830
rect 24216 11766 24268 11772
rect 23952 11694 23980 11766
rect 24504 11762 24532 12106
rect 24492 11756 24544 11762
rect 24492 11698 24544 11704
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 24596 11558 24624 12378
rect 24688 12374 24716 14350
rect 25412 13796 25464 13802
rect 25412 13738 25464 13744
rect 25424 13462 25452 13738
rect 28320 13628 28628 13637
rect 28320 13626 28326 13628
rect 28382 13626 28406 13628
rect 28462 13626 28486 13628
rect 28542 13626 28566 13628
rect 28622 13626 28628 13628
rect 28382 13574 28384 13626
rect 28564 13574 28566 13626
rect 28320 13572 28326 13574
rect 28382 13572 28406 13574
rect 28462 13572 28486 13574
rect 28542 13572 28566 13574
rect 28622 13572 28628 13574
rect 28320 13563 28628 13572
rect 25412 13456 25464 13462
rect 25412 13398 25464 13404
rect 32600 13394 32628 17070
rect 34152 16992 34204 16998
rect 34152 16934 34204 16940
rect 33692 16788 33744 16794
rect 33692 16730 33744 16736
rect 33704 14006 33732 16730
rect 33794 16348 34102 16357
rect 33794 16346 33800 16348
rect 33856 16346 33880 16348
rect 33936 16346 33960 16348
rect 34016 16346 34040 16348
rect 34096 16346 34102 16348
rect 33856 16294 33858 16346
rect 34038 16294 34040 16346
rect 33794 16292 33800 16294
rect 33856 16292 33880 16294
rect 33936 16292 33960 16294
rect 34016 16292 34040 16294
rect 34096 16292 34102 16294
rect 33794 16283 34102 16292
rect 33794 15260 34102 15269
rect 33794 15258 33800 15260
rect 33856 15258 33880 15260
rect 33936 15258 33960 15260
rect 34016 15258 34040 15260
rect 34096 15258 34102 15260
rect 33856 15206 33858 15258
rect 34038 15206 34040 15258
rect 33794 15204 33800 15206
rect 33856 15204 33880 15206
rect 33936 15204 33960 15206
rect 34016 15204 34040 15206
rect 34096 15204 34102 15206
rect 33794 15195 34102 15204
rect 33794 14172 34102 14181
rect 33794 14170 33800 14172
rect 33856 14170 33880 14172
rect 33936 14170 33960 14172
rect 34016 14170 34040 14172
rect 34096 14170 34102 14172
rect 33856 14118 33858 14170
rect 34038 14118 34040 14170
rect 33794 14116 33800 14118
rect 33856 14116 33880 14118
rect 33936 14116 33960 14118
rect 34016 14116 34040 14118
rect 34096 14116 34102 14118
rect 33794 14107 34102 14116
rect 33692 14000 33744 14006
rect 33692 13942 33744 13948
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 33244 13734 33272 13874
rect 33692 13796 33744 13802
rect 33692 13738 33744 13744
rect 33232 13728 33284 13734
rect 33232 13670 33284 13676
rect 32588 13388 32640 13394
rect 32588 13330 32640 13336
rect 26332 13320 26384 13326
rect 26332 13262 26384 13268
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 30288 13320 30340 13326
rect 30288 13262 30340 13268
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 33324 13320 33376 13326
rect 33324 13262 33376 13268
rect 25136 12912 25188 12918
rect 25136 12854 25188 12860
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 24676 12368 24728 12374
rect 24676 12310 24728 12316
rect 24688 11762 24716 12310
rect 25056 12102 25084 12582
rect 25148 12434 25176 12854
rect 25320 12776 25372 12782
rect 25320 12718 25372 12724
rect 25332 12442 25360 12718
rect 26344 12442 26372 13262
rect 26700 12708 26752 12714
rect 26700 12650 26752 12656
rect 26516 12640 26568 12646
rect 26516 12582 26568 12588
rect 25228 12436 25280 12442
rect 25148 12406 25228 12434
rect 25228 12378 25280 12384
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 26332 12436 26384 12442
rect 26332 12378 26384 12384
rect 25240 12306 25268 12378
rect 26240 12368 26292 12374
rect 26292 12316 26372 12322
rect 26240 12310 26372 12316
rect 25228 12300 25280 12306
rect 26252 12294 26372 12310
rect 26528 12306 26556 12582
rect 25228 12242 25280 12248
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 24676 11756 24728 11762
rect 24676 11698 24728 11704
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 22846 10908 23154 10917
rect 22846 10906 22852 10908
rect 22908 10906 22932 10908
rect 22988 10906 23012 10908
rect 23068 10906 23092 10908
rect 23148 10906 23154 10908
rect 22908 10854 22910 10906
rect 23090 10854 23092 10906
rect 22846 10852 22852 10854
rect 22908 10852 22932 10854
rect 22988 10852 23012 10854
rect 23068 10852 23092 10854
rect 23148 10852 23154 10854
rect 22846 10843 23154 10852
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 23032 10266 23060 10610
rect 23204 10464 23256 10470
rect 23204 10406 23256 10412
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 22846 9820 23154 9829
rect 22846 9818 22852 9820
rect 22908 9818 22932 9820
rect 22988 9818 23012 9820
rect 23068 9818 23092 9820
rect 23148 9818 23154 9820
rect 22908 9766 22910 9818
rect 23090 9766 23092 9818
rect 22846 9764 22852 9766
rect 22908 9764 22932 9766
rect 22988 9764 23012 9766
rect 23068 9764 23092 9766
rect 23148 9764 23154 9766
rect 22846 9755 23154 9764
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22664 7546 22692 7754
rect 22756 7546 22784 8774
rect 22846 8732 23154 8741
rect 22846 8730 22852 8732
rect 22908 8730 22932 8732
rect 22988 8730 23012 8732
rect 23068 8730 23092 8732
rect 23148 8730 23154 8732
rect 22908 8678 22910 8730
rect 23090 8678 23092 8730
rect 22846 8676 22852 8678
rect 22908 8676 22932 8678
rect 22988 8676 23012 8678
rect 23068 8676 23092 8678
rect 23148 8676 23154 8678
rect 22846 8667 23154 8676
rect 23216 8498 23244 10406
rect 23676 9654 23704 10950
rect 24688 10742 24716 11698
rect 24780 11150 24808 12038
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 24780 10742 24808 10950
rect 24676 10736 24728 10742
rect 24676 10678 24728 10684
rect 24768 10736 24820 10742
rect 24768 10678 24820 10684
rect 25148 9994 25176 11086
rect 25240 11014 25268 12242
rect 26344 11898 26372 12294
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 26332 11892 26384 11898
rect 26332 11834 26384 11840
rect 26436 11694 26464 12106
rect 26712 11762 26740 12650
rect 26804 12646 26832 13262
rect 27804 13252 27856 13258
rect 27804 13194 27856 13200
rect 27252 12776 27304 12782
rect 27252 12718 27304 12724
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 26804 11898 26832 12582
rect 27264 11898 27292 12718
rect 27816 12442 27844 13194
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 27988 12912 28040 12918
rect 27988 12854 28040 12860
rect 27804 12436 27856 12442
rect 27804 12378 27856 12384
rect 27436 12300 27488 12306
rect 27436 12242 27488 12248
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 27252 11892 27304 11898
rect 27252 11834 27304 11840
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 26148 11688 26200 11694
rect 26148 11630 26200 11636
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 25964 11620 26016 11626
rect 25964 11562 26016 11568
rect 25976 11354 26004 11562
rect 26160 11354 26188 11630
rect 26436 11370 26464 11630
rect 25964 11348 26016 11354
rect 25964 11290 26016 11296
rect 26148 11348 26200 11354
rect 26436 11342 26556 11370
rect 26148 11290 26200 11296
rect 26528 11218 26556 11342
rect 26516 11212 26568 11218
rect 26516 11154 26568 11160
rect 26976 11144 27028 11150
rect 26976 11086 27028 11092
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 25228 11008 25280 11014
rect 25228 10950 25280 10956
rect 26252 10810 26280 11018
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 25228 10736 25280 10742
rect 25228 10678 25280 10684
rect 25778 10704 25834 10713
rect 25240 10266 25268 10678
rect 25778 10639 25834 10648
rect 25792 10538 25820 10639
rect 25780 10532 25832 10538
rect 25780 10474 25832 10480
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 26988 10198 27016 11086
rect 27264 11014 27292 11698
rect 27344 11620 27396 11626
rect 27344 11562 27396 11568
rect 27252 11008 27304 11014
rect 27252 10950 27304 10956
rect 27264 10266 27292 10950
rect 27252 10260 27304 10266
rect 27252 10202 27304 10208
rect 26976 10192 27028 10198
rect 26976 10134 27028 10140
rect 26988 10062 27016 10134
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 26700 10056 26752 10062
rect 26700 9998 26752 10004
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 25136 9988 25188 9994
rect 25136 9930 25188 9936
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24964 9654 24992 9862
rect 25148 9722 25176 9930
rect 25240 9722 25268 9998
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 23664 9648 23716 9654
rect 23664 9590 23716 9596
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 25424 9586 25452 9998
rect 26332 9920 26384 9926
rect 26332 9862 26384 9868
rect 25412 9580 25464 9586
rect 25412 9522 25464 9528
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 26240 9512 26292 9518
rect 26240 9454 26292 9460
rect 23204 8492 23256 8498
rect 23204 8434 23256 8440
rect 23400 8090 23428 9454
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24492 8900 24544 8906
rect 24492 8842 24544 8848
rect 24504 8430 24532 8842
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 24504 7886 24532 8366
rect 24596 8090 24624 8910
rect 26252 8906 26280 9454
rect 26344 8906 26372 9862
rect 26240 8900 26292 8906
rect 26240 8842 26292 8848
rect 26332 8900 26384 8906
rect 26332 8842 26384 8848
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25056 8498 25084 8774
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 24584 8084 24636 8090
rect 24584 8026 24636 8032
rect 25240 7886 25268 8774
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25608 8430 25636 8570
rect 25596 8424 25648 8430
rect 25596 8366 25648 8372
rect 26252 7954 26280 8842
rect 26712 8838 26740 9998
rect 26700 8832 26752 8838
rect 26700 8774 26752 8780
rect 27356 8650 27384 11562
rect 27448 11286 27476 12242
rect 27620 12232 27672 12238
rect 27620 12174 27672 12180
rect 27632 11762 27660 12174
rect 28000 11898 28028 12854
rect 28320 12540 28628 12549
rect 28320 12538 28326 12540
rect 28382 12538 28406 12540
rect 28462 12538 28486 12540
rect 28542 12538 28566 12540
rect 28622 12538 28628 12540
rect 28382 12486 28384 12538
rect 28564 12486 28566 12538
rect 28320 12484 28326 12486
rect 28382 12484 28406 12486
rect 28462 12484 28486 12486
rect 28542 12484 28566 12486
rect 28622 12484 28628 12486
rect 28320 12475 28628 12484
rect 28736 12434 28764 13126
rect 29460 12776 29512 12782
rect 29460 12718 29512 12724
rect 30196 12776 30248 12782
rect 30196 12718 30248 12724
rect 29092 12640 29144 12646
rect 29092 12582 29144 12588
rect 29104 12442 29132 12582
rect 29472 12442 29500 12718
rect 30208 12646 30236 12718
rect 30196 12640 30248 12646
rect 30196 12582 30248 12588
rect 28644 12406 28764 12434
rect 29092 12436 29144 12442
rect 28644 12102 28672 12406
rect 29092 12378 29144 12384
rect 29460 12436 29512 12442
rect 29460 12378 29512 12384
rect 29920 12436 29972 12442
rect 29920 12378 29972 12384
rect 29104 12238 29132 12378
rect 29092 12232 29144 12238
rect 29092 12174 29144 12180
rect 29932 12102 29960 12378
rect 30208 12322 30236 12582
rect 30300 12434 30328 13262
rect 30472 13184 30524 13190
rect 30472 13126 30524 13132
rect 30484 12918 30512 13126
rect 30472 12912 30524 12918
rect 30472 12854 30524 12860
rect 30748 12844 30800 12850
rect 30748 12786 30800 12792
rect 30472 12640 30524 12646
rect 30472 12582 30524 12588
rect 30484 12442 30512 12582
rect 30472 12436 30524 12442
rect 30300 12406 30420 12434
rect 30392 12322 30420 12406
rect 30472 12378 30524 12384
rect 30564 12436 30616 12442
rect 30564 12378 30616 12384
rect 30576 12322 30604 12378
rect 30760 12374 30788 12786
rect 30208 12294 30328 12322
rect 30300 12238 30328 12294
rect 30392 12294 30604 12322
rect 30748 12368 30800 12374
rect 30748 12310 30800 12316
rect 31300 12300 31352 12306
rect 30012 12232 30064 12238
rect 30012 12174 30064 12180
rect 30288 12232 30340 12238
rect 30288 12174 30340 12180
rect 28632 12096 28684 12102
rect 28632 12038 28684 12044
rect 29920 12096 29972 12102
rect 29920 12038 29972 12044
rect 28644 11898 28672 12038
rect 27988 11892 28040 11898
rect 27988 11834 28040 11840
rect 28632 11892 28684 11898
rect 28632 11834 28684 11840
rect 29920 11892 29972 11898
rect 29920 11834 29972 11840
rect 29460 11824 29512 11830
rect 29458 11792 29460 11801
rect 29512 11792 29514 11801
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 28816 11756 28868 11762
rect 29458 11727 29514 11736
rect 29736 11756 29788 11762
rect 28816 11698 28868 11704
rect 29736 11698 29788 11704
rect 28320 11452 28628 11461
rect 28320 11450 28326 11452
rect 28382 11450 28406 11452
rect 28462 11450 28486 11452
rect 28542 11450 28566 11452
rect 28622 11450 28628 11452
rect 28382 11398 28384 11450
rect 28564 11398 28566 11450
rect 28320 11396 28326 11398
rect 28382 11396 28406 11398
rect 28462 11396 28486 11398
rect 28542 11396 28566 11398
rect 28622 11396 28628 11398
rect 28320 11387 28628 11396
rect 27436 11280 27488 11286
rect 27436 11222 27488 11228
rect 27620 11144 27672 11150
rect 27620 11086 27672 11092
rect 27528 10056 27580 10062
rect 27528 9998 27580 10004
rect 27436 9920 27488 9926
rect 27436 9862 27488 9868
rect 27448 8974 27476 9862
rect 27540 9722 27568 9998
rect 27632 9994 27660 11086
rect 28828 10674 28856 11698
rect 29748 11286 29776 11698
rect 29736 11280 29788 11286
rect 29736 11222 29788 11228
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 28816 10668 28868 10674
rect 28816 10610 28868 10616
rect 28320 10364 28628 10373
rect 28320 10362 28326 10364
rect 28382 10362 28406 10364
rect 28462 10362 28486 10364
rect 28542 10362 28566 10364
rect 28622 10362 28628 10364
rect 28382 10310 28384 10362
rect 28564 10310 28566 10362
rect 28320 10308 28326 10310
rect 28382 10308 28406 10310
rect 28462 10308 28486 10310
rect 28542 10308 28566 10310
rect 28622 10308 28628 10310
rect 28320 10299 28628 10308
rect 27620 9988 27672 9994
rect 27620 9930 27672 9936
rect 27528 9716 27580 9722
rect 27528 9658 27580 9664
rect 27632 8974 27660 9930
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 28460 9654 28488 9862
rect 28448 9648 28500 9654
rect 28448 9590 28500 9596
rect 27804 9512 27856 9518
rect 27804 9454 27856 9460
rect 27816 9178 27844 9454
rect 28320 9276 28628 9285
rect 28320 9274 28326 9276
rect 28382 9274 28406 9276
rect 28462 9274 28486 9276
rect 28542 9274 28566 9276
rect 28622 9274 28628 9276
rect 28382 9222 28384 9274
rect 28564 9222 28566 9274
rect 28320 9220 28326 9222
rect 28382 9220 28406 9222
rect 28462 9220 28486 9222
rect 28542 9220 28566 9222
rect 28622 9220 28628 9222
rect 28320 9211 28628 9220
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 28736 9042 28764 10610
rect 28828 10130 28856 10610
rect 28816 10124 28868 10130
rect 28816 10066 28868 10072
rect 29932 9994 29960 11834
rect 30024 11286 30052 12174
rect 30196 12164 30248 12170
rect 30196 12106 30248 12112
rect 30012 11280 30064 11286
rect 30012 11222 30064 11228
rect 30012 11144 30064 11150
rect 30012 11086 30064 11092
rect 29920 9988 29972 9994
rect 29920 9930 29972 9936
rect 30024 9926 30052 11086
rect 30208 11014 30236 12106
rect 30196 11008 30248 11014
rect 30196 10950 30248 10956
rect 30300 10606 30328 12174
rect 30392 12170 30420 12294
rect 31300 12242 31352 12248
rect 30380 12164 30432 12170
rect 30380 12106 30432 12112
rect 30656 12164 30708 12170
rect 30656 12106 30708 12112
rect 30668 11898 30696 12106
rect 30748 12096 30800 12102
rect 30748 12038 30800 12044
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 30656 11892 30708 11898
rect 30656 11834 30708 11840
rect 30656 11620 30708 11626
rect 30656 11562 30708 11568
rect 30668 11354 30696 11562
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30760 11150 30788 12038
rect 31220 11694 31248 12038
rect 31312 11694 31340 12242
rect 30840 11688 30892 11694
rect 30840 11630 30892 11636
rect 31208 11688 31260 11694
rect 31208 11630 31260 11636
rect 31300 11688 31352 11694
rect 31300 11630 31352 11636
rect 30852 11286 30880 11630
rect 31944 11552 31996 11558
rect 31944 11494 31996 11500
rect 30840 11280 30892 11286
rect 30840 11222 30892 11228
rect 31956 11150 31984 11494
rect 32324 11150 32352 13262
rect 33232 13252 33284 13258
rect 33232 13194 33284 13200
rect 33140 12436 33192 12442
rect 33140 12378 33192 12384
rect 33152 11694 33180 12378
rect 33244 11898 33272 13194
rect 33336 12238 33364 13262
rect 33600 12640 33652 12646
rect 33600 12582 33652 12588
rect 33324 12232 33376 12238
rect 33324 12174 33376 12180
rect 33508 12164 33560 12170
rect 33508 12106 33560 12112
rect 33520 11898 33548 12106
rect 33232 11892 33284 11898
rect 33232 11834 33284 11840
rect 33508 11892 33560 11898
rect 33508 11834 33560 11840
rect 33232 11756 33284 11762
rect 33232 11698 33284 11704
rect 33416 11756 33468 11762
rect 33416 11698 33468 11704
rect 32772 11688 32824 11694
rect 32772 11630 32824 11636
rect 33140 11688 33192 11694
rect 33140 11630 33192 11636
rect 30656 11144 30708 11150
rect 30656 11086 30708 11092
rect 30748 11144 30800 11150
rect 30748 11086 30800 11092
rect 31944 11144 31996 11150
rect 31944 11086 31996 11092
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32588 11144 32640 11150
rect 32588 11086 32640 11092
rect 30380 11076 30432 11082
rect 30380 11018 30432 11024
rect 30288 10600 30340 10606
rect 30288 10542 30340 10548
rect 30300 10130 30328 10542
rect 30288 10124 30340 10130
rect 30288 10066 30340 10072
rect 30392 9994 30420 11018
rect 30380 9988 30432 9994
rect 30380 9930 30432 9936
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 30024 9722 30052 9862
rect 30012 9716 30064 9722
rect 30012 9658 30064 9664
rect 30380 9580 30432 9586
rect 30380 9522 30432 9528
rect 29644 9512 29696 9518
rect 29644 9454 29696 9460
rect 28724 9036 28776 9042
rect 28724 8978 28776 8984
rect 27436 8968 27488 8974
rect 27436 8910 27488 8916
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 28448 8968 28500 8974
rect 28448 8910 28500 8916
rect 27620 8832 27672 8838
rect 27540 8780 27620 8786
rect 27540 8774 27672 8780
rect 27540 8758 27660 8774
rect 27356 8622 27476 8650
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 26240 7948 26292 7954
rect 26240 7890 26292 7896
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 26054 7848 26110 7857
rect 26054 7783 26110 7792
rect 22846 7644 23154 7653
rect 22846 7642 22852 7644
rect 22908 7642 22932 7644
rect 22988 7642 23012 7644
rect 23068 7642 23092 7644
rect 23148 7642 23154 7644
rect 22908 7590 22910 7642
rect 23090 7590 23092 7642
rect 22846 7588 22852 7590
rect 22908 7588 22932 7590
rect 22988 7588 23012 7590
rect 23068 7588 23092 7590
rect 23148 7588 23154 7590
rect 22846 7579 23154 7588
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 23308 7002 23336 7346
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 22846 6556 23154 6565
rect 22846 6554 22852 6556
rect 22908 6554 22932 6556
rect 22988 6554 23012 6556
rect 23068 6554 23092 6556
rect 23148 6554 23154 6556
rect 22908 6502 22910 6554
rect 23090 6502 23092 6554
rect 22846 6500 22852 6502
rect 22908 6500 22932 6502
rect 22988 6500 23012 6502
rect 23068 6500 23092 6502
rect 23148 6500 23154 6502
rect 22846 6491 23154 6500
rect 23308 6254 23336 6938
rect 24044 6322 24072 7346
rect 26068 7342 26096 7783
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 26160 7546 26188 7686
rect 26148 7540 26200 7546
rect 26148 7482 26200 7488
rect 26056 7336 26108 7342
rect 26056 7278 26108 7284
rect 25780 7200 25832 7206
rect 25780 7142 25832 7148
rect 25792 6798 25820 7142
rect 26068 7002 26096 7278
rect 26148 7268 26200 7274
rect 26148 7210 26200 7216
rect 26056 6996 26108 7002
rect 26056 6938 26108 6944
rect 26160 6798 26188 7210
rect 26252 6866 26280 7890
rect 26332 7812 26384 7818
rect 26332 7754 26384 7760
rect 26240 6860 26292 6866
rect 26240 6802 26292 6808
rect 25780 6792 25832 6798
rect 25780 6734 25832 6740
rect 26148 6792 26200 6798
rect 26344 6746 26372 7754
rect 26988 7410 27016 8230
rect 27356 7546 27384 8434
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 26976 7404 27028 7410
rect 26976 7346 27028 7352
rect 27448 6905 27476 8622
rect 27540 8430 27568 8758
rect 28460 8566 28488 8910
rect 27712 8560 27764 8566
rect 27712 8502 27764 8508
rect 28448 8560 28500 8566
rect 28448 8502 28500 8508
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 27434 6896 27490 6905
rect 26976 6860 27028 6866
rect 27434 6831 27490 6840
rect 26976 6802 27028 6808
rect 26148 6734 26200 6740
rect 26252 6718 26372 6746
rect 26252 6662 26280 6718
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 26424 6656 26476 6662
rect 26424 6598 26476 6604
rect 26436 6322 26464 6598
rect 26988 6322 27016 6802
rect 27344 6724 27396 6730
rect 27344 6666 27396 6672
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 26424 6316 26476 6322
rect 26424 6258 26476 6264
rect 26976 6316 27028 6322
rect 26976 6258 27028 6264
rect 23296 6248 23348 6254
rect 23296 6190 23348 6196
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 22940 5778 22968 6054
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22846 5468 23154 5477
rect 22846 5466 22852 5468
rect 22908 5466 22932 5468
rect 22988 5466 23012 5468
rect 23068 5466 23092 5468
rect 23148 5466 23154 5468
rect 22908 5414 22910 5466
rect 23090 5414 23092 5466
rect 22846 5412 22852 5414
rect 22908 5412 22932 5414
rect 22988 5412 23012 5414
rect 23068 5412 23092 5414
rect 23148 5412 23154 5414
rect 22846 5403 23154 5412
rect 23112 5228 23164 5234
rect 23112 5170 23164 5176
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22756 3942 22784 4966
rect 23124 4690 23152 5170
rect 23492 5166 23520 5850
rect 24044 5574 24072 6258
rect 26884 6248 26936 6254
rect 26884 6190 26936 6196
rect 24400 6112 24452 6118
rect 24400 6054 24452 6060
rect 24412 5710 24440 6054
rect 26896 5914 26924 6190
rect 26792 5908 26844 5914
rect 26792 5850 26844 5856
rect 26884 5908 26936 5914
rect 26884 5850 26936 5856
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 24676 5704 24728 5710
rect 26424 5704 26476 5710
rect 24676 5646 24728 5652
rect 26422 5672 26424 5681
rect 26476 5672 26478 5681
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 24308 5568 24360 5574
rect 24308 5510 24360 5516
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23112 4684 23164 4690
rect 23112 4626 23164 4632
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 22846 4380 23154 4389
rect 22846 4378 22852 4380
rect 22908 4378 22932 4380
rect 22988 4378 23012 4380
rect 23068 4378 23092 4380
rect 23148 4378 23154 4380
rect 22908 4326 22910 4378
rect 23090 4326 23092 4378
rect 22846 4324 22852 4326
rect 22908 4324 22932 4326
rect 22988 4324 23012 4326
rect 23068 4324 23092 4326
rect 23148 4324 23154 4326
rect 22846 4315 23154 4324
rect 22744 3936 22796 3942
rect 22744 3878 22796 3884
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22756 3058 22784 3470
rect 22846 3292 23154 3301
rect 22846 3290 22852 3292
rect 22908 3290 22932 3292
rect 22988 3290 23012 3292
rect 23068 3290 23092 3292
rect 23148 3290 23154 3292
rect 22908 3238 22910 3290
rect 23090 3238 23092 3290
rect 22846 3236 22852 3238
rect 22908 3236 22932 3238
rect 22988 3236 23012 3238
rect 23068 3236 23092 3238
rect 23148 3236 23154 3238
rect 22846 3227 23154 3236
rect 23216 3194 23244 4558
rect 23388 4072 23440 4078
rect 23388 4014 23440 4020
rect 23400 3194 23428 4014
rect 23584 3738 23612 4966
rect 23860 3942 23888 5170
rect 24320 4146 24348 5510
rect 24688 5098 24716 5646
rect 26422 5607 26478 5616
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 25136 5228 25188 5234
rect 25136 5170 25188 5176
rect 25320 5228 25372 5234
rect 25320 5170 25372 5176
rect 25504 5228 25556 5234
rect 25504 5170 25556 5176
rect 24860 5160 24912 5166
rect 24860 5102 24912 5108
rect 24676 5092 24728 5098
rect 24676 5034 24728 5040
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 24412 4826 24440 4966
rect 24872 4826 24900 5102
rect 25056 4826 25084 5170
rect 25148 4826 25176 5170
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 24860 4820 24912 4826
rect 24860 4762 24912 4768
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 24872 4214 24900 4762
rect 24400 4208 24452 4214
rect 24400 4150 24452 4156
rect 24860 4208 24912 4214
rect 24860 4150 24912 4156
rect 24308 4140 24360 4146
rect 24308 4082 24360 4088
rect 23848 3936 23900 3942
rect 23848 3878 23900 3884
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23756 3732 23808 3738
rect 23756 3674 23808 3680
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 23768 3058 23796 3674
rect 23860 3670 23888 3878
rect 24412 3738 24440 4150
rect 25056 4146 25084 4762
rect 25332 4282 25360 5170
rect 25320 4276 25372 4282
rect 25320 4218 25372 4224
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24780 3670 24808 4014
rect 25516 4010 25544 5170
rect 26804 4978 26832 5850
rect 26804 4950 26924 4978
rect 26896 4826 26924 4950
rect 26148 4820 26200 4826
rect 26148 4762 26200 4768
rect 26884 4820 26936 4826
rect 26884 4762 26936 4768
rect 26056 4616 26108 4622
rect 26056 4558 26108 4564
rect 26068 4146 26096 4558
rect 26160 4282 26188 4762
rect 26608 4548 26660 4554
rect 26608 4490 26660 4496
rect 26148 4276 26200 4282
rect 26148 4218 26200 4224
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 25504 4004 25556 4010
rect 25504 3946 25556 3952
rect 25044 3936 25096 3942
rect 25044 3878 25096 3884
rect 23848 3664 23900 3670
rect 23848 3606 23900 3612
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 25056 3466 25084 3878
rect 25044 3460 25096 3466
rect 25044 3402 25096 3408
rect 26620 3398 26648 4490
rect 26988 4146 27016 6258
rect 27356 5234 27384 6666
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 27252 4480 27304 4486
rect 27252 4422 27304 4428
rect 26976 4140 27028 4146
rect 26976 4082 27028 4088
rect 27264 3534 27292 4422
rect 27252 3528 27304 3534
rect 27252 3470 27304 3476
rect 26608 3392 26660 3398
rect 26608 3334 26660 3340
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 19720 2746 19840 2774
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 1582 1456 1638 1465
rect 1582 1391 1638 1400
rect 3252 800 3280 2382
rect 4540 800 4568 2382
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6472 800 6500 2246
rect 7760 800 7788 2382
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 800 9720 2246
rect 10980 800 11008 2382
rect 11898 2204 12206 2213
rect 11898 2202 11904 2204
rect 11960 2202 11984 2204
rect 12040 2202 12064 2204
rect 12120 2202 12144 2204
rect 12200 2202 12206 2204
rect 11960 2150 11962 2202
rect 12142 2150 12144 2202
rect 11898 2148 11904 2150
rect 11960 2148 11984 2150
rect 12040 2148 12064 2150
rect 12120 2148 12144 2150
rect 12200 2148 12206 2150
rect 11898 2139 12206 2148
rect 12912 800 12940 2382
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 800 14228 2246
rect 16132 800 16160 2382
rect 17420 800 17448 2382
rect 19352 800 19380 2382
rect 19720 2378 19748 2746
rect 22664 2446 22692 2790
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 19708 2372 19760 2378
rect 19708 2314 19760 2320
rect 20640 800 20668 2382
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22572 800 22600 2246
rect 22846 2204 23154 2213
rect 22846 2202 22852 2204
rect 22908 2202 22932 2204
rect 22988 2202 23012 2204
rect 23068 2202 23092 2204
rect 23148 2202 23154 2204
rect 22908 2150 22910 2202
rect 23090 2150 23092 2202
rect 22846 2148 22852 2150
rect 22908 2148 22932 2150
rect 22988 2148 23012 2150
rect 23068 2148 23092 2150
rect 23148 2148 23154 2150
rect 22846 2139 23154 2148
rect 23860 800 23888 2382
rect 25792 800 25820 2382
rect 27080 800 27108 2382
rect 27448 2310 27476 6831
rect 27540 5302 27568 8366
rect 27724 7954 27752 8502
rect 28320 8188 28628 8197
rect 28320 8186 28326 8188
rect 28382 8186 28406 8188
rect 28462 8186 28486 8188
rect 28542 8186 28566 8188
rect 28622 8186 28628 8188
rect 28382 8134 28384 8186
rect 28564 8134 28566 8186
rect 28320 8132 28326 8134
rect 28382 8132 28406 8134
rect 28462 8132 28486 8134
rect 28542 8132 28566 8134
rect 28622 8132 28628 8134
rect 28320 8123 28628 8132
rect 27712 7948 27764 7954
rect 27712 7890 27764 7896
rect 27724 7449 27752 7890
rect 28264 7744 28316 7750
rect 28264 7686 28316 7692
rect 28276 7478 28304 7686
rect 28264 7472 28316 7478
rect 27710 7440 27766 7449
rect 28264 7414 28316 7420
rect 28736 7410 28764 8978
rect 29552 8900 29604 8906
rect 29552 8842 29604 8848
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 29000 8832 29052 8838
rect 29000 8774 29052 8780
rect 28920 8566 28948 8774
rect 28908 8560 28960 8566
rect 28908 8502 28960 8508
rect 29012 8498 29040 8774
rect 29564 8498 29592 8842
rect 29000 8492 29052 8498
rect 29000 8434 29052 8440
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 28828 7954 28856 8366
rect 28816 7948 28868 7954
rect 28816 7890 28868 7896
rect 28816 7744 28868 7750
rect 28816 7686 28868 7692
rect 28828 7546 28856 7686
rect 29656 7546 29684 9454
rect 29828 9376 29880 9382
rect 29828 9318 29880 9324
rect 29840 8974 29868 9318
rect 30392 9178 30420 9522
rect 30668 9500 30696 11086
rect 31576 9648 31628 9654
rect 31576 9590 31628 9596
rect 31116 9580 31168 9586
rect 31116 9522 31168 9528
rect 30668 9472 30788 9500
rect 30380 9172 30432 9178
rect 30380 9114 30432 9120
rect 30760 8974 30788 9472
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 30748 8968 30800 8974
rect 30748 8910 30800 8916
rect 29828 8492 29880 8498
rect 29828 8434 29880 8440
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 29736 7880 29788 7886
rect 29736 7822 29788 7828
rect 28816 7540 28868 7546
rect 28816 7482 28868 7488
rect 29644 7540 29696 7546
rect 29644 7482 29696 7488
rect 27710 7375 27766 7384
rect 28724 7404 28776 7410
rect 27724 7342 27752 7375
rect 28724 7346 28776 7352
rect 27712 7336 27764 7342
rect 27712 7278 27764 7284
rect 28320 7100 28628 7109
rect 28320 7098 28326 7100
rect 28382 7098 28406 7100
rect 28462 7098 28486 7100
rect 28542 7098 28566 7100
rect 28622 7098 28628 7100
rect 28382 7046 28384 7098
rect 28564 7046 28566 7098
rect 28320 7044 28326 7046
rect 28382 7044 28406 7046
rect 28462 7044 28486 7046
rect 28542 7044 28566 7046
rect 28622 7044 28628 7046
rect 28320 7035 28628 7044
rect 28828 7002 28856 7482
rect 27712 6996 27764 7002
rect 27712 6938 27764 6944
rect 28816 6996 28868 7002
rect 28816 6938 28868 6944
rect 27620 5704 27672 5710
rect 27724 5692 27752 6938
rect 29748 6866 29776 7822
rect 29736 6860 29788 6866
rect 29736 6802 29788 6808
rect 29092 6656 29144 6662
rect 29092 6598 29144 6604
rect 29104 6118 29132 6598
rect 29000 6112 29052 6118
rect 29000 6054 29052 6060
rect 29092 6112 29144 6118
rect 29092 6054 29144 6060
rect 28320 6012 28628 6021
rect 28320 6010 28326 6012
rect 28382 6010 28406 6012
rect 28462 6010 28486 6012
rect 28542 6010 28566 6012
rect 28622 6010 28628 6012
rect 28382 5958 28384 6010
rect 28564 5958 28566 6010
rect 28320 5956 28326 5958
rect 28382 5956 28406 5958
rect 28462 5956 28486 5958
rect 28542 5956 28566 5958
rect 28622 5956 28628 5958
rect 28320 5947 28628 5956
rect 29012 5846 29040 6054
rect 28356 5840 28408 5846
rect 28356 5782 28408 5788
rect 29000 5840 29052 5846
rect 29000 5782 29052 5788
rect 29644 5840 29696 5846
rect 29644 5782 29696 5788
rect 28368 5710 28396 5782
rect 29012 5710 29040 5782
rect 27804 5704 27856 5710
rect 27724 5672 27804 5692
rect 28356 5704 28408 5710
rect 27856 5672 27858 5681
rect 27724 5664 27802 5672
rect 27620 5646 27672 5652
rect 27528 5296 27580 5302
rect 27528 5238 27580 5244
rect 27632 5098 27660 5646
rect 29000 5704 29052 5710
rect 28356 5646 28408 5652
rect 28630 5672 28686 5681
rect 27802 5607 27858 5616
rect 29000 5646 29052 5652
rect 29656 5642 29684 5782
rect 28630 5607 28686 5616
rect 29644 5636 29696 5642
rect 28644 5574 28672 5607
rect 29644 5578 29696 5584
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 28540 5568 28592 5574
rect 28540 5510 28592 5516
rect 28632 5568 28684 5574
rect 28632 5510 28684 5516
rect 27620 5092 27672 5098
rect 27620 5034 27672 5040
rect 28184 5030 28212 5510
rect 28552 5302 28580 5510
rect 28448 5296 28500 5302
rect 28448 5238 28500 5244
rect 28540 5296 28592 5302
rect 28540 5238 28592 5244
rect 28460 5166 28488 5238
rect 28448 5160 28500 5166
rect 28448 5102 28500 5108
rect 29276 5160 29328 5166
rect 29276 5102 29328 5108
rect 29368 5160 29420 5166
rect 29368 5102 29420 5108
rect 28172 5024 28224 5030
rect 28172 4966 28224 4972
rect 28320 4924 28628 4933
rect 28320 4922 28326 4924
rect 28382 4922 28406 4924
rect 28462 4922 28486 4924
rect 28542 4922 28566 4924
rect 28622 4922 28628 4924
rect 28382 4870 28384 4922
rect 28564 4870 28566 4922
rect 28320 4868 28326 4870
rect 28382 4868 28406 4870
rect 28462 4868 28486 4870
rect 28542 4868 28566 4870
rect 28622 4868 28628 4870
rect 28320 4859 28628 4868
rect 29092 4820 29144 4826
rect 29092 4762 29144 4768
rect 27620 4548 27672 4554
rect 27620 4490 27672 4496
rect 27632 4214 27660 4490
rect 29104 4282 29132 4762
rect 29288 4758 29316 5102
rect 29276 4752 29328 4758
rect 29276 4694 29328 4700
rect 29184 4480 29236 4486
rect 29184 4422 29236 4428
rect 29092 4276 29144 4282
rect 29092 4218 29144 4224
rect 27620 4208 27672 4214
rect 27620 4150 27672 4156
rect 28080 4208 28132 4214
rect 28080 4150 28132 4156
rect 27632 4078 27660 4150
rect 27528 4072 27580 4078
rect 27528 4014 27580 4020
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27540 3738 27568 4014
rect 28092 3738 28120 4150
rect 29092 3936 29144 3942
rect 29092 3878 29144 3884
rect 28320 3836 28628 3845
rect 28320 3834 28326 3836
rect 28382 3834 28406 3836
rect 28462 3834 28486 3836
rect 28542 3834 28566 3836
rect 28622 3834 28628 3836
rect 28382 3782 28384 3834
rect 28564 3782 28566 3834
rect 28320 3780 28326 3782
rect 28382 3780 28406 3782
rect 28462 3780 28486 3782
rect 28542 3780 28566 3782
rect 28622 3780 28628 3782
rect 28320 3771 28628 3780
rect 27528 3732 27580 3738
rect 27528 3674 27580 3680
rect 28080 3732 28132 3738
rect 28080 3674 28132 3680
rect 29104 3534 29132 3878
rect 29196 3534 29224 4422
rect 29380 4078 29408 5102
rect 29460 4820 29512 4826
rect 29460 4762 29512 4768
rect 29472 4622 29500 4762
rect 29552 4684 29604 4690
rect 29748 4672 29776 6802
rect 29840 6458 29868 8434
rect 30024 7750 30052 8434
rect 30288 8288 30340 8294
rect 30288 8230 30340 8236
rect 30300 7886 30328 8230
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 30012 7744 30064 7750
rect 30012 7686 30064 7692
rect 30024 7478 30052 7686
rect 30012 7472 30064 7478
rect 30012 7414 30064 7420
rect 30380 7404 30432 7410
rect 30380 7346 30432 7352
rect 29920 7336 29972 7342
rect 29920 7278 29972 7284
rect 29828 6452 29880 6458
rect 29828 6394 29880 6400
rect 29932 6254 29960 7278
rect 29920 6248 29972 6254
rect 29920 6190 29972 6196
rect 29828 5704 29880 5710
rect 29828 5646 29880 5652
rect 29840 5234 29868 5646
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 29932 5166 29960 6190
rect 30012 6180 30064 6186
rect 30012 6122 30064 6128
rect 30024 5710 30052 6122
rect 30392 5710 30420 7346
rect 31024 7200 31076 7206
rect 31024 7142 31076 7148
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30484 6322 30512 6598
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30012 5704 30064 5710
rect 30012 5646 30064 5652
rect 30380 5704 30432 5710
rect 30380 5646 30432 5652
rect 30484 5302 30512 6258
rect 30932 5908 30984 5914
rect 30932 5850 30984 5856
rect 30748 5636 30800 5642
rect 30748 5578 30800 5584
rect 30472 5296 30524 5302
rect 30472 5238 30524 5244
rect 30760 5234 30788 5578
rect 30944 5302 30972 5850
rect 31036 5846 31064 7142
rect 31128 6934 31156 9522
rect 31588 9110 31616 9590
rect 31576 9104 31628 9110
rect 31576 9046 31628 9052
rect 31668 9104 31720 9110
rect 31668 9046 31720 9052
rect 31588 8974 31616 9046
rect 31484 8968 31536 8974
rect 31484 8910 31536 8916
rect 31576 8968 31628 8974
rect 31576 8910 31628 8916
rect 31496 8362 31524 8910
rect 31680 8838 31708 9046
rect 31956 9042 31984 11086
rect 32324 10810 32352 11086
rect 32312 10804 32364 10810
rect 32312 10746 32364 10752
rect 32324 9042 32352 10746
rect 32600 10674 32628 11086
rect 32588 10668 32640 10674
rect 32588 10610 32640 10616
rect 32784 10470 32812 11630
rect 32496 10464 32548 10470
rect 32496 10406 32548 10412
rect 32772 10464 32824 10470
rect 32772 10406 32824 10412
rect 32508 9994 32536 10406
rect 33244 10266 33272 11698
rect 33428 11354 33456 11698
rect 33416 11348 33468 11354
rect 33416 11290 33468 11296
rect 33232 10260 33284 10266
rect 33232 10202 33284 10208
rect 32496 9988 32548 9994
rect 32496 9930 32548 9936
rect 33244 9586 33272 10202
rect 32680 9580 32732 9586
rect 32680 9522 32732 9528
rect 32772 9580 32824 9586
rect 32772 9522 32824 9528
rect 33232 9580 33284 9586
rect 33232 9522 33284 9528
rect 33416 9580 33468 9586
rect 33416 9522 33468 9528
rect 31944 9036 31996 9042
rect 31944 8978 31996 8984
rect 32312 9036 32364 9042
rect 32312 8978 32364 8984
rect 32692 8838 32720 9522
rect 32784 9178 32812 9522
rect 33140 9512 33192 9518
rect 33140 9454 33192 9460
rect 32772 9172 32824 9178
rect 32772 9114 32824 9120
rect 31668 8832 31720 8838
rect 31668 8774 31720 8780
rect 32680 8832 32732 8838
rect 32680 8774 32732 8780
rect 32402 8528 32458 8537
rect 32128 8492 32180 8498
rect 32402 8463 32404 8472
rect 32128 8434 32180 8440
rect 32456 8463 32458 8472
rect 33048 8492 33100 8498
rect 32404 8434 32456 8440
rect 33048 8434 33100 8440
rect 31484 8356 31536 8362
rect 31484 8298 31536 8304
rect 32140 7750 32168 8434
rect 32496 8356 32548 8362
rect 32496 8298 32548 8304
rect 32220 7880 32272 7886
rect 32220 7822 32272 7828
rect 32128 7744 32180 7750
rect 32128 7686 32180 7692
rect 32232 7410 32260 7822
rect 32508 7818 32536 8298
rect 32864 8288 32916 8294
rect 32864 8230 32916 8236
rect 32876 8090 32904 8230
rect 32864 8084 32916 8090
rect 32864 8026 32916 8032
rect 32312 7812 32364 7818
rect 32312 7754 32364 7760
rect 32496 7812 32548 7818
rect 32496 7754 32548 7760
rect 32324 7478 32352 7754
rect 32588 7540 32640 7546
rect 32588 7482 32640 7488
rect 32312 7472 32364 7478
rect 32312 7414 32364 7420
rect 32128 7404 32180 7410
rect 32128 7346 32180 7352
rect 32220 7404 32272 7410
rect 32220 7346 32272 7352
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 31116 6928 31168 6934
rect 31116 6870 31168 6876
rect 31312 6866 31340 7278
rect 31300 6860 31352 6866
rect 31300 6802 31352 6808
rect 32036 6724 32088 6730
rect 32036 6666 32088 6672
rect 31852 6452 31904 6458
rect 32048 6440 32076 6666
rect 31904 6412 32076 6440
rect 31852 6394 31904 6400
rect 31576 6384 31628 6390
rect 31576 6326 31628 6332
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 31116 6112 31168 6118
rect 31116 6054 31168 6060
rect 31128 5914 31156 6054
rect 31116 5908 31168 5914
rect 31116 5850 31168 5856
rect 31024 5840 31076 5846
rect 31024 5782 31076 5788
rect 30932 5296 30984 5302
rect 30932 5238 30984 5244
rect 30748 5228 30800 5234
rect 30748 5170 30800 5176
rect 29920 5160 29972 5166
rect 29920 5102 29972 5108
rect 30944 5098 30972 5238
rect 30932 5092 30984 5098
rect 30932 5034 30984 5040
rect 29604 4644 29776 4672
rect 29552 4626 29604 4632
rect 29460 4616 29512 4622
rect 29460 4558 29512 4564
rect 30932 4616 30984 4622
rect 30932 4558 30984 4564
rect 29472 4146 29500 4558
rect 29828 4548 29880 4554
rect 29828 4490 29880 4496
rect 29460 4140 29512 4146
rect 29460 4082 29512 4088
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 29092 3528 29144 3534
rect 29092 3470 29144 3476
rect 29184 3528 29236 3534
rect 29184 3470 29236 3476
rect 28000 3058 28028 3470
rect 29380 3398 29408 4014
rect 29840 3738 29868 4490
rect 30012 4480 30064 4486
rect 30012 4422 30064 4428
rect 30024 4146 30052 4422
rect 30564 4276 30616 4282
rect 30564 4218 30616 4224
rect 30012 4140 30064 4146
rect 30012 4082 30064 4088
rect 29828 3732 29880 3738
rect 29828 3674 29880 3680
rect 30576 3602 30604 4218
rect 30944 3738 30972 4558
rect 31312 4146 31340 6258
rect 31588 5642 31616 6326
rect 32140 6322 32168 7346
rect 32128 6316 32180 6322
rect 32128 6258 32180 6264
rect 32140 5794 32168 6258
rect 31956 5766 32168 5794
rect 31576 5636 31628 5642
rect 31576 5578 31628 5584
rect 31392 5568 31444 5574
rect 31392 5510 31444 5516
rect 31404 4486 31432 5510
rect 31956 5302 31984 5766
rect 32128 5704 32180 5710
rect 32128 5646 32180 5652
rect 31760 5296 31812 5302
rect 31760 5238 31812 5244
rect 31944 5296 31996 5302
rect 31944 5238 31996 5244
rect 31392 4480 31444 4486
rect 31392 4422 31444 4428
rect 31772 4214 31800 5238
rect 32140 5234 32168 5646
rect 32128 5228 32180 5234
rect 32128 5170 32180 5176
rect 31944 5024 31996 5030
rect 31944 4966 31996 4972
rect 31956 4554 31984 4966
rect 31944 4548 31996 4554
rect 31944 4490 31996 4496
rect 31760 4208 31812 4214
rect 31760 4150 31812 4156
rect 31300 4140 31352 4146
rect 31300 4082 31352 4088
rect 31312 3942 31340 4082
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 30932 3732 30984 3738
rect 30932 3674 30984 3680
rect 30564 3596 30616 3602
rect 30564 3538 30616 3544
rect 31772 3534 31800 4150
rect 30932 3528 30984 3534
rect 30932 3470 30984 3476
rect 31760 3528 31812 3534
rect 31760 3470 31812 3476
rect 29368 3392 29420 3398
rect 29368 3334 29420 3340
rect 30944 3058 30972 3470
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 30932 3052 30984 3058
rect 30932 2994 30984 3000
rect 28320 2748 28628 2757
rect 28320 2746 28326 2748
rect 28382 2746 28406 2748
rect 28462 2746 28486 2748
rect 28542 2746 28566 2748
rect 28622 2746 28628 2748
rect 28382 2694 28384 2746
rect 28564 2694 28566 2746
rect 28320 2692 28326 2694
rect 28382 2692 28406 2694
rect 28462 2692 28486 2694
rect 28542 2692 28566 2694
rect 28622 2692 28628 2694
rect 28320 2683 28628 2692
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 27436 2304 27488 2310
rect 27436 2246 27488 2252
rect 29012 800 29040 2382
rect 30300 800 30328 2382
rect 32220 2372 32272 2378
rect 32220 2314 32272 2320
rect 32232 800 32260 2314
rect 32324 2310 32352 7414
rect 32600 7002 32628 7482
rect 33060 7410 33088 8434
rect 32680 7404 32732 7410
rect 32680 7346 32732 7352
rect 33048 7404 33100 7410
rect 33048 7346 33100 7352
rect 32588 6996 32640 7002
rect 32588 6938 32640 6944
rect 32692 6866 32720 7346
rect 32772 7200 32824 7206
rect 32772 7142 32824 7148
rect 32680 6860 32732 6866
rect 32680 6802 32732 6808
rect 32692 6322 32720 6802
rect 32588 6316 32640 6322
rect 32588 6258 32640 6264
rect 32680 6316 32732 6322
rect 32680 6258 32732 6264
rect 32600 5030 32628 6258
rect 32692 5778 32720 6258
rect 32680 5772 32732 5778
rect 32680 5714 32732 5720
rect 32692 5234 32720 5714
rect 32680 5228 32732 5234
rect 32680 5170 32732 5176
rect 32588 5024 32640 5030
rect 32588 4966 32640 4972
rect 32600 3534 32628 4966
rect 32692 4214 32720 5170
rect 32784 4826 32812 7142
rect 33152 6905 33180 9454
rect 33232 8016 33284 8022
rect 33232 7958 33284 7964
rect 33138 6896 33194 6905
rect 33138 6831 33194 6840
rect 33244 6798 33272 7958
rect 33428 7478 33456 9522
rect 33612 9450 33640 12582
rect 33704 11218 33732 13738
rect 33794 13084 34102 13093
rect 33794 13082 33800 13084
rect 33856 13082 33880 13084
rect 33936 13082 33960 13084
rect 34016 13082 34040 13084
rect 34096 13082 34102 13084
rect 33856 13030 33858 13082
rect 34038 13030 34040 13082
rect 33794 13028 33800 13030
rect 33856 13028 33880 13030
rect 33936 13028 33960 13030
rect 34016 13028 34040 13030
rect 34096 13028 34102 13030
rect 33794 13019 34102 13028
rect 34164 12238 34192 16934
rect 34888 15496 34940 15502
rect 34888 15438 34940 15444
rect 34900 14074 34928 15438
rect 34888 14068 34940 14074
rect 34888 14010 34940 14016
rect 34520 13864 34572 13870
rect 34520 13806 34572 13812
rect 34532 12918 34560 13806
rect 37292 13394 37320 17274
rect 37384 17202 37412 19200
rect 38672 17270 38700 19200
rect 40604 17338 40632 19200
rect 40592 17332 40644 17338
rect 40592 17274 40644 17280
rect 38660 17264 38712 17270
rect 38660 17206 38712 17212
rect 41892 17202 41920 19200
rect 43442 19136 43498 19145
rect 43442 19071 43498 19080
rect 37372 17196 37424 17202
rect 37372 17138 37424 17144
rect 40684 17196 40736 17202
rect 40684 17138 40736 17144
rect 41880 17196 41932 17202
rect 41880 17138 41932 17144
rect 38936 16992 38988 16998
rect 38936 16934 38988 16940
rect 38948 13734 38976 16934
rect 39268 16892 39576 16901
rect 39268 16890 39274 16892
rect 39330 16890 39354 16892
rect 39410 16890 39434 16892
rect 39490 16890 39514 16892
rect 39570 16890 39576 16892
rect 39330 16838 39332 16890
rect 39512 16838 39514 16890
rect 39268 16836 39274 16838
rect 39330 16836 39354 16838
rect 39410 16836 39434 16838
rect 39490 16836 39514 16838
rect 39570 16836 39576 16838
rect 39268 16827 39576 16836
rect 40040 16584 40092 16590
rect 40040 16526 40092 16532
rect 39268 15804 39576 15813
rect 39268 15802 39274 15804
rect 39330 15802 39354 15804
rect 39410 15802 39434 15804
rect 39490 15802 39514 15804
rect 39570 15802 39576 15804
rect 39330 15750 39332 15802
rect 39512 15750 39514 15802
rect 39268 15748 39274 15750
rect 39330 15748 39354 15750
rect 39410 15748 39434 15750
rect 39490 15748 39514 15750
rect 39570 15748 39576 15750
rect 39268 15739 39576 15748
rect 39268 14716 39576 14725
rect 39268 14714 39274 14716
rect 39330 14714 39354 14716
rect 39410 14714 39434 14716
rect 39490 14714 39514 14716
rect 39570 14714 39576 14716
rect 39330 14662 39332 14714
rect 39512 14662 39514 14714
rect 39268 14660 39274 14662
rect 39330 14660 39354 14662
rect 39410 14660 39434 14662
rect 39490 14660 39514 14662
rect 39570 14660 39576 14662
rect 39268 14651 39576 14660
rect 38936 13728 38988 13734
rect 38936 13670 38988 13676
rect 39268 13628 39576 13637
rect 39268 13626 39274 13628
rect 39330 13626 39354 13628
rect 39410 13626 39434 13628
rect 39490 13626 39514 13628
rect 39570 13626 39576 13628
rect 39330 13574 39332 13626
rect 39512 13574 39514 13626
rect 39268 13572 39274 13574
rect 39330 13572 39354 13574
rect 39410 13572 39434 13574
rect 39490 13572 39514 13574
rect 39570 13572 39576 13574
rect 39268 13563 39576 13572
rect 37280 13388 37332 13394
rect 37280 13330 37332 13336
rect 38936 13388 38988 13394
rect 38936 13330 38988 13336
rect 37648 13320 37700 13326
rect 37648 13262 37700 13268
rect 38292 13320 38344 13326
rect 38292 13262 38344 13268
rect 38384 13320 38436 13326
rect 38384 13262 38436 13268
rect 35624 13184 35676 13190
rect 35624 13126 35676 13132
rect 35636 12986 35664 13126
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 34520 12912 34572 12918
rect 34520 12854 34572 12860
rect 34336 12844 34388 12850
rect 34336 12786 34388 12792
rect 34348 12442 34376 12786
rect 34532 12782 34560 12854
rect 37556 12844 37608 12850
rect 37556 12786 37608 12792
rect 34520 12776 34572 12782
rect 34520 12718 34572 12724
rect 37004 12776 37056 12782
rect 37004 12718 37056 12724
rect 34336 12436 34388 12442
rect 34336 12378 34388 12384
rect 34244 12300 34296 12306
rect 34244 12242 34296 12248
rect 36544 12300 36596 12306
rect 36544 12242 36596 12248
rect 34152 12232 34204 12238
rect 34152 12174 34204 12180
rect 33794 11996 34102 12005
rect 33794 11994 33800 11996
rect 33856 11994 33880 11996
rect 33936 11994 33960 11996
rect 34016 11994 34040 11996
rect 34096 11994 34102 11996
rect 33856 11942 33858 11994
rect 34038 11942 34040 11994
rect 33794 11940 33800 11942
rect 33856 11940 33880 11942
rect 33936 11940 33960 11942
rect 34016 11940 34040 11942
rect 34096 11940 34102 11942
rect 33794 11931 34102 11940
rect 34152 11756 34204 11762
rect 34152 11698 34204 11704
rect 33692 11212 33744 11218
rect 33692 11154 33744 11160
rect 33794 10908 34102 10917
rect 33794 10906 33800 10908
rect 33856 10906 33880 10908
rect 33936 10906 33960 10908
rect 34016 10906 34040 10908
rect 34096 10906 34102 10908
rect 33856 10854 33858 10906
rect 34038 10854 34040 10906
rect 33794 10852 33800 10854
rect 33856 10852 33880 10854
rect 33936 10852 33960 10854
rect 34016 10852 34040 10854
rect 34096 10852 34102 10854
rect 33794 10843 34102 10852
rect 34060 10532 34112 10538
rect 34060 10474 34112 10480
rect 34072 9908 34100 10474
rect 34164 10130 34192 11698
rect 34152 10124 34204 10130
rect 34152 10066 34204 10072
rect 34072 9880 34192 9908
rect 33794 9820 34102 9829
rect 33794 9818 33800 9820
rect 33856 9818 33880 9820
rect 33936 9818 33960 9820
rect 34016 9818 34040 9820
rect 34096 9818 34102 9820
rect 33856 9766 33858 9818
rect 34038 9766 34040 9818
rect 33794 9764 33800 9766
rect 33856 9764 33880 9766
rect 33936 9764 33960 9766
rect 34016 9764 34040 9766
rect 34096 9764 34102 9766
rect 33794 9755 34102 9764
rect 33600 9444 33652 9450
rect 33600 9386 33652 9392
rect 33692 8900 33744 8906
rect 33692 8842 33744 8848
rect 33704 8634 33732 8842
rect 33794 8732 34102 8741
rect 33794 8730 33800 8732
rect 33856 8730 33880 8732
rect 33936 8730 33960 8732
rect 34016 8730 34040 8732
rect 34096 8730 34102 8732
rect 33856 8678 33858 8730
rect 34038 8678 34040 8730
rect 33794 8676 33800 8678
rect 33856 8676 33880 8678
rect 33936 8676 33960 8678
rect 34016 8676 34040 8678
rect 34096 8676 34102 8678
rect 33794 8667 34102 8676
rect 33692 8628 33744 8634
rect 33692 8570 33744 8576
rect 33508 8356 33560 8362
rect 33508 8298 33560 8304
rect 33520 7954 33548 8298
rect 33508 7948 33560 7954
rect 33508 7890 33560 7896
rect 33704 7886 33732 8570
rect 33692 7880 33744 7886
rect 33692 7822 33744 7828
rect 33794 7644 34102 7653
rect 33794 7642 33800 7644
rect 33856 7642 33880 7644
rect 33936 7642 33960 7644
rect 34016 7642 34040 7644
rect 34096 7642 34102 7644
rect 33856 7590 33858 7642
rect 34038 7590 34040 7642
rect 33794 7588 33800 7590
rect 33856 7588 33880 7590
rect 33936 7588 33960 7590
rect 34016 7588 34040 7590
rect 34096 7588 34102 7590
rect 33794 7579 34102 7588
rect 33416 7472 33468 7478
rect 33416 7414 33468 7420
rect 33232 6792 33284 6798
rect 33232 6734 33284 6740
rect 33794 6556 34102 6565
rect 33794 6554 33800 6556
rect 33856 6554 33880 6556
rect 33936 6554 33960 6556
rect 34016 6554 34040 6556
rect 34096 6554 34102 6556
rect 33856 6502 33858 6554
rect 34038 6502 34040 6554
rect 33794 6500 33800 6502
rect 33856 6500 33880 6502
rect 33936 6500 33960 6502
rect 34016 6500 34040 6502
rect 34096 6500 34102 6502
rect 33794 6491 34102 6500
rect 33600 6112 33652 6118
rect 33600 6054 33652 6060
rect 33140 5636 33192 5642
rect 33140 5578 33192 5584
rect 33152 4826 33180 5578
rect 33508 5568 33560 5574
rect 33508 5510 33560 5516
rect 33324 5092 33376 5098
rect 33324 5034 33376 5040
rect 32772 4820 32824 4826
rect 32772 4762 32824 4768
rect 33140 4820 33192 4826
rect 33140 4762 33192 4768
rect 33232 4820 33284 4826
rect 33232 4762 33284 4768
rect 32680 4208 32732 4214
rect 32680 4150 32732 4156
rect 32864 4208 32916 4214
rect 32864 4150 32916 4156
rect 32588 3528 32640 3534
rect 32588 3470 32640 3476
rect 32876 3194 32904 4150
rect 33244 3738 33272 4762
rect 33336 4622 33364 5034
rect 33324 4616 33376 4622
rect 33324 4558 33376 4564
rect 33416 4548 33468 4554
rect 33416 4490 33468 4496
rect 33428 4282 33456 4490
rect 33520 4486 33548 5510
rect 33612 4554 33640 6054
rect 33692 5772 33744 5778
rect 33692 5714 33744 5720
rect 33704 4758 33732 5714
rect 33794 5468 34102 5477
rect 33794 5466 33800 5468
rect 33856 5466 33880 5468
rect 33936 5466 33960 5468
rect 34016 5466 34040 5468
rect 34096 5466 34102 5468
rect 33856 5414 33858 5466
rect 34038 5414 34040 5466
rect 33794 5412 33800 5414
rect 33856 5412 33880 5414
rect 33936 5412 33960 5414
rect 34016 5412 34040 5414
rect 34096 5412 34102 5414
rect 33794 5403 34102 5412
rect 33692 4752 33744 4758
rect 33692 4694 33744 4700
rect 33600 4548 33652 4554
rect 33600 4490 33652 4496
rect 33508 4480 33560 4486
rect 33508 4422 33560 4428
rect 33794 4380 34102 4389
rect 33794 4378 33800 4380
rect 33856 4378 33880 4380
rect 33936 4378 33960 4380
rect 34016 4378 34040 4380
rect 34096 4378 34102 4380
rect 33856 4326 33858 4378
rect 34038 4326 34040 4378
rect 33794 4324 33800 4326
rect 33856 4324 33880 4326
rect 33936 4324 33960 4326
rect 34016 4324 34040 4326
rect 34096 4324 34102 4326
rect 33794 4315 34102 4324
rect 33416 4276 33468 4282
rect 33416 4218 33468 4224
rect 33232 3732 33284 3738
rect 33232 3674 33284 3680
rect 33508 3392 33560 3398
rect 33508 3334 33560 3340
rect 32864 3188 32916 3194
rect 32864 3130 32916 3136
rect 32312 2304 32364 2310
rect 32312 2246 32364 2252
rect 33520 800 33548 3334
rect 33794 3292 34102 3301
rect 33794 3290 33800 3292
rect 33856 3290 33880 3292
rect 33936 3290 33960 3292
rect 34016 3290 34040 3292
rect 34096 3290 34102 3292
rect 33856 3238 33858 3290
rect 34038 3238 34040 3290
rect 33794 3236 33800 3238
rect 33856 3236 33880 3238
rect 33936 3236 33960 3238
rect 34016 3236 34040 3238
rect 34096 3236 34102 3238
rect 33794 3227 34102 3236
rect 34164 3194 34192 9880
rect 34256 9518 34284 12242
rect 34704 11892 34756 11898
rect 34704 11834 34756 11840
rect 34612 11756 34664 11762
rect 34612 11698 34664 11704
rect 34624 11218 34652 11698
rect 34612 11212 34664 11218
rect 34612 11154 34664 11160
rect 34520 10056 34572 10062
rect 34520 9998 34572 10004
rect 34532 9518 34560 9998
rect 34244 9512 34296 9518
rect 34244 9454 34296 9460
rect 34520 9512 34572 9518
rect 34716 9466 34744 11834
rect 36556 11762 36584 12242
rect 37016 12238 37044 12718
rect 37004 12232 37056 12238
rect 37004 12174 37056 12180
rect 36544 11756 36596 11762
rect 36544 11698 36596 11704
rect 37016 11218 37044 12174
rect 37188 12096 37240 12102
rect 37240 12044 37320 12050
rect 37188 12038 37320 12044
rect 37200 12022 37320 12038
rect 37292 11558 37320 12022
rect 37568 11898 37596 12786
rect 37660 12434 37688 13262
rect 37740 12436 37792 12442
rect 37660 12406 37740 12434
rect 37740 12378 37792 12384
rect 37556 11892 37608 11898
rect 37556 11834 37608 11840
rect 37648 11824 37700 11830
rect 37648 11766 37700 11772
rect 37280 11552 37332 11558
rect 37280 11494 37332 11500
rect 37556 11552 37608 11558
rect 37556 11494 37608 11500
rect 37464 11280 37516 11286
rect 37464 11222 37516 11228
rect 37004 11212 37056 11218
rect 37004 11154 37056 11160
rect 34980 11144 35032 11150
rect 34980 11086 35032 11092
rect 34992 10606 35020 11086
rect 35624 11076 35676 11082
rect 35624 11018 35676 11024
rect 34980 10600 35032 10606
rect 34980 10542 35032 10548
rect 35636 10266 35664 11018
rect 36728 11008 36780 11014
rect 36728 10950 36780 10956
rect 36740 10849 36768 10950
rect 36726 10840 36782 10849
rect 37016 10810 37044 11154
rect 37186 11112 37242 11121
rect 37186 11047 37188 11056
rect 37240 11047 37242 11056
rect 37188 11018 37240 11024
rect 36726 10775 36782 10784
rect 37004 10804 37056 10810
rect 37004 10746 37056 10752
rect 35808 10668 35860 10674
rect 35808 10610 35860 10616
rect 35992 10668 36044 10674
rect 35992 10610 36044 10616
rect 35820 10266 35848 10610
rect 35624 10260 35676 10266
rect 35624 10202 35676 10208
rect 35808 10260 35860 10266
rect 35808 10202 35860 10208
rect 34796 10056 34848 10062
rect 34796 9998 34848 10004
rect 34520 9454 34572 9460
rect 34428 9376 34480 9382
rect 34428 9318 34480 9324
rect 34440 8906 34468 9318
rect 34428 8900 34480 8906
rect 34428 8842 34480 8848
rect 34532 8838 34560 9454
rect 34624 9438 34744 9466
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34624 8294 34652 9438
rect 34808 9382 34836 9998
rect 35072 9920 35124 9926
rect 35072 9862 35124 9868
rect 35084 9722 35112 9862
rect 34888 9716 34940 9722
rect 34888 9658 34940 9664
rect 35072 9716 35124 9722
rect 35072 9658 35124 9664
rect 34704 9376 34756 9382
rect 34704 9318 34756 9324
rect 34796 9376 34848 9382
rect 34796 9318 34848 9324
rect 34716 8974 34744 9318
rect 34704 8968 34756 8974
rect 34704 8910 34756 8916
rect 34704 8832 34756 8838
rect 34704 8774 34756 8780
rect 34716 8498 34744 8774
rect 34808 8634 34836 9318
rect 34900 9110 34928 9658
rect 35084 9178 35112 9658
rect 35808 9580 35860 9586
rect 35808 9522 35860 9528
rect 35900 9580 35952 9586
rect 35900 9522 35952 9528
rect 35820 9450 35848 9522
rect 35808 9444 35860 9450
rect 35808 9386 35860 9392
rect 35072 9172 35124 9178
rect 35072 9114 35124 9120
rect 34888 9104 34940 9110
rect 34888 9046 34940 9052
rect 35912 9042 35940 9522
rect 34980 9036 35032 9042
rect 34980 8978 35032 8984
rect 35900 9036 35952 9042
rect 35900 8978 35952 8984
rect 34888 8968 34940 8974
rect 34888 8910 34940 8916
rect 34900 8634 34928 8910
rect 34796 8628 34848 8634
rect 34796 8570 34848 8576
rect 34888 8628 34940 8634
rect 34888 8570 34940 8576
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 34992 8362 35020 8978
rect 34980 8356 35032 8362
rect 34980 8298 35032 8304
rect 34612 8288 34664 8294
rect 34612 8230 34664 8236
rect 34624 7886 34652 8230
rect 34612 7880 34664 7886
rect 34612 7822 34664 7828
rect 34704 7744 34756 7750
rect 34704 7686 34756 7692
rect 34716 7546 34744 7686
rect 34704 7540 34756 7546
rect 34704 7482 34756 7488
rect 35808 7472 35860 7478
rect 35808 7414 35860 7420
rect 35348 7336 35400 7342
rect 35348 7278 35400 7284
rect 34796 7200 34848 7206
rect 34796 7142 34848 7148
rect 34520 6316 34572 6322
rect 34520 6258 34572 6264
rect 34532 5914 34560 6258
rect 34704 6248 34756 6254
rect 34704 6190 34756 6196
rect 34716 5914 34744 6190
rect 34520 5908 34572 5914
rect 34520 5850 34572 5856
rect 34704 5908 34756 5914
rect 34704 5850 34756 5856
rect 34808 4622 34836 7142
rect 35360 5914 35388 7278
rect 35820 6458 35848 7414
rect 35808 6452 35860 6458
rect 35808 6394 35860 6400
rect 35716 6316 35768 6322
rect 35716 6258 35768 6264
rect 35348 5908 35400 5914
rect 35348 5850 35400 5856
rect 35624 5704 35676 5710
rect 35624 5646 35676 5652
rect 35440 5568 35492 5574
rect 35440 5510 35492 5516
rect 35452 5166 35480 5510
rect 35440 5160 35492 5166
rect 35440 5102 35492 5108
rect 35636 4826 35664 5646
rect 35728 5234 35756 6258
rect 35716 5228 35768 5234
rect 35716 5170 35768 5176
rect 35624 4820 35676 4826
rect 35624 4762 35676 4768
rect 34796 4616 34848 4622
rect 34796 4558 34848 4564
rect 34152 3188 34204 3194
rect 34152 3130 34204 3136
rect 35532 2848 35584 2854
rect 35532 2790 35584 2796
rect 35544 2446 35572 2790
rect 36004 2650 36032 10610
rect 37476 10606 37504 11222
rect 37568 11150 37596 11494
rect 37556 11144 37608 11150
rect 37556 11086 37608 11092
rect 36544 10600 36596 10606
rect 37464 10600 37516 10606
rect 36544 10542 36596 10548
rect 37278 10568 37334 10577
rect 36176 10056 36228 10062
rect 36176 9998 36228 10004
rect 36188 8537 36216 9998
rect 36556 9994 36584 10542
rect 37464 10542 37516 10548
rect 37278 10503 37280 10512
rect 37332 10503 37334 10512
rect 37372 10532 37424 10538
rect 37280 10474 37332 10480
rect 37372 10474 37424 10480
rect 37384 10441 37412 10474
rect 37370 10432 37426 10441
rect 37370 10367 37426 10376
rect 37568 10198 37596 11086
rect 37660 10606 37688 11766
rect 37752 11762 37780 12378
rect 38016 12368 38068 12374
rect 38016 12310 38068 12316
rect 37740 11756 37792 11762
rect 37740 11698 37792 11704
rect 38028 11694 38056 12310
rect 38304 12102 38332 13262
rect 38396 12986 38424 13262
rect 38476 13252 38528 13258
rect 38476 13194 38528 13200
rect 38384 12980 38436 12986
rect 38384 12922 38436 12928
rect 38292 12096 38344 12102
rect 38292 12038 38344 12044
rect 38488 11914 38516 13194
rect 38568 13184 38620 13190
rect 38568 13126 38620 13132
rect 38580 12714 38608 13126
rect 38568 12708 38620 12714
rect 38568 12650 38620 12656
rect 38304 11886 38516 11914
rect 38106 11792 38162 11801
rect 38304 11762 38332 11886
rect 38580 11830 38608 12650
rect 38568 11824 38620 11830
rect 38568 11766 38620 11772
rect 38106 11727 38162 11736
rect 38292 11756 38344 11762
rect 38120 11694 38148 11727
rect 38292 11698 38344 11704
rect 38476 11756 38528 11762
rect 38476 11698 38528 11704
rect 38016 11688 38068 11694
rect 38016 11630 38068 11636
rect 38108 11688 38160 11694
rect 38108 11630 38160 11636
rect 38488 11558 38516 11698
rect 38476 11552 38528 11558
rect 38476 11494 38528 11500
rect 37924 11212 37976 11218
rect 37924 11154 37976 11160
rect 37740 11076 37792 11082
rect 37740 11018 37792 11024
rect 37648 10600 37700 10606
rect 37648 10542 37700 10548
rect 37556 10192 37608 10198
rect 37556 10134 37608 10140
rect 37660 9994 37688 10542
rect 37752 10441 37780 11018
rect 37832 11008 37884 11014
rect 37832 10950 37884 10956
rect 37844 10577 37872 10950
rect 37830 10568 37886 10577
rect 37830 10503 37886 10512
rect 37738 10432 37794 10441
rect 37738 10367 37794 10376
rect 37936 10130 37964 11154
rect 38290 10840 38346 10849
rect 38290 10775 38346 10784
rect 38304 10742 38332 10775
rect 38292 10736 38344 10742
rect 38292 10678 38344 10684
rect 38488 10606 38516 11494
rect 38580 11150 38608 11766
rect 38948 11762 38976 13330
rect 39672 13320 39724 13326
rect 39672 13262 39724 13268
rect 39120 12980 39172 12986
rect 39120 12922 39172 12928
rect 39028 12232 39080 12238
rect 39028 12174 39080 12180
rect 39040 11898 39068 12174
rect 39028 11892 39080 11898
rect 39028 11834 39080 11840
rect 38936 11756 38988 11762
rect 38936 11698 38988 11704
rect 39028 11756 39080 11762
rect 39028 11698 39080 11704
rect 39040 11558 39068 11698
rect 39028 11552 39080 11558
rect 39028 11494 39080 11500
rect 38568 11144 38620 11150
rect 38660 11144 38712 11150
rect 38568 11086 38620 11092
rect 38658 11112 38660 11121
rect 38712 11112 38714 11121
rect 38658 11047 38714 11056
rect 39132 10674 39160 12922
rect 39684 12646 39712 13262
rect 39764 12912 39816 12918
rect 39764 12854 39816 12860
rect 39672 12640 39724 12646
rect 39672 12582 39724 12588
rect 39268 12540 39576 12549
rect 39268 12538 39274 12540
rect 39330 12538 39354 12540
rect 39410 12538 39434 12540
rect 39490 12538 39514 12540
rect 39570 12538 39576 12540
rect 39330 12486 39332 12538
rect 39512 12486 39514 12538
rect 39268 12484 39274 12486
rect 39330 12484 39354 12486
rect 39410 12484 39434 12486
rect 39490 12484 39514 12486
rect 39570 12484 39576 12486
rect 39268 12475 39576 12484
rect 39684 12238 39712 12582
rect 39776 12434 39804 12854
rect 40052 12782 40080 16526
rect 40696 16454 40724 17138
rect 42524 17060 42576 17066
rect 42524 17002 42576 17008
rect 40684 16448 40736 16454
rect 40684 16390 40736 16396
rect 40960 13456 41012 13462
rect 40960 13398 41012 13404
rect 40224 13184 40276 13190
rect 40224 13126 40276 13132
rect 40500 13184 40552 13190
rect 40500 13126 40552 13132
rect 40040 12776 40092 12782
rect 40040 12718 40092 12724
rect 39776 12406 39988 12434
rect 39856 12368 39908 12374
rect 39856 12310 39908 12316
rect 39304 12232 39356 12238
rect 39304 12174 39356 12180
rect 39672 12232 39724 12238
rect 39672 12174 39724 12180
rect 39316 12102 39344 12174
rect 39304 12096 39356 12102
rect 39304 12038 39356 12044
rect 39316 11830 39344 12038
rect 39304 11824 39356 11830
rect 39304 11766 39356 11772
rect 39268 11452 39576 11461
rect 39268 11450 39274 11452
rect 39330 11450 39354 11452
rect 39410 11450 39434 11452
rect 39490 11450 39514 11452
rect 39570 11450 39576 11452
rect 39330 11398 39332 11450
rect 39512 11398 39514 11450
rect 39268 11396 39274 11398
rect 39330 11396 39354 11398
rect 39410 11396 39434 11398
rect 39490 11396 39514 11398
rect 39570 11396 39576 11398
rect 39268 11387 39576 11396
rect 39684 10810 39712 12174
rect 39868 12170 39896 12310
rect 39856 12164 39908 12170
rect 39856 12106 39908 12112
rect 39764 11756 39816 11762
rect 39764 11698 39816 11704
rect 39776 11082 39804 11698
rect 39764 11076 39816 11082
rect 39764 11018 39816 11024
rect 39672 10804 39724 10810
rect 39672 10746 39724 10752
rect 39120 10668 39172 10674
rect 39120 10610 39172 10616
rect 38476 10600 38528 10606
rect 38476 10542 38528 10548
rect 37924 10124 37976 10130
rect 37924 10066 37976 10072
rect 38476 10056 38528 10062
rect 38476 9998 38528 10004
rect 36544 9988 36596 9994
rect 36544 9930 36596 9936
rect 37648 9988 37700 9994
rect 37648 9930 37700 9936
rect 36556 9586 36584 9930
rect 36544 9580 36596 9586
rect 36544 9522 36596 9528
rect 38488 9450 38516 9998
rect 38844 9988 38896 9994
rect 38844 9930 38896 9936
rect 38660 9648 38712 9654
rect 38660 9590 38712 9596
rect 38568 9580 38620 9586
rect 38568 9522 38620 9528
rect 38476 9444 38528 9450
rect 38476 9386 38528 9392
rect 38200 9172 38252 9178
rect 38200 9114 38252 9120
rect 36174 8528 36230 8537
rect 38212 8498 38240 9114
rect 38488 8498 38516 9386
rect 38580 8974 38608 9522
rect 38568 8968 38620 8974
rect 38568 8910 38620 8916
rect 38672 8906 38700 9590
rect 38752 9580 38804 9586
rect 38752 9522 38804 9528
rect 38660 8900 38712 8906
rect 38660 8842 38712 8848
rect 36174 8463 36230 8472
rect 37372 8492 37424 8498
rect 37372 8434 37424 8440
rect 38200 8492 38252 8498
rect 38200 8434 38252 8440
rect 38476 8492 38528 8498
rect 38476 8434 38528 8440
rect 37384 2650 37412 8434
rect 38764 8362 38792 9522
rect 38856 9178 38884 9930
rect 39028 9920 39080 9926
rect 39028 9862 39080 9868
rect 38936 9512 38988 9518
rect 38936 9454 38988 9460
rect 38844 9172 38896 9178
rect 38844 9114 38896 9120
rect 38948 8634 38976 9454
rect 39040 8974 39068 9862
rect 39132 9722 39160 10610
rect 39268 10364 39576 10373
rect 39268 10362 39274 10364
rect 39330 10362 39354 10364
rect 39410 10362 39434 10364
rect 39490 10362 39514 10364
rect 39570 10362 39576 10364
rect 39330 10310 39332 10362
rect 39512 10310 39514 10362
rect 39268 10308 39274 10310
rect 39330 10308 39354 10310
rect 39410 10308 39434 10310
rect 39490 10308 39514 10310
rect 39570 10308 39576 10310
rect 39268 10299 39576 10308
rect 39672 10260 39724 10266
rect 39672 10202 39724 10208
rect 39120 9716 39172 9722
rect 39120 9658 39172 9664
rect 39684 9654 39712 10202
rect 39672 9648 39724 9654
rect 39670 9616 39672 9625
rect 39724 9616 39726 9625
rect 39670 9551 39726 9560
rect 39268 9276 39576 9285
rect 39268 9274 39274 9276
rect 39330 9274 39354 9276
rect 39410 9274 39434 9276
rect 39490 9274 39514 9276
rect 39570 9274 39576 9276
rect 39330 9222 39332 9274
rect 39512 9222 39514 9274
rect 39268 9220 39274 9222
rect 39330 9220 39354 9222
rect 39410 9220 39434 9222
rect 39490 9220 39514 9222
rect 39570 9220 39576 9222
rect 39268 9211 39576 9220
rect 39120 9104 39172 9110
rect 39120 9046 39172 9052
rect 39210 9072 39266 9081
rect 39028 8968 39080 8974
rect 39028 8910 39080 8916
rect 38936 8628 38988 8634
rect 38936 8570 38988 8576
rect 38936 8492 38988 8498
rect 38936 8434 38988 8440
rect 38752 8356 38804 8362
rect 38752 8298 38804 8304
rect 38948 7954 38976 8434
rect 38936 7948 38988 7954
rect 38936 7890 38988 7896
rect 39132 7886 39160 9046
rect 39210 9007 39266 9016
rect 39580 9036 39632 9042
rect 39224 8838 39252 9007
rect 39580 8978 39632 8984
rect 39212 8832 39264 8838
rect 39212 8774 39264 8780
rect 39304 8832 39356 8838
rect 39304 8774 39356 8780
rect 39316 8498 39344 8774
rect 39592 8498 39620 8978
rect 39684 8974 39712 9551
rect 39868 9518 39896 12106
rect 39960 11898 39988 12406
rect 39948 11892 40000 11898
rect 39948 11834 40000 11840
rect 39960 11762 39988 11834
rect 40132 11824 40184 11830
rect 40132 11766 40184 11772
rect 39948 11756 40000 11762
rect 39948 11698 40000 11704
rect 39960 11286 39988 11698
rect 39948 11280 40000 11286
rect 39948 11222 40000 11228
rect 40144 11014 40172 11766
rect 40236 11150 40264 13126
rect 40512 12442 40540 13126
rect 40592 12844 40644 12850
rect 40592 12786 40644 12792
rect 40500 12436 40552 12442
rect 40500 12378 40552 12384
rect 40408 12368 40460 12374
rect 40328 12328 40408 12356
rect 40328 12170 40356 12328
rect 40408 12310 40460 12316
rect 40316 12164 40368 12170
rect 40316 12106 40368 12112
rect 40512 11830 40540 12378
rect 40604 12306 40632 12786
rect 40592 12300 40644 12306
rect 40592 12242 40644 12248
rect 40776 12164 40828 12170
rect 40776 12106 40828 12112
rect 40500 11824 40552 11830
rect 40500 11766 40552 11772
rect 40788 11762 40816 12106
rect 40408 11756 40460 11762
rect 40408 11698 40460 11704
rect 40592 11756 40644 11762
rect 40592 11698 40644 11704
rect 40776 11756 40828 11762
rect 40776 11698 40828 11704
rect 40316 11620 40368 11626
rect 40316 11562 40368 11568
rect 40328 11529 40356 11562
rect 40314 11520 40370 11529
rect 40314 11455 40370 11464
rect 40420 11234 40448 11698
rect 40500 11552 40552 11558
rect 40500 11494 40552 11500
rect 40328 11206 40448 11234
rect 40224 11144 40276 11150
rect 40224 11086 40276 11092
rect 40132 11008 40184 11014
rect 40132 10950 40184 10956
rect 40328 10418 40356 11206
rect 40408 11144 40460 11150
rect 40408 11086 40460 11092
rect 40144 10390 40356 10418
rect 40144 10266 40172 10390
rect 40132 10260 40184 10266
rect 40132 10202 40184 10208
rect 40316 10260 40368 10266
rect 40316 10202 40368 10208
rect 40328 10169 40356 10202
rect 40314 10160 40370 10169
rect 40420 10146 40448 11086
rect 40512 10674 40540 11494
rect 40604 11354 40632 11698
rect 40592 11348 40644 11354
rect 40592 11290 40644 11296
rect 40972 11150 41000 13398
rect 41972 13252 42024 13258
rect 41972 13194 42024 13200
rect 41984 12646 42012 13194
rect 41972 12640 42024 12646
rect 41972 12582 42024 12588
rect 41052 12164 41104 12170
rect 41052 12106 41104 12112
rect 41064 11354 41092 12106
rect 41604 11892 41656 11898
rect 41604 11834 41656 11840
rect 41512 11824 41564 11830
rect 41512 11766 41564 11772
rect 41328 11552 41380 11558
rect 41328 11494 41380 11500
rect 41052 11348 41104 11354
rect 41052 11290 41104 11296
rect 41340 11218 41368 11494
rect 41524 11218 41552 11766
rect 41328 11212 41380 11218
rect 41328 11154 41380 11160
rect 41512 11212 41564 11218
rect 41512 11154 41564 11160
rect 40960 11144 41012 11150
rect 40960 11086 41012 11092
rect 41420 11144 41472 11150
rect 41420 11086 41472 11092
rect 41052 11008 41104 11014
rect 41052 10950 41104 10956
rect 40500 10668 40552 10674
rect 40500 10610 40552 10616
rect 41064 10606 41092 10950
rect 41432 10810 41460 11086
rect 41512 11076 41564 11082
rect 41512 11018 41564 11024
rect 41420 10804 41472 10810
rect 41420 10746 41472 10752
rect 41052 10600 41104 10606
rect 41052 10542 41104 10548
rect 40500 10532 40552 10538
rect 40500 10474 40552 10480
rect 41236 10532 41288 10538
rect 41236 10474 41288 10480
rect 40512 10266 40540 10474
rect 40592 10464 40644 10470
rect 40592 10406 40644 10412
rect 40776 10464 40828 10470
rect 40776 10406 40828 10412
rect 40604 10266 40632 10406
rect 40500 10260 40552 10266
rect 40500 10202 40552 10208
rect 40592 10260 40644 10266
rect 40592 10202 40644 10208
rect 40370 10118 40448 10146
rect 40314 10095 40370 10104
rect 40132 10056 40184 10062
rect 40316 10056 40368 10062
rect 40132 9998 40184 10004
rect 40314 10024 40316 10033
rect 40368 10024 40370 10033
rect 40144 9586 40172 9998
rect 40314 9959 40370 9968
rect 40328 9636 40356 9959
rect 40236 9608 40356 9636
rect 40132 9580 40184 9586
rect 40132 9522 40184 9528
rect 39856 9512 39908 9518
rect 39856 9454 39908 9460
rect 40144 9382 40172 9522
rect 40236 9450 40264 9608
rect 40224 9444 40276 9450
rect 40224 9386 40276 9392
rect 40132 9376 40184 9382
rect 40132 9318 40184 9324
rect 40132 9172 40184 9178
rect 40132 9114 40184 9120
rect 39856 9104 39908 9110
rect 39856 9046 39908 9052
rect 39672 8968 39724 8974
rect 39672 8910 39724 8916
rect 39868 8566 39896 9046
rect 40040 8968 40092 8974
rect 40040 8910 40092 8916
rect 39856 8560 39908 8566
rect 39856 8502 39908 8508
rect 39304 8492 39356 8498
rect 39304 8434 39356 8440
rect 39580 8492 39632 8498
rect 39580 8434 39632 8440
rect 39268 8188 39576 8197
rect 39268 8186 39274 8188
rect 39330 8186 39354 8188
rect 39410 8186 39434 8188
rect 39490 8186 39514 8188
rect 39570 8186 39576 8188
rect 39330 8134 39332 8186
rect 39512 8134 39514 8186
rect 39268 8132 39274 8134
rect 39330 8132 39354 8134
rect 39410 8132 39434 8134
rect 39490 8132 39514 8134
rect 39570 8132 39576 8134
rect 39268 8123 39576 8132
rect 39868 7954 39896 8502
rect 40052 8090 40080 8910
rect 40040 8084 40092 8090
rect 40040 8026 40092 8032
rect 39856 7948 39908 7954
rect 39856 7890 39908 7896
rect 39120 7880 39172 7886
rect 39120 7822 39172 7828
rect 39396 7880 39448 7886
rect 39396 7822 39448 7828
rect 39408 7410 39436 7822
rect 39856 7812 39908 7818
rect 39856 7754 39908 7760
rect 39868 7546 39896 7754
rect 39856 7540 39908 7546
rect 39856 7482 39908 7488
rect 39396 7404 39448 7410
rect 39396 7346 39448 7352
rect 39948 7404 40000 7410
rect 39948 7346 40000 7352
rect 39268 7100 39576 7109
rect 39268 7098 39274 7100
rect 39330 7098 39354 7100
rect 39410 7098 39434 7100
rect 39490 7098 39514 7100
rect 39570 7098 39576 7100
rect 39330 7046 39332 7098
rect 39512 7046 39514 7098
rect 39268 7044 39274 7046
rect 39330 7044 39354 7046
rect 39410 7044 39434 7046
rect 39490 7044 39514 7046
rect 39570 7044 39576 7046
rect 39268 7035 39576 7044
rect 39960 6866 39988 7346
rect 39948 6860 40000 6866
rect 39948 6802 40000 6808
rect 40144 6798 40172 9114
rect 40236 9081 40264 9386
rect 40222 9072 40278 9081
rect 40222 9007 40278 9016
rect 40236 8906 40264 9007
rect 40224 8900 40276 8906
rect 40224 8842 40276 8848
rect 40420 8430 40448 10118
rect 40684 10056 40736 10062
rect 40684 9998 40736 10004
rect 40696 9897 40724 9998
rect 40682 9888 40738 9897
rect 40682 9823 40738 9832
rect 40788 9722 40816 10406
rect 41144 10056 41196 10062
rect 41142 10024 41144 10033
rect 41196 10024 41198 10033
rect 41142 9959 41198 9968
rect 40868 9920 40920 9926
rect 40868 9862 40920 9868
rect 40776 9716 40828 9722
rect 40776 9658 40828 9664
rect 40880 9382 40908 9862
rect 41248 9722 41276 10474
rect 41326 10160 41382 10169
rect 41326 10095 41382 10104
rect 41340 10062 41368 10095
rect 41524 10062 41552 11018
rect 41616 10674 41644 11834
rect 41984 11762 42012 12582
rect 42432 12096 42484 12102
rect 42432 12038 42484 12044
rect 41972 11756 42024 11762
rect 41972 11698 42024 11704
rect 41984 11150 42012 11698
rect 42444 11694 42472 12038
rect 42432 11688 42484 11694
rect 42432 11630 42484 11636
rect 42062 11520 42118 11529
rect 42062 11455 42118 11464
rect 42076 11354 42104 11455
rect 42064 11348 42116 11354
rect 42064 11290 42116 11296
rect 42444 11150 42472 11630
rect 41972 11144 42024 11150
rect 41972 11086 42024 11092
rect 42432 11144 42484 11150
rect 42432 11086 42484 11092
rect 42536 11082 42564 17002
rect 43456 16794 43484 19071
rect 43824 16794 43852 19200
rect 44086 17776 44142 17785
rect 44086 17711 44142 17720
rect 44100 17338 44128 17711
rect 44742 17436 45050 17445
rect 44742 17434 44748 17436
rect 44804 17434 44828 17436
rect 44884 17434 44908 17436
rect 44964 17434 44988 17436
rect 45044 17434 45050 17436
rect 44804 17382 44806 17434
rect 44986 17382 44988 17434
rect 44742 17380 44748 17382
rect 44804 17380 44828 17382
rect 44884 17380 44908 17382
rect 44964 17380 44988 17382
rect 45044 17380 45050 17382
rect 44742 17371 45050 17380
rect 44088 17332 44140 17338
rect 44088 17274 44140 17280
rect 43904 17196 43956 17202
rect 43904 17138 43956 17144
rect 43444 16788 43496 16794
rect 43444 16730 43496 16736
rect 43812 16788 43864 16794
rect 43812 16730 43864 16736
rect 43916 15366 43944 17138
rect 45112 17134 45140 19200
rect 45100 17128 45152 17134
rect 45100 17070 45152 17076
rect 44742 16348 45050 16357
rect 44742 16346 44748 16348
rect 44804 16346 44828 16348
rect 44884 16346 44908 16348
rect 44964 16346 44988 16348
rect 45044 16346 45050 16348
rect 44804 16294 44806 16346
rect 44986 16294 44988 16346
rect 44742 16292 44748 16294
rect 44804 16292 44828 16294
rect 44884 16292 44908 16294
rect 44964 16292 44988 16294
rect 45044 16292 45050 16294
rect 44742 16283 45050 16292
rect 44180 15904 44232 15910
rect 44180 15846 44232 15852
rect 44192 15745 44220 15846
rect 44178 15736 44234 15745
rect 44178 15671 44234 15680
rect 43904 15360 43956 15366
rect 43904 15302 43956 15308
rect 44742 15260 45050 15269
rect 44742 15258 44748 15260
rect 44804 15258 44828 15260
rect 44884 15258 44908 15260
rect 44964 15258 44988 15260
rect 45044 15258 45050 15260
rect 44804 15206 44806 15258
rect 44986 15206 44988 15258
rect 44742 15204 44748 15206
rect 44804 15204 44828 15206
rect 44884 15204 44908 15206
rect 44964 15204 44988 15206
rect 45044 15204 45050 15206
rect 44742 15195 45050 15204
rect 42984 14408 43036 14414
rect 42984 14350 43036 14356
rect 44086 14376 44142 14385
rect 42996 14006 43024 14350
rect 44086 14311 44142 14320
rect 44100 14278 44128 14311
rect 44088 14272 44140 14278
rect 44088 14214 44140 14220
rect 44742 14172 45050 14181
rect 44742 14170 44748 14172
rect 44804 14170 44828 14172
rect 44884 14170 44908 14172
rect 44964 14170 44988 14172
rect 45044 14170 45050 14172
rect 44804 14118 44806 14170
rect 44986 14118 44988 14170
rect 44742 14116 44748 14118
rect 44804 14116 44828 14118
rect 44884 14116 44908 14118
rect 44964 14116 44988 14118
rect 45044 14116 45050 14118
rect 44742 14107 45050 14116
rect 42984 14000 43036 14006
rect 42984 13942 43036 13948
rect 42616 13456 42668 13462
rect 42616 13398 42668 13404
rect 42628 12306 42656 13398
rect 44742 13084 45050 13093
rect 44742 13082 44748 13084
rect 44804 13082 44828 13084
rect 44884 13082 44908 13084
rect 44964 13082 44988 13084
rect 45044 13082 45050 13084
rect 44804 13030 44806 13082
rect 44986 13030 44988 13082
rect 44742 13028 44748 13030
rect 44804 13028 44828 13030
rect 44884 13028 44908 13030
rect 44964 13028 44988 13030
rect 45044 13028 45050 13030
rect 44742 13019 45050 13028
rect 42708 12844 42760 12850
rect 42708 12786 42760 12792
rect 42720 12442 42748 12786
rect 44088 12640 44140 12646
rect 44088 12582 44140 12588
rect 42708 12436 42760 12442
rect 42708 12378 42760 12384
rect 44100 12345 44128 12582
rect 44086 12336 44142 12345
rect 42616 12300 42668 12306
rect 44086 12271 44142 12280
rect 42616 12242 42668 12248
rect 44742 11996 45050 12005
rect 44742 11994 44748 11996
rect 44804 11994 44828 11996
rect 44884 11994 44908 11996
rect 44964 11994 44988 11996
rect 45044 11994 45050 11996
rect 44804 11942 44806 11994
rect 44986 11942 44988 11994
rect 44742 11940 44748 11942
rect 44804 11940 44828 11942
rect 44884 11940 44908 11942
rect 44964 11940 44988 11942
rect 45044 11940 45050 11942
rect 44742 11931 45050 11940
rect 42708 11688 42760 11694
rect 42708 11630 42760 11636
rect 42720 11218 42748 11630
rect 42708 11212 42760 11218
rect 42708 11154 42760 11160
rect 42524 11076 42576 11082
rect 42524 11018 42576 11024
rect 42892 11008 42944 11014
rect 42892 10950 42944 10956
rect 43536 11008 43588 11014
rect 43536 10950 43588 10956
rect 42904 10742 42932 10950
rect 42892 10736 42944 10742
rect 42892 10678 42944 10684
rect 43548 10674 43576 10950
rect 44742 10908 45050 10917
rect 44742 10906 44748 10908
rect 44804 10906 44828 10908
rect 44884 10906 44908 10908
rect 44964 10906 44988 10908
rect 45044 10906 45050 10908
rect 44804 10854 44806 10906
rect 44986 10854 44988 10906
rect 44742 10852 44748 10854
rect 44804 10852 44828 10854
rect 44884 10852 44908 10854
rect 44964 10852 44988 10854
rect 45044 10852 45050 10854
rect 44742 10843 45050 10852
rect 44178 10704 44234 10713
rect 41604 10668 41656 10674
rect 41604 10610 41656 10616
rect 42800 10668 42852 10674
rect 42800 10610 42852 10616
rect 43536 10668 43588 10674
rect 44178 10639 44180 10648
rect 43536 10610 43588 10616
rect 44232 10639 44234 10648
rect 44180 10610 44232 10616
rect 42708 10464 42760 10470
rect 42708 10406 42760 10412
rect 41972 10124 42024 10130
rect 41972 10066 42024 10072
rect 41328 10056 41380 10062
rect 41328 9998 41380 10004
rect 41512 10056 41564 10062
rect 41512 9998 41564 10004
rect 41984 9994 42012 10066
rect 42064 10056 42116 10062
rect 42064 9998 42116 10004
rect 42340 10056 42392 10062
rect 42340 9998 42392 10004
rect 41972 9988 42024 9994
rect 41972 9930 42024 9936
rect 41694 9888 41750 9897
rect 41694 9823 41750 9832
rect 41236 9716 41288 9722
rect 41236 9658 41288 9664
rect 40958 9616 41014 9625
rect 41328 9580 41380 9586
rect 41014 9560 41328 9568
rect 40958 9551 40960 9560
rect 41012 9540 41328 9560
rect 40960 9522 41012 9528
rect 41328 9522 41380 9528
rect 41708 9382 41736 9823
rect 42076 9518 42104 9998
rect 42156 9920 42208 9926
rect 42156 9862 42208 9868
rect 42064 9512 42116 9518
rect 42064 9454 42116 9460
rect 40868 9376 40920 9382
rect 40868 9318 40920 9324
rect 41512 9376 41564 9382
rect 41512 9318 41564 9324
rect 41696 9376 41748 9382
rect 41696 9318 41748 9324
rect 41524 8974 41552 9318
rect 42168 9110 42196 9862
rect 42352 9722 42380 9998
rect 42340 9716 42392 9722
rect 42340 9658 42392 9664
rect 42720 9586 42748 10406
rect 42812 10266 42840 10610
rect 43352 10600 43404 10606
rect 43352 10542 43404 10548
rect 42800 10260 42852 10266
rect 42800 10202 42852 10208
rect 43364 9654 43392 10542
rect 43444 10056 43496 10062
rect 43444 9998 43496 10004
rect 43352 9648 43404 9654
rect 43352 9590 43404 9596
rect 43456 9586 43484 9998
rect 43628 9920 43680 9926
rect 43628 9862 43680 9868
rect 43640 9586 43668 9862
rect 44742 9820 45050 9829
rect 44742 9818 44748 9820
rect 44804 9818 44828 9820
rect 44884 9818 44908 9820
rect 44964 9818 44988 9820
rect 45044 9818 45050 9820
rect 44804 9766 44806 9818
rect 44986 9766 44988 9818
rect 44742 9764 44748 9766
rect 44804 9764 44828 9766
rect 44884 9764 44908 9766
rect 44964 9764 44988 9766
rect 45044 9764 45050 9766
rect 44742 9755 45050 9764
rect 42616 9580 42668 9586
rect 42616 9522 42668 9528
rect 42708 9580 42760 9586
rect 42708 9522 42760 9528
rect 43444 9580 43496 9586
rect 43444 9522 43496 9528
rect 43628 9580 43680 9586
rect 43628 9522 43680 9528
rect 42524 9512 42576 9518
rect 42524 9454 42576 9460
rect 42156 9104 42208 9110
rect 42156 9046 42208 9052
rect 40500 8968 40552 8974
rect 40500 8910 40552 8916
rect 41512 8968 41564 8974
rect 41512 8910 41564 8916
rect 40512 8634 40540 8910
rect 40776 8900 40828 8906
rect 40776 8842 40828 8848
rect 40500 8628 40552 8634
rect 40500 8570 40552 8576
rect 40408 8424 40460 8430
rect 40328 8372 40408 8378
rect 40328 8366 40460 8372
rect 40328 8350 40448 8366
rect 40328 7410 40356 8350
rect 40408 7744 40460 7750
rect 40408 7686 40460 7692
rect 40316 7404 40368 7410
rect 40316 7346 40368 7352
rect 40420 7342 40448 7686
rect 40788 7546 40816 8842
rect 41236 8492 41288 8498
rect 41236 8434 41288 8440
rect 41144 8424 41196 8430
rect 41144 8366 41196 8372
rect 41156 7954 41184 8366
rect 41248 8090 41276 8434
rect 41524 8430 41552 8910
rect 42536 8430 42564 9454
rect 42628 9058 42656 9522
rect 43352 9444 43404 9450
rect 43352 9386 43404 9392
rect 43364 9178 43392 9386
rect 43352 9172 43404 9178
rect 43352 9114 43404 9120
rect 42628 9030 42748 9058
rect 42616 8968 42668 8974
rect 42616 8910 42668 8916
rect 41512 8424 41564 8430
rect 41512 8366 41564 8372
rect 42524 8424 42576 8430
rect 42524 8366 42576 8372
rect 41236 8084 41288 8090
rect 41236 8026 41288 8032
rect 41144 7948 41196 7954
rect 41144 7890 41196 7896
rect 41144 7744 41196 7750
rect 41144 7686 41196 7692
rect 40776 7540 40828 7546
rect 40776 7482 40828 7488
rect 41156 7410 41184 7686
rect 41524 7410 41552 8366
rect 42628 8362 42656 8910
rect 42616 8356 42668 8362
rect 42616 8298 42668 8304
rect 42628 7886 42656 8298
rect 42720 8090 42748 9030
rect 42800 8832 42852 8838
rect 42800 8774 42852 8780
rect 42812 8566 42840 8774
rect 42800 8560 42852 8566
rect 42800 8502 42852 8508
rect 43260 8492 43312 8498
rect 43260 8434 43312 8440
rect 42708 8084 42760 8090
rect 42708 8026 42760 8032
rect 41880 7880 41932 7886
rect 41880 7822 41932 7828
rect 42616 7880 42668 7886
rect 42616 7822 42668 7828
rect 40960 7404 41012 7410
rect 40960 7346 41012 7352
rect 41144 7404 41196 7410
rect 41144 7346 41196 7352
rect 41512 7404 41564 7410
rect 41512 7346 41564 7352
rect 40408 7336 40460 7342
rect 40408 7278 40460 7284
rect 40972 7002 41000 7346
rect 41892 7206 41920 7822
rect 41880 7200 41932 7206
rect 41880 7142 41932 7148
rect 40960 6996 41012 7002
rect 40960 6938 41012 6944
rect 40132 6792 40184 6798
rect 40132 6734 40184 6740
rect 39268 6012 39576 6021
rect 39268 6010 39274 6012
rect 39330 6010 39354 6012
rect 39410 6010 39434 6012
rect 39490 6010 39514 6012
rect 39570 6010 39576 6012
rect 39330 5958 39332 6010
rect 39512 5958 39514 6010
rect 39268 5956 39274 5958
rect 39330 5956 39354 5958
rect 39410 5956 39434 5958
rect 39490 5956 39514 5958
rect 39570 5956 39576 5958
rect 39268 5947 39576 5956
rect 42800 5024 42852 5030
rect 42800 4966 42852 4972
rect 39268 4924 39576 4933
rect 39268 4922 39274 4924
rect 39330 4922 39354 4924
rect 39410 4922 39434 4924
rect 39490 4922 39514 4924
rect 39570 4922 39576 4924
rect 39330 4870 39332 4922
rect 39512 4870 39514 4922
rect 39268 4868 39274 4870
rect 39330 4868 39354 4870
rect 39410 4868 39434 4870
rect 39490 4868 39514 4870
rect 39570 4868 39576 4870
rect 39268 4859 39576 4868
rect 42812 4622 42840 4966
rect 42800 4616 42852 4622
rect 42800 4558 42852 4564
rect 39268 3836 39576 3845
rect 39268 3834 39274 3836
rect 39330 3834 39354 3836
rect 39410 3834 39434 3836
rect 39490 3834 39514 3836
rect 39570 3834 39576 3836
rect 39330 3782 39332 3834
rect 39512 3782 39514 3834
rect 39268 3780 39274 3782
rect 39330 3780 39354 3782
rect 39410 3780 39434 3782
rect 39490 3780 39514 3782
rect 39570 3780 39576 3782
rect 39268 3771 39576 3780
rect 43272 3194 43300 8434
rect 43456 3194 43484 9522
rect 44178 8936 44234 8945
rect 44178 8871 44234 8880
rect 44192 8498 44220 8871
rect 44742 8732 45050 8741
rect 44742 8730 44748 8732
rect 44804 8730 44828 8732
rect 44884 8730 44908 8732
rect 44964 8730 44988 8732
rect 45044 8730 45050 8732
rect 44804 8678 44806 8730
rect 44986 8678 44988 8730
rect 44742 8676 44748 8678
rect 44804 8676 44828 8678
rect 44884 8676 44908 8678
rect 44964 8676 44988 8678
rect 45044 8676 45050 8678
rect 44742 8667 45050 8676
rect 44180 8492 44232 8498
rect 44180 8434 44232 8440
rect 44180 7880 44232 7886
rect 44178 7848 44180 7857
rect 44232 7848 44234 7857
rect 44178 7783 44234 7792
rect 44742 7644 45050 7653
rect 44742 7642 44748 7644
rect 44804 7642 44828 7644
rect 44884 7642 44908 7644
rect 44964 7642 44988 7644
rect 45044 7642 45050 7644
rect 44804 7590 44806 7642
rect 44986 7590 44988 7642
rect 44742 7588 44748 7590
rect 44804 7588 44828 7590
rect 44884 7588 44908 7590
rect 44964 7588 44988 7590
rect 45044 7588 45050 7590
rect 44742 7579 45050 7588
rect 43904 7336 43956 7342
rect 43904 7278 43956 7284
rect 43916 5710 43944 7278
rect 44742 6556 45050 6565
rect 44742 6554 44748 6556
rect 44804 6554 44828 6556
rect 44884 6554 44908 6556
rect 44964 6554 44988 6556
rect 45044 6554 45050 6556
rect 44804 6502 44806 6554
rect 44986 6502 44988 6554
rect 44742 6500 44748 6502
rect 44804 6500 44828 6502
rect 44884 6500 44908 6502
rect 44964 6500 44988 6502
rect 45044 6500 45050 6502
rect 44742 6491 45050 6500
rect 43904 5704 43956 5710
rect 43904 5646 43956 5652
rect 44088 5568 44140 5574
rect 44088 5510 44140 5516
rect 44100 5273 44128 5510
rect 44742 5468 45050 5477
rect 44742 5466 44748 5468
rect 44804 5466 44828 5468
rect 44884 5466 44908 5468
rect 44964 5466 44988 5468
rect 45044 5466 45050 5468
rect 44804 5414 44806 5466
rect 44986 5414 44988 5466
rect 44742 5412 44748 5414
rect 44804 5412 44828 5414
rect 44884 5412 44908 5414
rect 44964 5412 44988 5414
rect 45044 5412 45050 5414
rect 44742 5403 45050 5412
rect 44086 5264 44142 5273
rect 44086 5199 44142 5208
rect 44088 4480 44140 4486
rect 44088 4422 44140 4428
rect 44100 4185 44128 4422
rect 44742 4380 45050 4389
rect 44742 4378 44748 4380
rect 44804 4378 44828 4380
rect 44884 4378 44908 4380
rect 44964 4378 44988 4380
rect 45044 4378 45050 4380
rect 44804 4326 44806 4378
rect 44986 4326 44988 4378
rect 44742 4324 44748 4326
rect 44804 4324 44828 4326
rect 44884 4324 44908 4326
rect 44964 4324 44988 4326
rect 45044 4324 45050 4326
rect 44742 4315 45050 4324
rect 44086 4176 44142 4185
rect 44086 4111 44142 4120
rect 43904 3936 43956 3942
rect 43904 3878 43956 3884
rect 43260 3188 43312 3194
rect 43260 3130 43312 3136
rect 43444 3188 43496 3194
rect 43444 3130 43496 3136
rect 43812 3052 43864 3058
rect 43812 2994 43864 3000
rect 39268 2748 39576 2757
rect 39268 2746 39274 2748
rect 39330 2746 39354 2748
rect 39410 2746 39434 2748
rect 39490 2746 39514 2748
rect 39570 2746 39576 2748
rect 39330 2694 39332 2746
rect 39512 2694 39514 2746
rect 39268 2692 39274 2694
rect 39330 2692 39354 2694
rect 39410 2692 39434 2694
rect 39490 2692 39514 2694
rect 39570 2692 39576 2694
rect 39268 2683 39576 2692
rect 35992 2644 36044 2650
rect 35992 2586 36044 2592
rect 37372 2644 37424 2650
rect 37372 2586 37424 2592
rect 35532 2440 35584 2446
rect 35532 2382 35584 2388
rect 36728 2440 36780 2446
rect 36728 2382 36780 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 39948 2440 40000 2446
rect 39948 2382 40000 2388
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 33794 2204 34102 2213
rect 33794 2202 33800 2204
rect 33856 2202 33880 2204
rect 33936 2202 33960 2204
rect 34016 2202 34040 2204
rect 34096 2202 34102 2204
rect 33856 2150 33858 2202
rect 34038 2150 34040 2202
rect 33794 2148 33800 2150
rect 33856 2148 33880 2150
rect 33936 2148 33960 2150
rect 34016 2148 34040 2150
rect 34096 2148 34102 2150
rect 33794 2139 34102 2148
rect 35452 800 35480 2246
rect 36740 800 36768 2382
rect 38672 800 38700 2382
rect 39960 800 39988 2382
rect 41880 2372 41932 2378
rect 41880 2314 41932 2320
rect 41892 800 41920 2314
rect 43824 800 43852 2994
rect 43916 2446 43944 3878
rect 44180 3528 44232 3534
rect 44180 3470 44232 3476
rect 43904 2440 43956 2446
rect 43904 2382 43956 2388
rect 44086 2408 44142 2417
rect 44086 2343 44142 2352
rect 44100 2310 44128 2343
rect 44088 2304 44140 2310
rect 44088 2246 44140 2252
rect -10 0 102 800
rect 1278 0 1390 800
rect 3210 0 3322 800
rect 4498 0 4610 800
rect 6430 0 6542 800
rect 7718 0 7830 800
rect 9650 0 9762 800
rect 10938 0 11050 800
rect 12870 0 12982 800
rect 14158 0 14270 800
rect 16090 0 16202 800
rect 17378 0 17490 800
rect 19310 0 19422 800
rect 20598 0 20710 800
rect 22530 0 22642 800
rect 23818 0 23930 800
rect 25750 0 25862 800
rect 27038 0 27150 800
rect 28970 0 29082 800
rect 30258 0 30370 800
rect 32190 0 32302 800
rect 33478 0 33590 800
rect 35410 0 35522 800
rect 36698 0 36810 800
rect 38630 0 38742 800
rect 39918 0 40030 800
rect 41850 0 41962 800
rect 43782 0 43894 800
rect 44192 785 44220 3470
rect 44742 3292 45050 3301
rect 44742 3290 44748 3292
rect 44804 3290 44828 3292
rect 44884 3290 44908 3292
rect 44964 3290 44988 3292
rect 45044 3290 45050 3292
rect 44804 3238 44806 3290
rect 44986 3238 44988 3290
rect 44742 3236 44748 3238
rect 44804 3236 44828 3238
rect 44884 3236 44908 3238
rect 44964 3236 44988 3238
rect 45044 3236 45050 3238
rect 44742 3227 45050 3236
rect 45100 2984 45152 2990
rect 45100 2926 45152 2932
rect 44742 2204 45050 2213
rect 44742 2202 44748 2204
rect 44804 2202 44828 2204
rect 44884 2202 44908 2204
rect 44964 2202 44988 2204
rect 45044 2202 45050 2204
rect 44804 2150 44806 2202
rect 44986 2150 44988 2202
rect 44742 2148 44748 2150
rect 44804 2148 44828 2150
rect 44884 2148 44908 2150
rect 44964 2148 44988 2150
rect 45044 2148 45050 2150
rect 44742 2139 45050 2148
rect 45112 800 45140 2926
rect 44178 776 44234 785
rect 44178 711 44234 720
rect 45070 0 45182 800
<< via2 >>
rect 3974 18400 4030 18456
rect 2226 17040 2282 17096
rect 1582 15000 1638 15056
rect 11904 17434 11960 17436
rect 11984 17434 12040 17436
rect 12064 17434 12120 17436
rect 12144 17434 12200 17436
rect 11904 17382 11950 17434
rect 11950 17382 11960 17434
rect 11984 17382 12014 17434
rect 12014 17382 12026 17434
rect 12026 17382 12040 17434
rect 12064 17382 12078 17434
rect 12078 17382 12090 17434
rect 12090 17382 12120 17434
rect 12144 17382 12154 17434
rect 12154 17382 12200 17434
rect 11904 17380 11960 17382
rect 11984 17380 12040 17382
rect 12064 17380 12120 17382
rect 12144 17380 12200 17382
rect 22852 17434 22908 17436
rect 22932 17434 22988 17436
rect 23012 17434 23068 17436
rect 23092 17434 23148 17436
rect 22852 17382 22898 17434
rect 22898 17382 22908 17434
rect 22932 17382 22962 17434
rect 22962 17382 22974 17434
rect 22974 17382 22988 17434
rect 23012 17382 23026 17434
rect 23026 17382 23038 17434
rect 23038 17382 23068 17434
rect 23092 17382 23102 17434
rect 23102 17382 23148 17434
rect 22852 17380 22908 17382
rect 22932 17380 22988 17382
rect 23012 17380 23068 17382
rect 23092 17380 23148 17382
rect 33800 17434 33856 17436
rect 33880 17434 33936 17436
rect 33960 17434 34016 17436
rect 34040 17434 34096 17436
rect 33800 17382 33846 17434
rect 33846 17382 33856 17434
rect 33880 17382 33910 17434
rect 33910 17382 33922 17434
rect 33922 17382 33936 17434
rect 33960 17382 33974 17434
rect 33974 17382 33986 17434
rect 33986 17382 34016 17434
rect 34040 17382 34050 17434
rect 34050 17382 34096 17434
rect 33800 17380 33856 17382
rect 33880 17380 33936 17382
rect 33960 17380 34016 17382
rect 34040 17380 34096 17382
rect 1582 13640 1638 13696
rect 1582 10240 1638 10296
rect 4066 11620 4122 11656
rect 4066 11600 4068 11620
rect 4068 11600 4120 11620
rect 4120 11600 4122 11620
rect 6430 16890 6486 16892
rect 6510 16890 6566 16892
rect 6590 16890 6646 16892
rect 6670 16890 6726 16892
rect 6430 16838 6476 16890
rect 6476 16838 6486 16890
rect 6510 16838 6540 16890
rect 6540 16838 6552 16890
rect 6552 16838 6566 16890
rect 6590 16838 6604 16890
rect 6604 16838 6616 16890
rect 6616 16838 6646 16890
rect 6670 16838 6680 16890
rect 6680 16838 6726 16890
rect 6430 16836 6486 16838
rect 6510 16836 6566 16838
rect 6590 16836 6646 16838
rect 6670 16836 6726 16838
rect 6430 15802 6486 15804
rect 6510 15802 6566 15804
rect 6590 15802 6646 15804
rect 6670 15802 6726 15804
rect 6430 15750 6476 15802
rect 6476 15750 6486 15802
rect 6510 15750 6540 15802
rect 6540 15750 6552 15802
rect 6552 15750 6566 15802
rect 6590 15750 6604 15802
rect 6604 15750 6616 15802
rect 6616 15750 6646 15802
rect 6670 15750 6680 15802
rect 6680 15750 6726 15802
rect 6430 15748 6486 15750
rect 6510 15748 6566 15750
rect 6590 15748 6646 15750
rect 6670 15748 6726 15750
rect 6430 14714 6486 14716
rect 6510 14714 6566 14716
rect 6590 14714 6646 14716
rect 6670 14714 6726 14716
rect 6430 14662 6476 14714
rect 6476 14662 6486 14714
rect 6510 14662 6540 14714
rect 6540 14662 6552 14714
rect 6552 14662 6566 14714
rect 6590 14662 6604 14714
rect 6604 14662 6616 14714
rect 6616 14662 6646 14714
rect 6670 14662 6680 14714
rect 6680 14662 6726 14714
rect 6430 14660 6486 14662
rect 6510 14660 6566 14662
rect 6590 14660 6646 14662
rect 6670 14660 6726 14662
rect 6430 13626 6486 13628
rect 6510 13626 6566 13628
rect 6590 13626 6646 13628
rect 6670 13626 6726 13628
rect 6430 13574 6476 13626
rect 6476 13574 6486 13626
rect 6510 13574 6540 13626
rect 6540 13574 6552 13626
rect 6552 13574 6566 13626
rect 6590 13574 6604 13626
rect 6604 13574 6616 13626
rect 6616 13574 6646 13626
rect 6670 13574 6680 13626
rect 6680 13574 6726 13626
rect 6430 13572 6486 13574
rect 6510 13572 6566 13574
rect 6590 13572 6646 13574
rect 6670 13572 6726 13574
rect 1582 8200 1638 8256
rect 1582 6840 1638 6896
rect 6430 12538 6486 12540
rect 6510 12538 6566 12540
rect 6590 12538 6646 12540
rect 6670 12538 6726 12540
rect 6430 12486 6476 12538
rect 6476 12486 6486 12538
rect 6510 12486 6540 12538
rect 6540 12486 6552 12538
rect 6552 12486 6566 12538
rect 6590 12486 6604 12538
rect 6604 12486 6616 12538
rect 6616 12486 6646 12538
rect 6670 12486 6680 12538
rect 6680 12486 6726 12538
rect 6430 12484 6486 12486
rect 6510 12484 6566 12486
rect 6590 12484 6646 12486
rect 6670 12484 6726 12486
rect 6430 11450 6486 11452
rect 6510 11450 6566 11452
rect 6590 11450 6646 11452
rect 6670 11450 6726 11452
rect 6430 11398 6476 11450
rect 6476 11398 6486 11450
rect 6510 11398 6540 11450
rect 6540 11398 6552 11450
rect 6552 11398 6566 11450
rect 6590 11398 6604 11450
rect 6604 11398 6616 11450
rect 6616 11398 6646 11450
rect 6670 11398 6680 11450
rect 6680 11398 6726 11450
rect 6430 11396 6486 11398
rect 6510 11396 6566 11398
rect 6590 11396 6646 11398
rect 6670 11396 6726 11398
rect 6430 10362 6486 10364
rect 6510 10362 6566 10364
rect 6590 10362 6646 10364
rect 6670 10362 6726 10364
rect 6430 10310 6476 10362
rect 6476 10310 6486 10362
rect 6510 10310 6540 10362
rect 6540 10310 6552 10362
rect 6552 10310 6566 10362
rect 6590 10310 6604 10362
rect 6604 10310 6616 10362
rect 6616 10310 6646 10362
rect 6670 10310 6680 10362
rect 6680 10310 6726 10362
rect 6430 10308 6486 10310
rect 6510 10308 6566 10310
rect 6590 10308 6646 10310
rect 6670 10308 6726 10310
rect 6430 9274 6486 9276
rect 6510 9274 6566 9276
rect 6590 9274 6646 9276
rect 6670 9274 6726 9276
rect 6430 9222 6476 9274
rect 6476 9222 6486 9274
rect 6510 9222 6540 9274
rect 6540 9222 6552 9274
rect 6552 9222 6566 9274
rect 6590 9222 6604 9274
rect 6604 9222 6616 9274
rect 6616 9222 6646 9274
rect 6670 9222 6680 9274
rect 6680 9222 6726 9274
rect 6430 9220 6486 9222
rect 6510 9220 6566 9222
rect 6590 9220 6646 9222
rect 6670 9220 6726 9222
rect 6430 8186 6486 8188
rect 6510 8186 6566 8188
rect 6590 8186 6646 8188
rect 6670 8186 6726 8188
rect 6430 8134 6476 8186
rect 6476 8134 6486 8186
rect 6510 8134 6540 8186
rect 6540 8134 6552 8186
rect 6552 8134 6566 8186
rect 6590 8134 6604 8186
rect 6604 8134 6616 8186
rect 6616 8134 6646 8186
rect 6670 8134 6680 8186
rect 6680 8134 6726 8186
rect 6430 8132 6486 8134
rect 6510 8132 6566 8134
rect 6590 8132 6646 8134
rect 6670 8132 6726 8134
rect 6430 7098 6486 7100
rect 6510 7098 6566 7100
rect 6590 7098 6646 7100
rect 6670 7098 6726 7100
rect 6430 7046 6476 7098
rect 6476 7046 6486 7098
rect 6510 7046 6540 7098
rect 6540 7046 6552 7098
rect 6552 7046 6566 7098
rect 6590 7046 6604 7098
rect 6604 7046 6616 7098
rect 6616 7046 6646 7098
rect 6670 7046 6680 7098
rect 6680 7046 6726 7098
rect 6430 7044 6486 7046
rect 6510 7044 6566 7046
rect 6590 7044 6646 7046
rect 6670 7044 6726 7046
rect 6430 6010 6486 6012
rect 6510 6010 6566 6012
rect 6590 6010 6646 6012
rect 6670 6010 6726 6012
rect 6430 5958 6476 6010
rect 6476 5958 6486 6010
rect 6510 5958 6540 6010
rect 6540 5958 6552 6010
rect 6552 5958 6566 6010
rect 6590 5958 6604 6010
rect 6604 5958 6616 6010
rect 6616 5958 6646 6010
rect 6670 5958 6680 6010
rect 6680 5958 6726 6010
rect 6430 5956 6486 5958
rect 6510 5956 6566 5958
rect 6590 5956 6646 5958
rect 6670 5956 6726 5958
rect 1398 4800 1454 4856
rect 6430 4922 6486 4924
rect 6510 4922 6566 4924
rect 6590 4922 6646 4924
rect 6670 4922 6726 4924
rect 6430 4870 6476 4922
rect 6476 4870 6486 4922
rect 6510 4870 6540 4922
rect 6540 4870 6552 4922
rect 6552 4870 6566 4922
rect 6590 4870 6604 4922
rect 6604 4870 6616 4922
rect 6616 4870 6646 4922
rect 6670 4870 6680 4922
rect 6680 4870 6726 4922
rect 6430 4868 6486 4870
rect 6510 4868 6566 4870
rect 6590 4868 6646 4870
rect 6670 4868 6726 4870
rect 6430 3834 6486 3836
rect 6510 3834 6566 3836
rect 6590 3834 6646 3836
rect 6670 3834 6726 3836
rect 6430 3782 6476 3834
rect 6476 3782 6486 3834
rect 6510 3782 6540 3834
rect 6540 3782 6552 3834
rect 6552 3782 6566 3834
rect 6590 3782 6604 3834
rect 6604 3782 6616 3834
rect 6616 3782 6646 3834
rect 6670 3782 6680 3834
rect 6680 3782 6726 3834
rect 6430 3780 6486 3782
rect 6510 3780 6566 3782
rect 6590 3780 6646 3782
rect 6670 3780 6726 3782
rect 1582 3476 1584 3496
rect 1584 3476 1636 3496
rect 1636 3476 1638 3496
rect 1582 3440 1638 3476
rect 11904 16346 11960 16348
rect 11984 16346 12040 16348
rect 12064 16346 12120 16348
rect 12144 16346 12200 16348
rect 11904 16294 11950 16346
rect 11950 16294 11960 16346
rect 11984 16294 12014 16346
rect 12014 16294 12026 16346
rect 12026 16294 12040 16346
rect 12064 16294 12078 16346
rect 12078 16294 12090 16346
rect 12090 16294 12120 16346
rect 12144 16294 12154 16346
rect 12154 16294 12200 16346
rect 11904 16292 11960 16294
rect 11984 16292 12040 16294
rect 12064 16292 12120 16294
rect 12144 16292 12200 16294
rect 11904 15258 11960 15260
rect 11984 15258 12040 15260
rect 12064 15258 12120 15260
rect 12144 15258 12200 15260
rect 11904 15206 11950 15258
rect 11950 15206 11960 15258
rect 11984 15206 12014 15258
rect 12014 15206 12026 15258
rect 12026 15206 12040 15258
rect 12064 15206 12078 15258
rect 12078 15206 12090 15258
rect 12090 15206 12120 15258
rect 12144 15206 12154 15258
rect 12154 15206 12200 15258
rect 11904 15204 11960 15206
rect 11984 15204 12040 15206
rect 12064 15204 12120 15206
rect 12144 15204 12200 15206
rect 11904 14170 11960 14172
rect 11984 14170 12040 14172
rect 12064 14170 12120 14172
rect 12144 14170 12200 14172
rect 11904 14118 11950 14170
rect 11950 14118 11960 14170
rect 11984 14118 12014 14170
rect 12014 14118 12026 14170
rect 12026 14118 12040 14170
rect 12064 14118 12078 14170
rect 12078 14118 12090 14170
rect 12090 14118 12120 14170
rect 12144 14118 12154 14170
rect 12154 14118 12200 14170
rect 11904 14116 11960 14118
rect 11984 14116 12040 14118
rect 12064 14116 12120 14118
rect 12144 14116 12200 14118
rect 11904 13082 11960 13084
rect 11984 13082 12040 13084
rect 12064 13082 12120 13084
rect 12144 13082 12200 13084
rect 11904 13030 11950 13082
rect 11950 13030 11960 13082
rect 11984 13030 12014 13082
rect 12014 13030 12026 13082
rect 12026 13030 12040 13082
rect 12064 13030 12078 13082
rect 12078 13030 12090 13082
rect 12090 13030 12120 13082
rect 12144 13030 12154 13082
rect 12154 13030 12200 13082
rect 11904 13028 11960 13030
rect 11984 13028 12040 13030
rect 12064 13028 12120 13030
rect 12144 13028 12200 13030
rect 12070 12144 12126 12200
rect 11904 11994 11960 11996
rect 11984 11994 12040 11996
rect 12064 11994 12120 11996
rect 12144 11994 12200 11996
rect 11904 11942 11950 11994
rect 11950 11942 11960 11994
rect 11984 11942 12014 11994
rect 12014 11942 12026 11994
rect 12026 11942 12040 11994
rect 12064 11942 12078 11994
rect 12078 11942 12090 11994
rect 12090 11942 12120 11994
rect 12144 11942 12154 11994
rect 12154 11942 12200 11994
rect 11904 11940 11960 11942
rect 11984 11940 12040 11942
rect 12064 11940 12120 11942
rect 12144 11940 12200 11942
rect 8206 5636 8262 5672
rect 8206 5616 8208 5636
rect 8208 5616 8260 5636
rect 8260 5616 8262 5636
rect 6430 2746 6486 2748
rect 6510 2746 6566 2748
rect 6590 2746 6646 2748
rect 6670 2746 6726 2748
rect 6430 2694 6476 2746
rect 6476 2694 6486 2746
rect 6510 2694 6540 2746
rect 6540 2694 6552 2746
rect 6552 2694 6566 2746
rect 6590 2694 6604 2746
rect 6604 2694 6616 2746
rect 6616 2694 6646 2746
rect 6670 2694 6680 2746
rect 6680 2694 6726 2746
rect 6430 2692 6486 2694
rect 6510 2692 6566 2694
rect 6590 2692 6646 2694
rect 6670 2692 6726 2694
rect 11904 10906 11960 10908
rect 11984 10906 12040 10908
rect 12064 10906 12120 10908
rect 12144 10906 12200 10908
rect 11904 10854 11950 10906
rect 11950 10854 11960 10906
rect 11984 10854 12014 10906
rect 12014 10854 12026 10906
rect 12026 10854 12040 10906
rect 12064 10854 12078 10906
rect 12078 10854 12090 10906
rect 12090 10854 12120 10906
rect 12144 10854 12154 10906
rect 12154 10854 12200 10906
rect 11904 10852 11960 10854
rect 11984 10852 12040 10854
rect 12064 10852 12120 10854
rect 12144 10852 12200 10854
rect 11904 9818 11960 9820
rect 11984 9818 12040 9820
rect 12064 9818 12120 9820
rect 12144 9818 12200 9820
rect 11904 9766 11950 9818
rect 11950 9766 11960 9818
rect 11984 9766 12014 9818
rect 12014 9766 12026 9818
rect 12026 9766 12040 9818
rect 12064 9766 12078 9818
rect 12078 9766 12090 9818
rect 12090 9766 12120 9818
rect 12144 9766 12154 9818
rect 12154 9766 12200 9818
rect 11904 9764 11960 9766
rect 11984 9764 12040 9766
rect 12064 9764 12120 9766
rect 12144 9764 12200 9766
rect 11904 8730 11960 8732
rect 11984 8730 12040 8732
rect 12064 8730 12120 8732
rect 12144 8730 12200 8732
rect 11904 8678 11950 8730
rect 11950 8678 11960 8730
rect 11984 8678 12014 8730
rect 12014 8678 12026 8730
rect 12026 8678 12040 8730
rect 12064 8678 12078 8730
rect 12078 8678 12090 8730
rect 12090 8678 12120 8730
rect 12144 8678 12154 8730
rect 12154 8678 12200 8730
rect 11904 8676 11960 8678
rect 11984 8676 12040 8678
rect 12064 8676 12120 8678
rect 12144 8676 12200 8678
rect 11904 7642 11960 7644
rect 11984 7642 12040 7644
rect 12064 7642 12120 7644
rect 12144 7642 12200 7644
rect 11904 7590 11950 7642
rect 11950 7590 11960 7642
rect 11984 7590 12014 7642
rect 12014 7590 12026 7642
rect 12026 7590 12040 7642
rect 12064 7590 12078 7642
rect 12078 7590 12090 7642
rect 12090 7590 12120 7642
rect 12144 7590 12154 7642
rect 12154 7590 12200 7642
rect 11904 7588 11960 7590
rect 11984 7588 12040 7590
rect 12064 7588 12120 7590
rect 12144 7588 12200 7590
rect 11904 6554 11960 6556
rect 11984 6554 12040 6556
rect 12064 6554 12120 6556
rect 12144 6554 12200 6556
rect 11904 6502 11950 6554
rect 11950 6502 11960 6554
rect 11984 6502 12014 6554
rect 12014 6502 12026 6554
rect 12026 6502 12040 6554
rect 12064 6502 12078 6554
rect 12078 6502 12090 6554
rect 12090 6502 12120 6554
rect 12144 6502 12154 6554
rect 12154 6502 12200 6554
rect 11904 6500 11960 6502
rect 11984 6500 12040 6502
rect 12064 6500 12120 6502
rect 12144 6500 12200 6502
rect 11904 5466 11960 5468
rect 11984 5466 12040 5468
rect 12064 5466 12120 5468
rect 12144 5466 12200 5468
rect 11904 5414 11950 5466
rect 11950 5414 11960 5466
rect 11984 5414 12014 5466
rect 12014 5414 12026 5466
rect 12026 5414 12040 5466
rect 12064 5414 12078 5466
rect 12078 5414 12090 5466
rect 12090 5414 12120 5466
rect 12144 5414 12154 5466
rect 12154 5414 12200 5466
rect 11904 5412 11960 5414
rect 11984 5412 12040 5414
rect 12064 5412 12120 5414
rect 12144 5412 12200 5414
rect 11904 4378 11960 4380
rect 11984 4378 12040 4380
rect 12064 4378 12120 4380
rect 12144 4378 12200 4380
rect 11904 4326 11950 4378
rect 11950 4326 11960 4378
rect 11984 4326 12014 4378
rect 12014 4326 12026 4378
rect 12026 4326 12040 4378
rect 12064 4326 12078 4378
rect 12078 4326 12090 4378
rect 12090 4326 12120 4378
rect 12144 4326 12154 4378
rect 12154 4326 12200 4378
rect 11904 4324 11960 4326
rect 11984 4324 12040 4326
rect 12064 4324 12120 4326
rect 12144 4324 12200 4326
rect 13450 11736 13506 11792
rect 15474 11736 15530 11792
rect 14278 10004 14280 10024
rect 14280 10004 14332 10024
rect 14332 10004 14334 10024
rect 14278 9968 14334 10004
rect 12714 5616 12770 5672
rect 17378 16890 17434 16892
rect 17458 16890 17514 16892
rect 17538 16890 17594 16892
rect 17618 16890 17674 16892
rect 17378 16838 17424 16890
rect 17424 16838 17434 16890
rect 17458 16838 17488 16890
rect 17488 16838 17500 16890
rect 17500 16838 17514 16890
rect 17538 16838 17552 16890
rect 17552 16838 17564 16890
rect 17564 16838 17594 16890
rect 17618 16838 17628 16890
rect 17628 16838 17674 16890
rect 17378 16836 17434 16838
rect 17458 16836 17514 16838
rect 17538 16836 17594 16838
rect 17618 16836 17674 16838
rect 22852 16346 22908 16348
rect 22932 16346 22988 16348
rect 23012 16346 23068 16348
rect 23092 16346 23148 16348
rect 22852 16294 22898 16346
rect 22898 16294 22908 16346
rect 22932 16294 22962 16346
rect 22962 16294 22974 16346
rect 22974 16294 22988 16346
rect 23012 16294 23026 16346
rect 23026 16294 23038 16346
rect 23038 16294 23068 16346
rect 23092 16294 23102 16346
rect 23102 16294 23148 16346
rect 22852 16292 22908 16294
rect 22932 16292 22988 16294
rect 23012 16292 23068 16294
rect 23092 16292 23148 16294
rect 17378 15802 17434 15804
rect 17458 15802 17514 15804
rect 17538 15802 17594 15804
rect 17618 15802 17674 15804
rect 17378 15750 17424 15802
rect 17424 15750 17434 15802
rect 17458 15750 17488 15802
rect 17488 15750 17500 15802
rect 17500 15750 17514 15802
rect 17538 15750 17552 15802
rect 17552 15750 17564 15802
rect 17564 15750 17594 15802
rect 17618 15750 17628 15802
rect 17628 15750 17674 15802
rect 17378 15748 17434 15750
rect 17458 15748 17514 15750
rect 17538 15748 17594 15750
rect 17618 15748 17674 15750
rect 17378 14714 17434 14716
rect 17458 14714 17514 14716
rect 17538 14714 17594 14716
rect 17618 14714 17674 14716
rect 17378 14662 17424 14714
rect 17424 14662 17434 14714
rect 17458 14662 17488 14714
rect 17488 14662 17500 14714
rect 17500 14662 17514 14714
rect 17538 14662 17552 14714
rect 17552 14662 17564 14714
rect 17564 14662 17594 14714
rect 17618 14662 17628 14714
rect 17628 14662 17674 14714
rect 17378 14660 17434 14662
rect 17458 14660 17514 14662
rect 17538 14660 17594 14662
rect 17618 14660 17674 14662
rect 17378 13626 17434 13628
rect 17458 13626 17514 13628
rect 17538 13626 17594 13628
rect 17618 13626 17674 13628
rect 17378 13574 17424 13626
rect 17424 13574 17434 13626
rect 17458 13574 17488 13626
rect 17488 13574 17500 13626
rect 17500 13574 17514 13626
rect 17538 13574 17552 13626
rect 17552 13574 17564 13626
rect 17564 13574 17594 13626
rect 17618 13574 17628 13626
rect 17628 13574 17674 13626
rect 17378 13572 17434 13574
rect 17458 13572 17514 13574
rect 17538 13572 17594 13574
rect 17618 13572 17674 13574
rect 22852 15258 22908 15260
rect 22932 15258 22988 15260
rect 23012 15258 23068 15260
rect 23092 15258 23148 15260
rect 22852 15206 22898 15258
rect 22898 15206 22908 15258
rect 22932 15206 22962 15258
rect 22962 15206 22974 15258
rect 22974 15206 22988 15258
rect 23012 15206 23026 15258
rect 23026 15206 23038 15258
rect 23038 15206 23068 15258
rect 23092 15206 23102 15258
rect 23102 15206 23148 15258
rect 22852 15204 22908 15206
rect 22932 15204 22988 15206
rect 23012 15204 23068 15206
rect 23092 15204 23148 15206
rect 22852 14170 22908 14172
rect 22932 14170 22988 14172
rect 23012 14170 23068 14172
rect 23092 14170 23148 14172
rect 22852 14118 22898 14170
rect 22898 14118 22908 14170
rect 22932 14118 22962 14170
rect 22962 14118 22974 14170
rect 22974 14118 22988 14170
rect 23012 14118 23026 14170
rect 23026 14118 23038 14170
rect 23038 14118 23068 14170
rect 23092 14118 23102 14170
rect 23102 14118 23148 14170
rect 22852 14116 22908 14118
rect 22932 14116 22988 14118
rect 23012 14116 23068 14118
rect 23092 14116 23148 14118
rect 17378 12538 17434 12540
rect 17458 12538 17514 12540
rect 17538 12538 17594 12540
rect 17618 12538 17674 12540
rect 17378 12486 17424 12538
rect 17424 12486 17434 12538
rect 17458 12486 17488 12538
rect 17488 12486 17500 12538
rect 17500 12486 17514 12538
rect 17538 12486 17552 12538
rect 17552 12486 17564 12538
rect 17564 12486 17594 12538
rect 17618 12486 17628 12538
rect 17628 12486 17674 12538
rect 17378 12484 17434 12486
rect 17458 12484 17514 12486
rect 17538 12484 17594 12486
rect 17618 12484 17674 12486
rect 18326 12144 18382 12200
rect 17378 11450 17434 11452
rect 17458 11450 17514 11452
rect 17538 11450 17594 11452
rect 17618 11450 17674 11452
rect 17378 11398 17424 11450
rect 17424 11398 17434 11450
rect 17458 11398 17488 11450
rect 17488 11398 17500 11450
rect 17500 11398 17514 11450
rect 17538 11398 17552 11450
rect 17552 11398 17564 11450
rect 17564 11398 17594 11450
rect 17618 11398 17628 11450
rect 17628 11398 17674 11450
rect 17378 11396 17434 11398
rect 17458 11396 17514 11398
rect 17538 11396 17594 11398
rect 17618 11396 17674 11398
rect 17378 10362 17434 10364
rect 17458 10362 17514 10364
rect 17538 10362 17594 10364
rect 17618 10362 17674 10364
rect 17378 10310 17424 10362
rect 17424 10310 17434 10362
rect 17458 10310 17488 10362
rect 17488 10310 17500 10362
rect 17500 10310 17514 10362
rect 17538 10310 17552 10362
rect 17552 10310 17564 10362
rect 17564 10310 17594 10362
rect 17618 10310 17628 10362
rect 17628 10310 17674 10362
rect 17378 10308 17434 10310
rect 17458 10308 17514 10310
rect 17538 10308 17594 10310
rect 17618 10308 17674 10310
rect 17378 9274 17434 9276
rect 17458 9274 17514 9276
rect 17538 9274 17594 9276
rect 17618 9274 17674 9276
rect 17378 9222 17424 9274
rect 17424 9222 17434 9274
rect 17458 9222 17488 9274
rect 17488 9222 17500 9274
rect 17500 9222 17514 9274
rect 17538 9222 17552 9274
rect 17552 9222 17564 9274
rect 17564 9222 17594 9274
rect 17618 9222 17628 9274
rect 17628 9222 17674 9274
rect 17378 9220 17434 9222
rect 17458 9220 17514 9222
rect 17538 9220 17594 9222
rect 17618 9220 17674 9222
rect 19246 11736 19302 11792
rect 18694 9968 18750 10024
rect 17378 8186 17434 8188
rect 17458 8186 17514 8188
rect 17538 8186 17594 8188
rect 17618 8186 17674 8188
rect 17378 8134 17424 8186
rect 17424 8134 17434 8186
rect 17458 8134 17488 8186
rect 17488 8134 17500 8186
rect 17500 8134 17514 8186
rect 17538 8134 17552 8186
rect 17552 8134 17564 8186
rect 17564 8134 17594 8186
rect 17618 8134 17628 8186
rect 17628 8134 17674 8186
rect 17378 8132 17434 8134
rect 17458 8132 17514 8134
rect 17538 8132 17594 8134
rect 17618 8132 17674 8134
rect 17378 7098 17434 7100
rect 17458 7098 17514 7100
rect 17538 7098 17594 7100
rect 17618 7098 17674 7100
rect 17378 7046 17424 7098
rect 17424 7046 17434 7098
rect 17458 7046 17488 7098
rect 17488 7046 17500 7098
rect 17500 7046 17514 7098
rect 17538 7046 17552 7098
rect 17552 7046 17564 7098
rect 17564 7046 17594 7098
rect 17618 7046 17628 7098
rect 17628 7046 17674 7098
rect 17378 7044 17434 7046
rect 17458 7044 17514 7046
rect 17538 7044 17594 7046
rect 17618 7044 17674 7046
rect 17378 6010 17434 6012
rect 17458 6010 17514 6012
rect 17538 6010 17594 6012
rect 17618 6010 17674 6012
rect 17378 5958 17424 6010
rect 17424 5958 17434 6010
rect 17458 5958 17488 6010
rect 17488 5958 17500 6010
rect 17500 5958 17514 6010
rect 17538 5958 17552 6010
rect 17552 5958 17564 6010
rect 17564 5958 17594 6010
rect 17618 5958 17628 6010
rect 17628 5958 17674 6010
rect 17378 5956 17434 5958
rect 17458 5956 17514 5958
rect 17538 5956 17594 5958
rect 17618 5956 17674 5958
rect 22006 10648 22062 10704
rect 20442 7792 20498 7848
rect 11904 3290 11960 3292
rect 11984 3290 12040 3292
rect 12064 3290 12120 3292
rect 12144 3290 12200 3292
rect 11904 3238 11950 3290
rect 11950 3238 11960 3290
rect 11984 3238 12014 3290
rect 12014 3238 12026 3290
rect 12026 3238 12040 3290
rect 12064 3238 12078 3290
rect 12078 3238 12090 3290
rect 12090 3238 12120 3290
rect 12144 3238 12154 3290
rect 12154 3238 12200 3290
rect 11904 3236 11960 3238
rect 11984 3236 12040 3238
rect 12064 3236 12120 3238
rect 12144 3236 12200 3238
rect 17378 4922 17434 4924
rect 17458 4922 17514 4924
rect 17538 4922 17594 4924
rect 17618 4922 17674 4924
rect 17378 4870 17424 4922
rect 17424 4870 17434 4922
rect 17458 4870 17488 4922
rect 17488 4870 17500 4922
rect 17500 4870 17514 4922
rect 17538 4870 17552 4922
rect 17552 4870 17564 4922
rect 17564 4870 17594 4922
rect 17618 4870 17628 4922
rect 17628 4870 17674 4922
rect 17378 4868 17434 4870
rect 17458 4868 17514 4870
rect 17538 4868 17594 4870
rect 17618 4868 17674 4870
rect 17378 3834 17434 3836
rect 17458 3834 17514 3836
rect 17538 3834 17594 3836
rect 17618 3834 17674 3836
rect 17378 3782 17424 3834
rect 17424 3782 17434 3834
rect 17458 3782 17488 3834
rect 17488 3782 17500 3834
rect 17500 3782 17514 3834
rect 17538 3782 17552 3834
rect 17552 3782 17564 3834
rect 17564 3782 17594 3834
rect 17618 3782 17628 3834
rect 17628 3782 17674 3834
rect 17378 3780 17434 3782
rect 17458 3780 17514 3782
rect 17538 3780 17594 3782
rect 17618 3780 17674 3782
rect 17378 2746 17434 2748
rect 17458 2746 17514 2748
rect 17538 2746 17594 2748
rect 17618 2746 17674 2748
rect 17378 2694 17424 2746
rect 17424 2694 17434 2746
rect 17458 2694 17488 2746
rect 17488 2694 17500 2746
rect 17500 2694 17514 2746
rect 17538 2694 17552 2746
rect 17552 2694 17564 2746
rect 17564 2694 17594 2746
rect 17618 2694 17628 2746
rect 17628 2694 17674 2746
rect 17378 2692 17434 2694
rect 17458 2692 17514 2694
rect 17538 2692 17594 2694
rect 17618 2692 17674 2694
rect 20626 5616 20682 5672
rect 22374 7384 22430 7440
rect 22852 13082 22908 13084
rect 22932 13082 22988 13084
rect 23012 13082 23068 13084
rect 23092 13082 23148 13084
rect 22852 13030 22898 13082
rect 22898 13030 22908 13082
rect 22932 13030 22962 13082
rect 22962 13030 22974 13082
rect 22974 13030 22988 13082
rect 23012 13030 23026 13082
rect 23026 13030 23038 13082
rect 23038 13030 23068 13082
rect 23092 13030 23102 13082
rect 23102 13030 23148 13082
rect 22852 13028 22908 13030
rect 22932 13028 22988 13030
rect 23012 13028 23068 13030
rect 23092 13028 23148 13030
rect 22852 11994 22908 11996
rect 22932 11994 22988 11996
rect 23012 11994 23068 11996
rect 23092 11994 23148 11996
rect 22852 11942 22898 11994
rect 22898 11942 22908 11994
rect 22932 11942 22962 11994
rect 22962 11942 22974 11994
rect 22974 11942 22988 11994
rect 23012 11942 23026 11994
rect 23026 11942 23038 11994
rect 23038 11942 23068 11994
rect 23092 11942 23102 11994
rect 23102 11942 23148 11994
rect 22852 11940 22908 11942
rect 22932 11940 22988 11942
rect 23012 11940 23068 11942
rect 23092 11940 23148 11942
rect 28326 16890 28382 16892
rect 28406 16890 28462 16892
rect 28486 16890 28542 16892
rect 28566 16890 28622 16892
rect 28326 16838 28372 16890
rect 28372 16838 28382 16890
rect 28406 16838 28436 16890
rect 28436 16838 28448 16890
rect 28448 16838 28462 16890
rect 28486 16838 28500 16890
rect 28500 16838 28512 16890
rect 28512 16838 28542 16890
rect 28566 16838 28576 16890
rect 28576 16838 28622 16890
rect 28326 16836 28382 16838
rect 28406 16836 28462 16838
rect 28486 16836 28542 16838
rect 28566 16836 28622 16838
rect 28326 15802 28382 15804
rect 28406 15802 28462 15804
rect 28486 15802 28542 15804
rect 28566 15802 28622 15804
rect 28326 15750 28372 15802
rect 28372 15750 28382 15802
rect 28406 15750 28436 15802
rect 28436 15750 28448 15802
rect 28448 15750 28462 15802
rect 28486 15750 28500 15802
rect 28500 15750 28512 15802
rect 28512 15750 28542 15802
rect 28566 15750 28576 15802
rect 28576 15750 28622 15802
rect 28326 15748 28382 15750
rect 28406 15748 28462 15750
rect 28486 15748 28542 15750
rect 28566 15748 28622 15750
rect 28326 14714 28382 14716
rect 28406 14714 28462 14716
rect 28486 14714 28542 14716
rect 28566 14714 28622 14716
rect 28326 14662 28372 14714
rect 28372 14662 28382 14714
rect 28406 14662 28436 14714
rect 28436 14662 28448 14714
rect 28448 14662 28462 14714
rect 28486 14662 28500 14714
rect 28500 14662 28512 14714
rect 28512 14662 28542 14714
rect 28566 14662 28576 14714
rect 28576 14662 28622 14714
rect 28326 14660 28382 14662
rect 28406 14660 28462 14662
rect 28486 14660 28542 14662
rect 28566 14660 28622 14662
rect 28326 13626 28382 13628
rect 28406 13626 28462 13628
rect 28486 13626 28542 13628
rect 28566 13626 28622 13628
rect 28326 13574 28372 13626
rect 28372 13574 28382 13626
rect 28406 13574 28436 13626
rect 28436 13574 28448 13626
rect 28448 13574 28462 13626
rect 28486 13574 28500 13626
rect 28500 13574 28512 13626
rect 28512 13574 28542 13626
rect 28566 13574 28576 13626
rect 28576 13574 28622 13626
rect 28326 13572 28382 13574
rect 28406 13572 28462 13574
rect 28486 13572 28542 13574
rect 28566 13572 28622 13574
rect 33800 16346 33856 16348
rect 33880 16346 33936 16348
rect 33960 16346 34016 16348
rect 34040 16346 34096 16348
rect 33800 16294 33846 16346
rect 33846 16294 33856 16346
rect 33880 16294 33910 16346
rect 33910 16294 33922 16346
rect 33922 16294 33936 16346
rect 33960 16294 33974 16346
rect 33974 16294 33986 16346
rect 33986 16294 34016 16346
rect 34040 16294 34050 16346
rect 34050 16294 34096 16346
rect 33800 16292 33856 16294
rect 33880 16292 33936 16294
rect 33960 16292 34016 16294
rect 34040 16292 34096 16294
rect 33800 15258 33856 15260
rect 33880 15258 33936 15260
rect 33960 15258 34016 15260
rect 34040 15258 34096 15260
rect 33800 15206 33846 15258
rect 33846 15206 33856 15258
rect 33880 15206 33910 15258
rect 33910 15206 33922 15258
rect 33922 15206 33936 15258
rect 33960 15206 33974 15258
rect 33974 15206 33986 15258
rect 33986 15206 34016 15258
rect 34040 15206 34050 15258
rect 34050 15206 34096 15258
rect 33800 15204 33856 15206
rect 33880 15204 33936 15206
rect 33960 15204 34016 15206
rect 34040 15204 34096 15206
rect 33800 14170 33856 14172
rect 33880 14170 33936 14172
rect 33960 14170 34016 14172
rect 34040 14170 34096 14172
rect 33800 14118 33846 14170
rect 33846 14118 33856 14170
rect 33880 14118 33910 14170
rect 33910 14118 33922 14170
rect 33922 14118 33936 14170
rect 33960 14118 33974 14170
rect 33974 14118 33986 14170
rect 33986 14118 34016 14170
rect 34040 14118 34050 14170
rect 34050 14118 34096 14170
rect 33800 14116 33856 14118
rect 33880 14116 33936 14118
rect 33960 14116 34016 14118
rect 34040 14116 34096 14118
rect 22852 10906 22908 10908
rect 22932 10906 22988 10908
rect 23012 10906 23068 10908
rect 23092 10906 23148 10908
rect 22852 10854 22898 10906
rect 22898 10854 22908 10906
rect 22932 10854 22962 10906
rect 22962 10854 22974 10906
rect 22974 10854 22988 10906
rect 23012 10854 23026 10906
rect 23026 10854 23038 10906
rect 23038 10854 23068 10906
rect 23092 10854 23102 10906
rect 23102 10854 23148 10906
rect 22852 10852 22908 10854
rect 22932 10852 22988 10854
rect 23012 10852 23068 10854
rect 23092 10852 23148 10854
rect 22852 9818 22908 9820
rect 22932 9818 22988 9820
rect 23012 9818 23068 9820
rect 23092 9818 23148 9820
rect 22852 9766 22898 9818
rect 22898 9766 22908 9818
rect 22932 9766 22962 9818
rect 22962 9766 22974 9818
rect 22974 9766 22988 9818
rect 23012 9766 23026 9818
rect 23026 9766 23038 9818
rect 23038 9766 23068 9818
rect 23092 9766 23102 9818
rect 23102 9766 23148 9818
rect 22852 9764 22908 9766
rect 22932 9764 22988 9766
rect 23012 9764 23068 9766
rect 23092 9764 23148 9766
rect 22852 8730 22908 8732
rect 22932 8730 22988 8732
rect 23012 8730 23068 8732
rect 23092 8730 23148 8732
rect 22852 8678 22898 8730
rect 22898 8678 22908 8730
rect 22932 8678 22962 8730
rect 22962 8678 22974 8730
rect 22974 8678 22988 8730
rect 23012 8678 23026 8730
rect 23026 8678 23038 8730
rect 23038 8678 23068 8730
rect 23092 8678 23102 8730
rect 23102 8678 23148 8730
rect 22852 8676 22908 8678
rect 22932 8676 22988 8678
rect 23012 8676 23068 8678
rect 23092 8676 23148 8678
rect 25778 10648 25834 10704
rect 28326 12538 28382 12540
rect 28406 12538 28462 12540
rect 28486 12538 28542 12540
rect 28566 12538 28622 12540
rect 28326 12486 28372 12538
rect 28372 12486 28382 12538
rect 28406 12486 28436 12538
rect 28436 12486 28448 12538
rect 28448 12486 28462 12538
rect 28486 12486 28500 12538
rect 28500 12486 28512 12538
rect 28512 12486 28542 12538
rect 28566 12486 28576 12538
rect 28576 12486 28622 12538
rect 28326 12484 28382 12486
rect 28406 12484 28462 12486
rect 28486 12484 28542 12486
rect 28566 12484 28622 12486
rect 29458 11772 29460 11792
rect 29460 11772 29512 11792
rect 29512 11772 29514 11792
rect 29458 11736 29514 11772
rect 28326 11450 28382 11452
rect 28406 11450 28462 11452
rect 28486 11450 28542 11452
rect 28566 11450 28622 11452
rect 28326 11398 28372 11450
rect 28372 11398 28382 11450
rect 28406 11398 28436 11450
rect 28436 11398 28448 11450
rect 28448 11398 28462 11450
rect 28486 11398 28500 11450
rect 28500 11398 28512 11450
rect 28512 11398 28542 11450
rect 28566 11398 28576 11450
rect 28576 11398 28622 11450
rect 28326 11396 28382 11398
rect 28406 11396 28462 11398
rect 28486 11396 28542 11398
rect 28566 11396 28622 11398
rect 28326 10362 28382 10364
rect 28406 10362 28462 10364
rect 28486 10362 28542 10364
rect 28566 10362 28622 10364
rect 28326 10310 28372 10362
rect 28372 10310 28382 10362
rect 28406 10310 28436 10362
rect 28436 10310 28448 10362
rect 28448 10310 28462 10362
rect 28486 10310 28500 10362
rect 28500 10310 28512 10362
rect 28512 10310 28542 10362
rect 28566 10310 28576 10362
rect 28576 10310 28622 10362
rect 28326 10308 28382 10310
rect 28406 10308 28462 10310
rect 28486 10308 28542 10310
rect 28566 10308 28622 10310
rect 28326 9274 28382 9276
rect 28406 9274 28462 9276
rect 28486 9274 28542 9276
rect 28566 9274 28622 9276
rect 28326 9222 28372 9274
rect 28372 9222 28382 9274
rect 28406 9222 28436 9274
rect 28436 9222 28448 9274
rect 28448 9222 28462 9274
rect 28486 9222 28500 9274
rect 28500 9222 28512 9274
rect 28512 9222 28542 9274
rect 28566 9222 28576 9274
rect 28576 9222 28622 9274
rect 28326 9220 28382 9222
rect 28406 9220 28462 9222
rect 28486 9220 28542 9222
rect 28566 9220 28622 9222
rect 26054 7792 26110 7848
rect 22852 7642 22908 7644
rect 22932 7642 22988 7644
rect 23012 7642 23068 7644
rect 23092 7642 23148 7644
rect 22852 7590 22898 7642
rect 22898 7590 22908 7642
rect 22932 7590 22962 7642
rect 22962 7590 22974 7642
rect 22974 7590 22988 7642
rect 23012 7590 23026 7642
rect 23026 7590 23038 7642
rect 23038 7590 23068 7642
rect 23092 7590 23102 7642
rect 23102 7590 23148 7642
rect 22852 7588 22908 7590
rect 22932 7588 22988 7590
rect 23012 7588 23068 7590
rect 23092 7588 23148 7590
rect 22852 6554 22908 6556
rect 22932 6554 22988 6556
rect 23012 6554 23068 6556
rect 23092 6554 23148 6556
rect 22852 6502 22898 6554
rect 22898 6502 22908 6554
rect 22932 6502 22962 6554
rect 22962 6502 22974 6554
rect 22974 6502 22988 6554
rect 23012 6502 23026 6554
rect 23026 6502 23038 6554
rect 23038 6502 23068 6554
rect 23092 6502 23102 6554
rect 23102 6502 23148 6554
rect 22852 6500 22908 6502
rect 22932 6500 22988 6502
rect 23012 6500 23068 6502
rect 23092 6500 23148 6502
rect 27434 6840 27490 6896
rect 22852 5466 22908 5468
rect 22932 5466 22988 5468
rect 23012 5466 23068 5468
rect 23092 5466 23148 5468
rect 22852 5414 22898 5466
rect 22898 5414 22908 5466
rect 22932 5414 22962 5466
rect 22962 5414 22974 5466
rect 22974 5414 22988 5466
rect 23012 5414 23026 5466
rect 23026 5414 23038 5466
rect 23038 5414 23068 5466
rect 23092 5414 23102 5466
rect 23102 5414 23148 5466
rect 22852 5412 22908 5414
rect 22932 5412 22988 5414
rect 23012 5412 23068 5414
rect 23092 5412 23148 5414
rect 26422 5652 26424 5672
rect 26424 5652 26476 5672
rect 26476 5652 26478 5672
rect 22852 4378 22908 4380
rect 22932 4378 22988 4380
rect 23012 4378 23068 4380
rect 23092 4378 23148 4380
rect 22852 4326 22898 4378
rect 22898 4326 22908 4378
rect 22932 4326 22962 4378
rect 22962 4326 22974 4378
rect 22974 4326 22988 4378
rect 23012 4326 23026 4378
rect 23026 4326 23038 4378
rect 23038 4326 23068 4378
rect 23092 4326 23102 4378
rect 23102 4326 23148 4378
rect 22852 4324 22908 4326
rect 22932 4324 22988 4326
rect 23012 4324 23068 4326
rect 23092 4324 23148 4326
rect 22852 3290 22908 3292
rect 22932 3290 22988 3292
rect 23012 3290 23068 3292
rect 23092 3290 23148 3292
rect 22852 3238 22898 3290
rect 22898 3238 22908 3290
rect 22932 3238 22962 3290
rect 22962 3238 22974 3290
rect 22974 3238 22988 3290
rect 23012 3238 23026 3290
rect 23026 3238 23038 3290
rect 23038 3238 23068 3290
rect 23092 3238 23102 3290
rect 23102 3238 23148 3290
rect 22852 3236 22908 3238
rect 22932 3236 22988 3238
rect 23012 3236 23068 3238
rect 23092 3236 23148 3238
rect 26422 5616 26478 5652
rect 1582 1400 1638 1456
rect 11904 2202 11960 2204
rect 11984 2202 12040 2204
rect 12064 2202 12120 2204
rect 12144 2202 12200 2204
rect 11904 2150 11950 2202
rect 11950 2150 11960 2202
rect 11984 2150 12014 2202
rect 12014 2150 12026 2202
rect 12026 2150 12040 2202
rect 12064 2150 12078 2202
rect 12078 2150 12090 2202
rect 12090 2150 12120 2202
rect 12144 2150 12154 2202
rect 12154 2150 12200 2202
rect 11904 2148 11960 2150
rect 11984 2148 12040 2150
rect 12064 2148 12120 2150
rect 12144 2148 12200 2150
rect 22852 2202 22908 2204
rect 22932 2202 22988 2204
rect 23012 2202 23068 2204
rect 23092 2202 23148 2204
rect 22852 2150 22898 2202
rect 22898 2150 22908 2202
rect 22932 2150 22962 2202
rect 22962 2150 22974 2202
rect 22974 2150 22988 2202
rect 23012 2150 23026 2202
rect 23026 2150 23038 2202
rect 23038 2150 23068 2202
rect 23092 2150 23102 2202
rect 23102 2150 23148 2202
rect 22852 2148 22908 2150
rect 22932 2148 22988 2150
rect 23012 2148 23068 2150
rect 23092 2148 23148 2150
rect 28326 8186 28382 8188
rect 28406 8186 28462 8188
rect 28486 8186 28542 8188
rect 28566 8186 28622 8188
rect 28326 8134 28372 8186
rect 28372 8134 28382 8186
rect 28406 8134 28436 8186
rect 28436 8134 28448 8186
rect 28448 8134 28462 8186
rect 28486 8134 28500 8186
rect 28500 8134 28512 8186
rect 28512 8134 28542 8186
rect 28566 8134 28576 8186
rect 28576 8134 28622 8186
rect 28326 8132 28382 8134
rect 28406 8132 28462 8134
rect 28486 8132 28542 8134
rect 28566 8132 28622 8134
rect 27710 7384 27766 7440
rect 28326 7098 28382 7100
rect 28406 7098 28462 7100
rect 28486 7098 28542 7100
rect 28566 7098 28622 7100
rect 28326 7046 28372 7098
rect 28372 7046 28382 7098
rect 28406 7046 28436 7098
rect 28436 7046 28448 7098
rect 28448 7046 28462 7098
rect 28486 7046 28500 7098
rect 28500 7046 28512 7098
rect 28512 7046 28542 7098
rect 28566 7046 28576 7098
rect 28576 7046 28622 7098
rect 28326 7044 28382 7046
rect 28406 7044 28462 7046
rect 28486 7044 28542 7046
rect 28566 7044 28622 7046
rect 28326 6010 28382 6012
rect 28406 6010 28462 6012
rect 28486 6010 28542 6012
rect 28566 6010 28622 6012
rect 28326 5958 28372 6010
rect 28372 5958 28382 6010
rect 28406 5958 28436 6010
rect 28436 5958 28448 6010
rect 28448 5958 28462 6010
rect 28486 5958 28500 6010
rect 28500 5958 28512 6010
rect 28512 5958 28542 6010
rect 28566 5958 28576 6010
rect 28576 5958 28622 6010
rect 28326 5956 28382 5958
rect 28406 5956 28462 5958
rect 28486 5956 28542 5958
rect 28566 5956 28622 5958
rect 27802 5652 27804 5672
rect 27804 5652 27856 5672
rect 27856 5652 27858 5672
rect 27802 5616 27858 5652
rect 28630 5616 28686 5672
rect 28326 4922 28382 4924
rect 28406 4922 28462 4924
rect 28486 4922 28542 4924
rect 28566 4922 28622 4924
rect 28326 4870 28372 4922
rect 28372 4870 28382 4922
rect 28406 4870 28436 4922
rect 28436 4870 28448 4922
rect 28448 4870 28462 4922
rect 28486 4870 28500 4922
rect 28500 4870 28512 4922
rect 28512 4870 28542 4922
rect 28566 4870 28576 4922
rect 28576 4870 28622 4922
rect 28326 4868 28382 4870
rect 28406 4868 28462 4870
rect 28486 4868 28542 4870
rect 28566 4868 28622 4870
rect 28326 3834 28382 3836
rect 28406 3834 28462 3836
rect 28486 3834 28542 3836
rect 28566 3834 28622 3836
rect 28326 3782 28372 3834
rect 28372 3782 28382 3834
rect 28406 3782 28436 3834
rect 28436 3782 28448 3834
rect 28448 3782 28462 3834
rect 28486 3782 28500 3834
rect 28500 3782 28512 3834
rect 28512 3782 28542 3834
rect 28566 3782 28576 3834
rect 28576 3782 28622 3834
rect 28326 3780 28382 3782
rect 28406 3780 28462 3782
rect 28486 3780 28542 3782
rect 28566 3780 28622 3782
rect 32402 8492 32458 8528
rect 32402 8472 32404 8492
rect 32404 8472 32456 8492
rect 32456 8472 32458 8492
rect 28326 2746 28382 2748
rect 28406 2746 28462 2748
rect 28486 2746 28542 2748
rect 28566 2746 28622 2748
rect 28326 2694 28372 2746
rect 28372 2694 28382 2746
rect 28406 2694 28436 2746
rect 28436 2694 28448 2746
rect 28448 2694 28462 2746
rect 28486 2694 28500 2746
rect 28500 2694 28512 2746
rect 28512 2694 28542 2746
rect 28566 2694 28576 2746
rect 28576 2694 28622 2746
rect 28326 2692 28382 2694
rect 28406 2692 28462 2694
rect 28486 2692 28542 2694
rect 28566 2692 28622 2694
rect 33138 6840 33194 6896
rect 33800 13082 33856 13084
rect 33880 13082 33936 13084
rect 33960 13082 34016 13084
rect 34040 13082 34096 13084
rect 33800 13030 33846 13082
rect 33846 13030 33856 13082
rect 33880 13030 33910 13082
rect 33910 13030 33922 13082
rect 33922 13030 33936 13082
rect 33960 13030 33974 13082
rect 33974 13030 33986 13082
rect 33986 13030 34016 13082
rect 34040 13030 34050 13082
rect 34050 13030 34096 13082
rect 33800 13028 33856 13030
rect 33880 13028 33936 13030
rect 33960 13028 34016 13030
rect 34040 13028 34096 13030
rect 43442 19080 43498 19136
rect 39274 16890 39330 16892
rect 39354 16890 39410 16892
rect 39434 16890 39490 16892
rect 39514 16890 39570 16892
rect 39274 16838 39320 16890
rect 39320 16838 39330 16890
rect 39354 16838 39384 16890
rect 39384 16838 39396 16890
rect 39396 16838 39410 16890
rect 39434 16838 39448 16890
rect 39448 16838 39460 16890
rect 39460 16838 39490 16890
rect 39514 16838 39524 16890
rect 39524 16838 39570 16890
rect 39274 16836 39330 16838
rect 39354 16836 39410 16838
rect 39434 16836 39490 16838
rect 39514 16836 39570 16838
rect 39274 15802 39330 15804
rect 39354 15802 39410 15804
rect 39434 15802 39490 15804
rect 39514 15802 39570 15804
rect 39274 15750 39320 15802
rect 39320 15750 39330 15802
rect 39354 15750 39384 15802
rect 39384 15750 39396 15802
rect 39396 15750 39410 15802
rect 39434 15750 39448 15802
rect 39448 15750 39460 15802
rect 39460 15750 39490 15802
rect 39514 15750 39524 15802
rect 39524 15750 39570 15802
rect 39274 15748 39330 15750
rect 39354 15748 39410 15750
rect 39434 15748 39490 15750
rect 39514 15748 39570 15750
rect 39274 14714 39330 14716
rect 39354 14714 39410 14716
rect 39434 14714 39490 14716
rect 39514 14714 39570 14716
rect 39274 14662 39320 14714
rect 39320 14662 39330 14714
rect 39354 14662 39384 14714
rect 39384 14662 39396 14714
rect 39396 14662 39410 14714
rect 39434 14662 39448 14714
rect 39448 14662 39460 14714
rect 39460 14662 39490 14714
rect 39514 14662 39524 14714
rect 39524 14662 39570 14714
rect 39274 14660 39330 14662
rect 39354 14660 39410 14662
rect 39434 14660 39490 14662
rect 39514 14660 39570 14662
rect 39274 13626 39330 13628
rect 39354 13626 39410 13628
rect 39434 13626 39490 13628
rect 39514 13626 39570 13628
rect 39274 13574 39320 13626
rect 39320 13574 39330 13626
rect 39354 13574 39384 13626
rect 39384 13574 39396 13626
rect 39396 13574 39410 13626
rect 39434 13574 39448 13626
rect 39448 13574 39460 13626
rect 39460 13574 39490 13626
rect 39514 13574 39524 13626
rect 39524 13574 39570 13626
rect 39274 13572 39330 13574
rect 39354 13572 39410 13574
rect 39434 13572 39490 13574
rect 39514 13572 39570 13574
rect 33800 11994 33856 11996
rect 33880 11994 33936 11996
rect 33960 11994 34016 11996
rect 34040 11994 34096 11996
rect 33800 11942 33846 11994
rect 33846 11942 33856 11994
rect 33880 11942 33910 11994
rect 33910 11942 33922 11994
rect 33922 11942 33936 11994
rect 33960 11942 33974 11994
rect 33974 11942 33986 11994
rect 33986 11942 34016 11994
rect 34040 11942 34050 11994
rect 34050 11942 34096 11994
rect 33800 11940 33856 11942
rect 33880 11940 33936 11942
rect 33960 11940 34016 11942
rect 34040 11940 34096 11942
rect 33800 10906 33856 10908
rect 33880 10906 33936 10908
rect 33960 10906 34016 10908
rect 34040 10906 34096 10908
rect 33800 10854 33846 10906
rect 33846 10854 33856 10906
rect 33880 10854 33910 10906
rect 33910 10854 33922 10906
rect 33922 10854 33936 10906
rect 33960 10854 33974 10906
rect 33974 10854 33986 10906
rect 33986 10854 34016 10906
rect 34040 10854 34050 10906
rect 34050 10854 34096 10906
rect 33800 10852 33856 10854
rect 33880 10852 33936 10854
rect 33960 10852 34016 10854
rect 34040 10852 34096 10854
rect 33800 9818 33856 9820
rect 33880 9818 33936 9820
rect 33960 9818 34016 9820
rect 34040 9818 34096 9820
rect 33800 9766 33846 9818
rect 33846 9766 33856 9818
rect 33880 9766 33910 9818
rect 33910 9766 33922 9818
rect 33922 9766 33936 9818
rect 33960 9766 33974 9818
rect 33974 9766 33986 9818
rect 33986 9766 34016 9818
rect 34040 9766 34050 9818
rect 34050 9766 34096 9818
rect 33800 9764 33856 9766
rect 33880 9764 33936 9766
rect 33960 9764 34016 9766
rect 34040 9764 34096 9766
rect 33800 8730 33856 8732
rect 33880 8730 33936 8732
rect 33960 8730 34016 8732
rect 34040 8730 34096 8732
rect 33800 8678 33846 8730
rect 33846 8678 33856 8730
rect 33880 8678 33910 8730
rect 33910 8678 33922 8730
rect 33922 8678 33936 8730
rect 33960 8678 33974 8730
rect 33974 8678 33986 8730
rect 33986 8678 34016 8730
rect 34040 8678 34050 8730
rect 34050 8678 34096 8730
rect 33800 8676 33856 8678
rect 33880 8676 33936 8678
rect 33960 8676 34016 8678
rect 34040 8676 34096 8678
rect 33800 7642 33856 7644
rect 33880 7642 33936 7644
rect 33960 7642 34016 7644
rect 34040 7642 34096 7644
rect 33800 7590 33846 7642
rect 33846 7590 33856 7642
rect 33880 7590 33910 7642
rect 33910 7590 33922 7642
rect 33922 7590 33936 7642
rect 33960 7590 33974 7642
rect 33974 7590 33986 7642
rect 33986 7590 34016 7642
rect 34040 7590 34050 7642
rect 34050 7590 34096 7642
rect 33800 7588 33856 7590
rect 33880 7588 33936 7590
rect 33960 7588 34016 7590
rect 34040 7588 34096 7590
rect 33800 6554 33856 6556
rect 33880 6554 33936 6556
rect 33960 6554 34016 6556
rect 34040 6554 34096 6556
rect 33800 6502 33846 6554
rect 33846 6502 33856 6554
rect 33880 6502 33910 6554
rect 33910 6502 33922 6554
rect 33922 6502 33936 6554
rect 33960 6502 33974 6554
rect 33974 6502 33986 6554
rect 33986 6502 34016 6554
rect 34040 6502 34050 6554
rect 34050 6502 34096 6554
rect 33800 6500 33856 6502
rect 33880 6500 33936 6502
rect 33960 6500 34016 6502
rect 34040 6500 34096 6502
rect 33800 5466 33856 5468
rect 33880 5466 33936 5468
rect 33960 5466 34016 5468
rect 34040 5466 34096 5468
rect 33800 5414 33846 5466
rect 33846 5414 33856 5466
rect 33880 5414 33910 5466
rect 33910 5414 33922 5466
rect 33922 5414 33936 5466
rect 33960 5414 33974 5466
rect 33974 5414 33986 5466
rect 33986 5414 34016 5466
rect 34040 5414 34050 5466
rect 34050 5414 34096 5466
rect 33800 5412 33856 5414
rect 33880 5412 33936 5414
rect 33960 5412 34016 5414
rect 34040 5412 34096 5414
rect 33800 4378 33856 4380
rect 33880 4378 33936 4380
rect 33960 4378 34016 4380
rect 34040 4378 34096 4380
rect 33800 4326 33846 4378
rect 33846 4326 33856 4378
rect 33880 4326 33910 4378
rect 33910 4326 33922 4378
rect 33922 4326 33936 4378
rect 33960 4326 33974 4378
rect 33974 4326 33986 4378
rect 33986 4326 34016 4378
rect 34040 4326 34050 4378
rect 34050 4326 34096 4378
rect 33800 4324 33856 4326
rect 33880 4324 33936 4326
rect 33960 4324 34016 4326
rect 34040 4324 34096 4326
rect 33800 3290 33856 3292
rect 33880 3290 33936 3292
rect 33960 3290 34016 3292
rect 34040 3290 34096 3292
rect 33800 3238 33846 3290
rect 33846 3238 33856 3290
rect 33880 3238 33910 3290
rect 33910 3238 33922 3290
rect 33922 3238 33936 3290
rect 33960 3238 33974 3290
rect 33974 3238 33986 3290
rect 33986 3238 34016 3290
rect 34040 3238 34050 3290
rect 34050 3238 34096 3290
rect 33800 3236 33856 3238
rect 33880 3236 33936 3238
rect 33960 3236 34016 3238
rect 34040 3236 34096 3238
rect 36726 10784 36782 10840
rect 37186 11076 37242 11112
rect 37186 11056 37188 11076
rect 37188 11056 37240 11076
rect 37240 11056 37242 11076
rect 37278 10532 37334 10568
rect 37278 10512 37280 10532
rect 37280 10512 37332 10532
rect 37332 10512 37334 10532
rect 37370 10376 37426 10432
rect 38106 11736 38162 11792
rect 37830 10512 37886 10568
rect 37738 10376 37794 10432
rect 38290 10784 38346 10840
rect 38658 11092 38660 11112
rect 38660 11092 38712 11112
rect 38712 11092 38714 11112
rect 38658 11056 38714 11092
rect 39274 12538 39330 12540
rect 39354 12538 39410 12540
rect 39434 12538 39490 12540
rect 39514 12538 39570 12540
rect 39274 12486 39320 12538
rect 39320 12486 39330 12538
rect 39354 12486 39384 12538
rect 39384 12486 39396 12538
rect 39396 12486 39410 12538
rect 39434 12486 39448 12538
rect 39448 12486 39460 12538
rect 39460 12486 39490 12538
rect 39514 12486 39524 12538
rect 39524 12486 39570 12538
rect 39274 12484 39330 12486
rect 39354 12484 39410 12486
rect 39434 12484 39490 12486
rect 39514 12484 39570 12486
rect 39274 11450 39330 11452
rect 39354 11450 39410 11452
rect 39434 11450 39490 11452
rect 39514 11450 39570 11452
rect 39274 11398 39320 11450
rect 39320 11398 39330 11450
rect 39354 11398 39384 11450
rect 39384 11398 39396 11450
rect 39396 11398 39410 11450
rect 39434 11398 39448 11450
rect 39448 11398 39460 11450
rect 39460 11398 39490 11450
rect 39514 11398 39524 11450
rect 39524 11398 39570 11450
rect 39274 11396 39330 11398
rect 39354 11396 39410 11398
rect 39434 11396 39490 11398
rect 39514 11396 39570 11398
rect 36174 8472 36230 8528
rect 39274 10362 39330 10364
rect 39354 10362 39410 10364
rect 39434 10362 39490 10364
rect 39514 10362 39570 10364
rect 39274 10310 39320 10362
rect 39320 10310 39330 10362
rect 39354 10310 39384 10362
rect 39384 10310 39396 10362
rect 39396 10310 39410 10362
rect 39434 10310 39448 10362
rect 39448 10310 39460 10362
rect 39460 10310 39490 10362
rect 39514 10310 39524 10362
rect 39524 10310 39570 10362
rect 39274 10308 39330 10310
rect 39354 10308 39410 10310
rect 39434 10308 39490 10310
rect 39514 10308 39570 10310
rect 39670 9596 39672 9616
rect 39672 9596 39724 9616
rect 39724 9596 39726 9616
rect 39670 9560 39726 9596
rect 39274 9274 39330 9276
rect 39354 9274 39410 9276
rect 39434 9274 39490 9276
rect 39514 9274 39570 9276
rect 39274 9222 39320 9274
rect 39320 9222 39330 9274
rect 39354 9222 39384 9274
rect 39384 9222 39396 9274
rect 39396 9222 39410 9274
rect 39434 9222 39448 9274
rect 39448 9222 39460 9274
rect 39460 9222 39490 9274
rect 39514 9222 39524 9274
rect 39524 9222 39570 9274
rect 39274 9220 39330 9222
rect 39354 9220 39410 9222
rect 39434 9220 39490 9222
rect 39514 9220 39570 9222
rect 39210 9016 39266 9072
rect 40314 11464 40370 11520
rect 40314 10104 40370 10160
rect 40314 10004 40316 10024
rect 40316 10004 40368 10024
rect 40368 10004 40370 10024
rect 40314 9968 40370 10004
rect 39274 8186 39330 8188
rect 39354 8186 39410 8188
rect 39434 8186 39490 8188
rect 39514 8186 39570 8188
rect 39274 8134 39320 8186
rect 39320 8134 39330 8186
rect 39354 8134 39384 8186
rect 39384 8134 39396 8186
rect 39396 8134 39410 8186
rect 39434 8134 39448 8186
rect 39448 8134 39460 8186
rect 39460 8134 39490 8186
rect 39514 8134 39524 8186
rect 39524 8134 39570 8186
rect 39274 8132 39330 8134
rect 39354 8132 39410 8134
rect 39434 8132 39490 8134
rect 39514 8132 39570 8134
rect 39274 7098 39330 7100
rect 39354 7098 39410 7100
rect 39434 7098 39490 7100
rect 39514 7098 39570 7100
rect 39274 7046 39320 7098
rect 39320 7046 39330 7098
rect 39354 7046 39384 7098
rect 39384 7046 39396 7098
rect 39396 7046 39410 7098
rect 39434 7046 39448 7098
rect 39448 7046 39460 7098
rect 39460 7046 39490 7098
rect 39514 7046 39524 7098
rect 39524 7046 39570 7098
rect 39274 7044 39330 7046
rect 39354 7044 39410 7046
rect 39434 7044 39490 7046
rect 39514 7044 39570 7046
rect 40222 9016 40278 9072
rect 40682 9832 40738 9888
rect 41142 10004 41144 10024
rect 41144 10004 41196 10024
rect 41196 10004 41198 10024
rect 41142 9968 41198 10004
rect 41326 10104 41382 10160
rect 42062 11464 42118 11520
rect 44086 17720 44142 17776
rect 44748 17434 44804 17436
rect 44828 17434 44884 17436
rect 44908 17434 44964 17436
rect 44988 17434 45044 17436
rect 44748 17382 44794 17434
rect 44794 17382 44804 17434
rect 44828 17382 44858 17434
rect 44858 17382 44870 17434
rect 44870 17382 44884 17434
rect 44908 17382 44922 17434
rect 44922 17382 44934 17434
rect 44934 17382 44964 17434
rect 44988 17382 44998 17434
rect 44998 17382 45044 17434
rect 44748 17380 44804 17382
rect 44828 17380 44884 17382
rect 44908 17380 44964 17382
rect 44988 17380 45044 17382
rect 44748 16346 44804 16348
rect 44828 16346 44884 16348
rect 44908 16346 44964 16348
rect 44988 16346 45044 16348
rect 44748 16294 44794 16346
rect 44794 16294 44804 16346
rect 44828 16294 44858 16346
rect 44858 16294 44870 16346
rect 44870 16294 44884 16346
rect 44908 16294 44922 16346
rect 44922 16294 44934 16346
rect 44934 16294 44964 16346
rect 44988 16294 44998 16346
rect 44998 16294 45044 16346
rect 44748 16292 44804 16294
rect 44828 16292 44884 16294
rect 44908 16292 44964 16294
rect 44988 16292 45044 16294
rect 44178 15680 44234 15736
rect 44748 15258 44804 15260
rect 44828 15258 44884 15260
rect 44908 15258 44964 15260
rect 44988 15258 45044 15260
rect 44748 15206 44794 15258
rect 44794 15206 44804 15258
rect 44828 15206 44858 15258
rect 44858 15206 44870 15258
rect 44870 15206 44884 15258
rect 44908 15206 44922 15258
rect 44922 15206 44934 15258
rect 44934 15206 44964 15258
rect 44988 15206 44998 15258
rect 44998 15206 45044 15258
rect 44748 15204 44804 15206
rect 44828 15204 44884 15206
rect 44908 15204 44964 15206
rect 44988 15204 45044 15206
rect 44086 14320 44142 14376
rect 44748 14170 44804 14172
rect 44828 14170 44884 14172
rect 44908 14170 44964 14172
rect 44988 14170 45044 14172
rect 44748 14118 44794 14170
rect 44794 14118 44804 14170
rect 44828 14118 44858 14170
rect 44858 14118 44870 14170
rect 44870 14118 44884 14170
rect 44908 14118 44922 14170
rect 44922 14118 44934 14170
rect 44934 14118 44964 14170
rect 44988 14118 44998 14170
rect 44998 14118 45044 14170
rect 44748 14116 44804 14118
rect 44828 14116 44884 14118
rect 44908 14116 44964 14118
rect 44988 14116 45044 14118
rect 44748 13082 44804 13084
rect 44828 13082 44884 13084
rect 44908 13082 44964 13084
rect 44988 13082 45044 13084
rect 44748 13030 44794 13082
rect 44794 13030 44804 13082
rect 44828 13030 44858 13082
rect 44858 13030 44870 13082
rect 44870 13030 44884 13082
rect 44908 13030 44922 13082
rect 44922 13030 44934 13082
rect 44934 13030 44964 13082
rect 44988 13030 44998 13082
rect 44998 13030 45044 13082
rect 44748 13028 44804 13030
rect 44828 13028 44884 13030
rect 44908 13028 44964 13030
rect 44988 13028 45044 13030
rect 44086 12280 44142 12336
rect 44748 11994 44804 11996
rect 44828 11994 44884 11996
rect 44908 11994 44964 11996
rect 44988 11994 45044 11996
rect 44748 11942 44794 11994
rect 44794 11942 44804 11994
rect 44828 11942 44858 11994
rect 44858 11942 44870 11994
rect 44870 11942 44884 11994
rect 44908 11942 44922 11994
rect 44922 11942 44934 11994
rect 44934 11942 44964 11994
rect 44988 11942 44998 11994
rect 44998 11942 45044 11994
rect 44748 11940 44804 11942
rect 44828 11940 44884 11942
rect 44908 11940 44964 11942
rect 44988 11940 45044 11942
rect 44748 10906 44804 10908
rect 44828 10906 44884 10908
rect 44908 10906 44964 10908
rect 44988 10906 45044 10908
rect 44748 10854 44794 10906
rect 44794 10854 44804 10906
rect 44828 10854 44858 10906
rect 44858 10854 44870 10906
rect 44870 10854 44884 10906
rect 44908 10854 44922 10906
rect 44922 10854 44934 10906
rect 44934 10854 44964 10906
rect 44988 10854 44998 10906
rect 44998 10854 45044 10906
rect 44748 10852 44804 10854
rect 44828 10852 44884 10854
rect 44908 10852 44964 10854
rect 44988 10852 45044 10854
rect 44178 10668 44234 10704
rect 44178 10648 44180 10668
rect 44180 10648 44232 10668
rect 44232 10648 44234 10668
rect 41694 9832 41750 9888
rect 40958 9580 41014 9616
rect 40958 9560 40960 9580
rect 40960 9560 41012 9580
rect 41012 9560 41014 9580
rect 44748 9818 44804 9820
rect 44828 9818 44884 9820
rect 44908 9818 44964 9820
rect 44988 9818 45044 9820
rect 44748 9766 44794 9818
rect 44794 9766 44804 9818
rect 44828 9766 44858 9818
rect 44858 9766 44870 9818
rect 44870 9766 44884 9818
rect 44908 9766 44922 9818
rect 44922 9766 44934 9818
rect 44934 9766 44964 9818
rect 44988 9766 44998 9818
rect 44998 9766 45044 9818
rect 44748 9764 44804 9766
rect 44828 9764 44884 9766
rect 44908 9764 44964 9766
rect 44988 9764 45044 9766
rect 39274 6010 39330 6012
rect 39354 6010 39410 6012
rect 39434 6010 39490 6012
rect 39514 6010 39570 6012
rect 39274 5958 39320 6010
rect 39320 5958 39330 6010
rect 39354 5958 39384 6010
rect 39384 5958 39396 6010
rect 39396 5958 39410 6010
rect 39434 5958 39448 6010
rect 39448 5958 39460 6010
rect 39460 5958 39490 6010
rect 39514 5958 39524 6010
rect 39524 5958 39570 6010
rect 39274 5956 39330 5958
rect 39354 5956 39410 5958
rect 39434 5956 39490 5958
rect 39514 5956 39570 5958
rect 39274 4922 39330 4924
rect 39354 4922 39410 4924
rect 39434 4922 39490 4924
rect 39514 4922 39570 4924
rect 39274 4870 39320 4922
rect 39320 4870 39330 4922
rect 39354 4870 39384 4922
rect 39384 4870 39396 4922
rect 39396 4870 39410 4922
rect 39434 4870 39448 4922
rect 39448 4870 39460 4922
rect 39460 4870 39490 4922
rect 39514 4870 39524 4922
rect 39524 4870 39570 4922
rect 39274 4868 39330 4870
rect 39354 4868 39410 4870
rect 39434 4868 39490 4870
rect 39514 4868 39570 4870
rect 39274 3834 39330 3836
rect 39354 3834 39410 3836
rect 39434 3834 39490 3836
rect 39514 3834 39570 3836
rect 39274 3782 39320 3834
rect 39320 3782 39330 3834
rect 39354 3782 39384 3834
rect 39384 3782 39396 3834
rect 39396 3782 39410 3834
rect 39434 3782 39448 3834
rect 39448 3782 39460 3834
rect 39460 3782 39490 3834
rect 39514 3782 39524 3834
rect 39524 3782 39570 3834
rect 39274 3780 39330 3782
rect 39354 3780 39410 3782
rect 39434 3780 39490 3782
rect 39514 3780 39570 3782
rect 44178 8880 44234 8936
rect 44748 8730 44804 8732
rect 44828 8730 44884 8732
rect 44908 8730 44964 8732
rect 44988 8730 45044 8732
rect 44748 8678 44794 8730
rect 44794 8678 44804 8730
rect 44828 8678 44858 8730
rect 44858 8678 44870 8730
rect 44870 8678 44884 8730
rect 44908 8678 44922 8730
rect 44922 8678 44934 8730
rect 44934 8678 44964 8730
rect 44988 8678 44998 8730
rect 44998 8678 45044 8730
rect 44748 8676 44804 8678
rect 44828 8676 44884 8678
rect 44908 8676 44964 8678
rect 44988 8676 45044 8678
rect 44178 7828 44180 7848
rect 44180 7828 44232 7848
rect 44232 7828 44234 7848
rect 44178 7792 44234 7828
rect 44748 7642 44804 7644
rect 44828 7642 44884 7644
rect 44908 7642 44964 7644
rect 44988 7642 45044 7644
rect 44748 7590 44794 7642
rect 44794 7590 44804 7642
rect 44828 7590 44858 7642
rect 44858 7590 44870 7642
rect 44870 7590 44884 7642
rect 44908 7590 44922 7642
rect 44922 7590 44934 7642
rect 44934 7590 44964 7642
rect 44988 7590 44998 7642
rect 44998 7590 45044 7642
rect 44748 7588 44804 7590
rect 44828 7588 44884 7590
rect 44908 7588 44964 7590
rect 44988 7588 45044 7590
rect 44748 6554 44804 6556
rect 44828 6554 44884 6556
rect 44908 6554 44964 6556
rect 44988 6554 45044 6556
rect 44748 6502 44794 6554
rect 44794 6502 44804 6554
rect 44828 6502 44858 6554
rect 44858 6502 44870 6554
rect 44870 6502 44884 6554
rect 44908 6502 44922 6554
rect 44922 6502 44934 6554
rect 44934 6502 44964 6554
rect 44988 6502 44998 6554
rect 44998 6502 45044 6554
rect 44748 6500 44804 6502
rect 44828 6500 44884 6502
rect 44908 6500 44964 6502
rect 44988 6500 45044 6502
rect 44748 5466 44804 5468
rect 44828 5466 44884 5468
rect 44908 5466 44964 5468
rect 44988 5466 45044 5468
rect 44748 5414 44794 5466
rect 44794 5414 44804 5466
rect 44828 5414 44858 5466
rect 44858 5414 44870 5466
rect 44870 5414 44884 5466
rect 44908 5414 44922 5466
rect 44922 5414 44934 5466
rect 44934 5414 44964 5466
rect 44988 5414 44998 5466
rect 44998 5414 45044 5466
rect 44748 5412 44804 5414
rect 44828 5412 44884 5414
rect 44908 5412 44964 5414
rect 44988 5412 45044 5414
rect 44086 5208 44142 5264
rect 44748 4378 44804 4380
rect 44828 4378 44884 4380
rect 44908 4378 44964 4380
rect 44988 4378 45044 4380
rect 44748 4326 44794 4378
rect 44794 4326 44804 4378
rect 44828 4326 44858 4378
rect 44858 4326 44870 4378
rect 44870 4326 44884 4378
rect 44908 4326 44922 4378
rect 44922 4326 44934 4378
rect 44934 4326 44964 4378
rect 44988 4326 44998 4378
rect 44998 4326 45044 4378
rect 44748 4324 44804 4326
rect 44828 4324 44884 4326
rect 44908 4324 44964 4326
rect 44988 4324 45044 4326
rect 44086 4120 44142 4176
rect 39274 2746 39330 2748
rect 39354 2746 39410 2748
rect 39434 2746 39490 2748
rect 39514 2746 39570 2748
rect 39274 2694 39320 2746
rect 39320 2694 39330 2746
rect 39354 2694 39384 2746
rect 39384 2694 39396 2746
rect 39396 2694 39410 2746
rect 39434 2694 39448 2746
rect 39448 2694 39460 2746
rect 39460 2694 39490 2746
rect 39514 2694 39524 2746
rect 39524 2694 39570 2746
rect 39274 2692 39330 2694
rect 39354 2692 39410 2694
rect 39434 2692 39490 2694
rect 39514 2692 39570 2694
rect 33800 2202 33856 2204
rect 33880 2202 33936 2204
rect 33960 2202 34016 2204
rect 34040 2202 34096 2204
rect 33800 2150 33846 2202
rect 33846 2150 33856 2202
rect 33880 2150 33910 2202
rect 33910 2150 33922 2202
rect 33922 2150 33936 2202
rect 33960 2150 33974 2202
rect 33974 2150 33986 2202
rect 33986 2150 34016 2202
rect 34040 2150 34050 2202
rect 34050 2150 34096 2202
rect 33800 2148 33856 2150
rect 33880 2148 33936 2150
rect 33960 2148 34016 2150
rect 34040 2148 34096 2150
rect 44086 2352 44142 2408
rect 44748 3290 44804 3292
rect 44828 3290 44884 3292
rect 44908 3290 44964 3292
rect 44988 3290 45044 3292
rect 44748 3238 44794 3290
rect 44794 3238 44804 3290
rect 44828 3238 44858 3290
rect 44858 3238 44870 3290
rect 44870 3238 44884 3290
rect 44908 3238 44922 3290
rect 44922 3238 44934 3290
rect 44934 3238 44964 3290
rect 44988 3238 44998 3290
rect 44998 3238 45044 3290
rect 44748 3236 44804 3238
rect 44828 3236 44884 3238
rect 44908 3236 44964 3238
rect 44988 3236 45044 3238
rect 44748 2202 44804 2204
rect 44828 2202 44884 2204
rect 44908 2202 44964 2204
rect 44988 2202 45044 2204
rect 44748 2150 44794 2202
rect 44794 2150 44804 2202
rect 44828 2150 44858 2202
rect 44858 2150 44870 2202
rect 44870 2150 44884 2202
rect 44908 2150 44922 2202
rect 44922 2150 44934 2202
rect 44934 2150 44964 2202
rect 44988 2150 44998 2202
rect 44998 2150 45044 2202
rect 44748 2148 44804 2150
rect 44828 2148 44884 2150
rect 44908 2148 44964 2150
rect 44988 2148 45044 2150
rect 44178 720 44234 776
<< metal3 >>
rect 43437 19138 43503 19141
rect 45200 19138 46000 19228
rect 43437 19136 46000 19138
rect 43437 19080 43442 19136
rect 43498 19080 46000 19136
rect 43437 19078 46000 19080
rect 43437 19075 43503 19078
rect 45200 18988 46000 19078
rect 0 18458 800 18548
rect 3969 18458 4035 18461
rect 0 18456 4035 18458
rect 0 18400 3974 18456
rect 4030 18400 4035 18456
rect 0 18398 4035 18400
rect 0 18308 800 18398
rect 3969 18395 4035 18398
rect 44081 17778 44147 17781
rect 45200 17778 46000 17868
rect 44081 17776 46000 17778
rect 44081 17720 44086 17776
rect 44142 17720 46000 17776
rect 44081 17718 46000 17720
rect 44081 17715 44147 17718
rect 45200 17628 46000 17718
rect 11894 17440 12210 17441
rect 11894 17376 11900 17440
rect 11964 17376 11980 17440
rect 12044 17376 12060 17440
rect 12124 17376 12140 17440
rect 12204 17376 12210 17440
rect 11894 17375 12210 17376
rect 22842 17440 23158 17441
rect 22842 17376 22848 17440
rect 22912 17376 22928 17440
rect 22992 17376 23008 17440
rect 23072 17376 23088 17440
rect 23152 17376 23158 17440
rect 22842 17375 23158 17376
rect 33790 17440 34106 17441
rect 33790 17376 33796 17440
rect 33860 17376 33876 17440
rect 33940 17376 33956 17440
rect 34020 17376 34036 17440
rect 34100 17376 34106 17440
rect 33790 17375 34106 17376
rect 44738 17440 45054 17441
rect 44738 17376 44744 17440
rect 44808 17376 44824 17440
rect 44888 17376 44904 17440
rect 44968 17376 44984 17440
rect 45048 17376 45054 17440
rect 44738 17375 45054 17376
rect 0 17098 800 17188
rect 2221 17098 2287 17101
rect 0 17096 2287 17098
rect 0 17040 2226 17096
rect 2282 17040 2287 17096
rect 0 17038 2287 17040
rect 0 16948 800 17038
rect 2221 17035 2287 17038
rect 6420 16896 6736 16897
rect 6420 16832 6426 16896
rect 6490 16832 6506 16896
rect 6570 16832 6586 16896
rect 6650 16832 6666 16896
rect 6730 16832 6736 16896
rect 6420 16831 6736 16832
rect 17368 16896 17684 16897
rect 17368 16832 17374 16896
rect 17438 16832 17454 16896
rect 17518 16832 17534 16896
rect 17598 16832 17614 16896
rect 17678 16832 17684 16896
rect 17368 16831 17684 16832
rect 28316 16896 28632 16897
rect 28316 16832 28322 16896
rect 28386 16832 28402 16896
rect 28466 16832 28482 16896
rect 28546 16832 28562 16896
rect 28626 16832 28632 16896
rect 28316 16831 28632 16832
rect 39264 16896 39580 16897
rect 39264 16832 39270 16896
rect 39334 16832 39350 16896
rect 39414 16832 39430 16896
rect 39494 16832 39510 16896
rect 39574 16832 39580 16896
rect 39264 16831 39580 16832
rect 11894 16352 12210 16353
rect 11894 16288 11900 16352
rect 11964 16288 11980 16352
rect 12044 16288 12060 16352
rect 12124 16288 12140 16352
rect 12204 16288 12210 16352
rect 11894 16287 12210 16288
rect 22842 16352 23158 16353
rect 22842 16288 22848 16352
rect 22912 16288 22928 16352
rect 22992 16288 23008 16352
rect 23072 16288 23088 16352
rect 23152 16288 23158 16352
rect 22842 16287 23158 16288
rect 33790 16352 34106 16353
rect 33790 16288 33796 16352
rect 33860 16288 33876 16352
rect 33940 16288 33956 16352
rect 34020 16288 34036 16352
rect 34100 16288 34106 16352
rect 33790 16287 34106 16288
rect 44738 16352 45054 16353
rect 44738 16288 44744 16352
rect 44808 16288 44824 16352
rect 44888 16288 44904 16352
rect 44968 16288 44984 16352
rect 45048 16288 45054 16352
rect 44738 16287 45054 16288
rect 6420 15808 6736 15809
rect 6420 15744 6426 15808
rect 6490 15744 6506 15808
rect 6570 15744 6586 15808
rect 6650 15744 6666 15808
rect 6730 15744 6736 15808
rect 6420 15743 6736 15744
rect 17368 15808 17684 15809
rect 17368 15744 17374 15808
rect 17438 15744 17454 15808
rect 17518 15744 17534 15808
rect 17598 15744 17614 15808
rect 17678 15744 17684 15808
rect 17368 15743 17684 15744
rect 28316 15808 28632 15809
rect 28316 15744 28322 15808
rect 28386 15744 28402 15808
rect 28466 15744 28482 15808
rect 28546 15744 28562 15808
rect 28626 15744 28632 15808
rect 28316 15743 28632 15744
rect 39264 15808 39580 15809
rect 39264 15744 39270 15808
rect 39334 15744 39350 15808
rect 39414 15744 39430 15808
rect 39494 15744 39510 15808
rect 39574 15744 39580 15808
rect 39264 15743 39580 15744
rect 44173 15738 44239 15741
rect 45200 15738 46000 15828
rect 44173 15736 46000 15738
rect 44173 15680 44178 15736
rect 44234 15680 46000 15736
rect 44173 15678 46000 15680
rect 44173 15675 44239 15678
rect 45200 15588 46000 15678
rect 11894 15264 12210 15265
rect 11894 15200 11900 15264
rect 11964 15200 11980 15264
rect 12044 15200 12060 15264
rect 12124 15200 12140 15264
rect 12204 15200 12210 15264
rect 11894 15199 12210 15200
rect 22842 15264 23158 15265
rect 22842 15200 22848 15264
rect 22912 15200 22928 15264
rect 22992 15200 23008 15264
rect 23072 15200 23088 15264
rect 23152 15200 23158 15264
rect 22842 15199 23158 15200
rect 33790 15264 34106 15265
rect 33790 15200 33796 15264
rect 33860 15200 33876 15264
rect 33940 15200 33956 15264
rect 34020 15200 34036 15264
rect 34100 15200 34106 15264
rect 33790 15199 34106 15200
rect 44738 15264 45054 15265
rect 44738 15200 44744 15264
rect 44808 15200 44824 15264
rect 44888 15200 44904 15264
rect 44968 15200 44984 15264
rect 45048 15200 45054 15264
rect 44738 15199 45054 15200
rect 0 15058 800 15148
rect 1577 15058 1643 15061
rect 0 15056 1643 15058
rect 0 15000 1582 15056
rect 1638 15000 1643 15056
rect 0 14998 1643 15000
rect 0 14908 800 14998
rect 1577 14995 1643 14998
rect 6420 14720 6736 14721
rect 6420 14656 6426 14720
rect 6490 14656 6506 14720
rect 6570 14656 6586 14720
rect 6650 14656 6666 14720
rect 6730 14656 6736 14720
rect 6420 14655 6736 14656
rect 17368 14720 17684 14721
rect 17368 14656 17374 14720
rect 17438 14656 17454 14720
rect 17518 14656 17534 14720
rect 17598 14656 17614 14720
rect 17678 14656 17684 14720
rect 17368 14655 17684 14656
rect 28316 14720 28632 14721
rect 28316 14656 28322 14720
rect 28386 14656 28402 14720
rect 28466 14656 28482 14720
rect 28546 14656 28562 14720
rect 28626 14656 28632 14720
rect 28316 14655 28632 14656
rect 39264 14720 39580 14721
rect 39264 14656 39270 14720
rect 39334 14656 39350 14720
rect 39414 14656 39430 14720
rect 39494 14656 39510 14720
rect 39574 14656 39580 14720
rect 39264 14655 39580 14656
rect 44081 14378 44147 14381
rect 45200 14378 46000 14468
rect 44081 14376 46000 14378
rect 44081 14320 44086 14376
rect 44142 14320 46000 14376
rect 44081 14318 46000 14320
rect 44081 14315 44147 14318
rect 45200 14228 46000 14318
rect 11894 14176 12210 14177
rect 11894 14112 11900 14176
rect 11964 14112 11980 14176
rect 12044 14112 12060 14176
rect 12124 14112 12140 14176
rect 12204 14112 12210 14176
rect 11894 14111 12210 14112
rect 22842 14176 23158 14177
rect 22842 14112 22848 14176
rect 22912 14112 22928 14176
rect 22992 14112 23008 14176
rect 23072 14112 23088 14176
rect 23152 14112 23158 14176
rect 22842 14111 23158 14112
rect 33790 14176 34106 14177
rect 33790 14112 33796 14176
rect 33860 14112 33876 14176
rect 33940 14112 33956 14176
rect 34020 14112 34036 14176
rect 34100 14112 34106 14176
rect 33790 14111 34106 14112
rect 44738 14176 45054 14177
rect 44738 14112 44744 14176
rect 44808 14112 44824 14176
rect 44888 14112 44904 14176
rect 44968 14112 44984 14176
rect 45048 14112 45054 14176
rect 44738 14111 45054 14112
rect 0 13698 800 13788
rect 1577 13698 1643 13701
rect 0 13696 1643 13698
rect 0 13640 1582 13696
rect 1638 13640 1643 13696
rect 0 13638 1643 13640
rect 0 13548 800 13638
rect 1577 13635 1643 13638
rect 6420 13632 6736 13633
rect 6420 13568 6426 13632
rect 6490 13568 6506 13632
rect 6570 13568 6586 13632
rect 6650 13568 6666 13632
rect 6730 13568 6736 13632
rect 6420 13567 6736 13568
rect 17368 13632 17684 13633
rect 17368 13568 17374 13632
rect 17438 13568 17454 13632
rect 17518 13568 17534 13632
rect 17598 13568 17614 13632
rect 17678 13568 17684 13632
rect 17368 13567 17684 13568
rect 28316 13632 28632 13633
rect 28316 13568 28322 13632
rect 28386 13568 28402 13632
rect 28466 13568 28482 13632
rect 28546 13568 28562 13632
rect 28626 13568 28632 13632
rect 28316 13567 28632 13568
rect 39264 13632 39580 13633
rect 39264 13568 39270 13632
rect 39334 13568 39350 13632
rect 39414 13568 39430 13632
rect 39494 13568 39510 13632
rect 39574 13568 39580 13632
rect 39264 13567 39580 13568
rect 11894 13088 12210 13089
rect 11894 13024 11900 13088
rect 11964 13024 11980 13088
rect 12044 13024 12060 13088
rect 12124 13024 12140 13088
rect 12204 13024 12210 13088
rect 11894 13023 12210 13024
rect 22842 13088 23158 13089
rect 22842 13024 22848 13088
rect 22912 13024 22928 13088
rect 22992 13024 23008 13088
rect 23072 13024 23088 13088
rect 23152 13024 23158 13088
rect 22842 13023 23158 13024
rect 33790 13088 34106 13089
rect 33790 13024 33796 13088
rect 33860 13024 33876 13088
rect 33940 13024 33956 13088
rect 34020 13024 34036 13088
rect 34100 13024 34106 13088
rect 33790 13023 34106 13024
rect 44738 13088 45054 13089
rect 44738 13024 44744 13088
rect 44808 13024 44824 13088
rect 44888 13024 44904 13088
rect 44968 13024 44984 13088
rect 45048 13024 45054 13088
rect 44738 13023 45054 13024
rect 6420 12544 6736 12545
rect 6420 12480 6426 12544
rect 6490 12480 6506 12544
rect 6570 12480 6586 12544
rect 6650 12480 6666 12544
rect 6730 12480 6736 12544
rect 6420 12479 6736 12480
rect 17368 12544 17684 12545
rect 17368 12480 17374 12544
rect 17438 12480 17454 12544
rect 17518 12480 17534 12544
rect 17598 12480 17614 12544
rect 17678 12480 17684 12544
rect 17368 12479 17684 12480
rect 28316 12544 28632 12545
rect 28316 12480 28322 12544
rect 28386 12480 28402 12544
rect 28466 12480 28482 12544
rect 28546 12480 28562 12544
rect 28626 12480 28632 12544
rect 28316 12479 28632 12480
rect 39264 12544 39580 12545
rect 39264 12480 39270 12544
rect 39334 12480 39350 12544
rect 39414 12480 39430 12544
rect 39494 12480 39510 12544
rect 39574 12480 39580 12544
rect 39264 12479 39580 12480
rect 44081 12338 44147 12341
rect 45200 12338 46000 12428
rect 44081 12336 46000 12338
rect 44081 12280 44086 12336
rect 44142 12280 46000 12336
rect 44081 12278 46000 12280
rect 44081 12275 44147 12278
rect 12065 12202 12131 12205
rect 18321 12202 18387 12205
rect 12065 12200 18387 12202
rect 12065 12144 12070 12200
rect 12126 12144 18326 12200
rect 18382 12144 18387 12200
rect 45200 12188 46000 12278
rect 12065 12142 18387 12144
rect 12065 12139 12131 12142
rect 18321 12139 18387 12142
rect 11894 12000 12210 12001
rect 11894 11936 11900 12000
rect 11964 11936 11980 12000
rect 12044 11936 12060 12000
rect 12124 11936 12140 12000
rect 12204 11936 12210 12000
rect 11894 11935 12210 11936
rect 22842 12000 23158 12001
rect 22842 11936 22848 12000
rect 22912 11936 22928 12000
rect 22992 11936 23008 12000
rect 23072 11936 23088 12000
rect 23152 11936 23158 12000
rect 22842 11935 23158 11936
rect 33790 12000 34106 12001
rect 33790 11936 33796 12000
rect 33860 11936 33876 12000
rect 33940 11936 33956 12000
rect 34020 11936 34036 12000
rect 34100 11936 34106 12000
rect 33790 11935 34106 11936
rect 44738 12000 45054 12001
rect 44738 11936 44744 12000
rect 44808 11936 44824 12000
rect 44888 11936 44904 12000
rect 44968 11936 44984 12000
rect 45048 11936 45054 12000
rect 44738 11935 45054 11936
rect 13445 11794 13511 11797
rect 15469 11794 15535 11797
rect 19241 11794 19307 11797
rect 13445 11792 19307 11794
rect 0 11658 800 11748
rect 13445 11736 13450 11792
rect 13506 11736 15474 11792
rect 15530 11736 19246 11792
rect 19302 11736 19307 11792
rect 13445 11734 19307 11736
rect 13445 11731 13511 11734
rect 15469 11731 15535 11734
rect 19241 11731 19307 11734
rect 29453 11794 29519 11797
rect 38101 11794 38167 11797
rect 29453 11792 38167 11794
rect 29453 11736 29458 11792
rect 29514 11736 38106 11792
rect 38162 11736 38167 11792
rect 29453 11734 38167 11736
rect 29453 11731 29519 11734
rect 38101 11731 38167 11734
rect 4061 11658 4127 11661
rect 0 11656 4127 11658
rect 0 11600 4066 11656
rect 4122 11600 4127 11656
rect 0 11598 4127 11600
rect 0 11508 800 11598
rect 4061 11595 4127 11598
rect 40309 11522 40375 11525
rect 42057 11522 42123 11525
rect 40309 11520 42123 11522
rect 40309 11464 40314 11520
rect 40370 11464 42062 11520
rect 42118 11464 42123 11520
rect 40309 11462 42123 11464
rect 40309 11459 40375 11462
rect 42057 11459 42123 11462
rect 6420 11456 6736 11457
rect 6420 11392 6426 11456
rect 6490 11392 6506 11456
rect 6570 11392 6586 11456
rect 6650 11392 6666 11456
rect 6730 11392 6736 11456
rect 6420 11391 6736 11392
rect 17368 11456 17684 11457
rect 17368 11392 17374 11456
rect 17438 11392 17454 11456
rect 17518 11392 17534 11456
rect 17598 11392 17614 11456
rect 17678 11392 17684 11456
rect 17368 11391 17684 11392
rect 28316 11456 28632 11457
rect 28316 11392 28322 11456
rect 28386 11392 28402 11456
rect 28466 11392 28482 11456
rect 28546 11392 28562 11456
rect 28626 11392 28632 11456
rect 28316 11391 28632 11392
rect 39264 11456 39580 11457
rect 39264 11392 39270 11456
rect 39334 11392 39350 11456
rect 39414 11392 39430 11456
rect 39494 11392 39510 11456
rect 39574 11392 39580 11456
rect 39264 11391 39580 11392
rect 37181 11114 37247 11117
rect 38653 11114 38719 11117
rect 37181 11112 38719 11114
rect 37181 11056 37186 11112
rect 37242 11056 38658 11112
rect 38714 11056 38719 11112
rect 37181 11054 38719 11056
rect 37181 11051 37247 11054
rect 38653 11051 38719 11054
rect 45200 10978 46000 11068
rect 11894 10912 12210 10913
rect 11894 10848 11900 10912
rect 11964 10848 11980 10912
rect 12044 10848 12060 10912
rect 12124 10848 12140 10912
rect 12204 10848 12210 10912
rect 11894 10847 12210 10848
rect 22842 10912 23158 10913
rect 22842 10848 22848 10912
rect 22912 10848 22928 10912
rect 22992 10848 23008 10912
rect 23072 10848 23088 10912
rect 23152 10848 23158 10912
rect 22842 10847 23158 10848
rect 33790 10912 34106 10913
rect 33790 10848 33796 10912
rect 33860 10848 33876 10912
rect 33940 10848 33956 10912
rect 34020 10848 34036 10912
rect 34100 10848 34106 10912
rect 33790 10847 34106 10848
rect 44738 10912 45054 10913
rect 44738 10848 44744 10912
rect 44808 10848 44824 10912
rect 44888 10848 44904 10912
rect 44968 10848 44984 10912
rect 45048 10848 45054 10912
rect 44738 10847 45054 10848
rect 36721 10842 36787 10845
rect 38285 10842 38351 10845
rect 36721 10840 38351 10842
rect 36721 10784 36726 10840
rect 36782 10784 38290 10840
rect 38346 10784 38351 10840
rect 36721 10782 38351 10784
rect 36721 10779 36787 10782
rect 38285 10779 38351 10782
rect 45142 10828 46000 10978
rect 22001 10706 22067 10709
rect 25773 10706 25839 10709
rect 22001 10704 25839 10706
rect 22001 10648 22006 10704
rect 22062 10648 25778 10704
rect 25834 10648 25839 10704
rect 22001 10646 25839 10648
rect 22001 10643 22067 10646
rect 25773 10643 25839 10646
rect 44173 10706 44239 10709
rect 45142 10706 45202 10828
rect 44173 10704 45202 10706
rect 44173 10648 44178 10704
rect 44234 10648 45202 10704
rect 44173 10646 45202 10648
rect 44173 10643 44239 10646
rect 37273 10570 37339 10573
rect 37825 10570 37891 10573
rect 37273 10568 37891 10570
rect 37273 10512 37278 10568
rect 37334 10512 37830 10568
rect 37886 10512 37891 10568
rect 37273 10510 37891 10512
rect 37273 10507 37339 10510
rect 37825 10507 37891 10510
rect 37365 10434 37431 10437
rect 37733 10434 37799 10437
rect 37365 10432 37799 10434
rect 0 10298 800 10388
rect 37365 10376 37370 10432
rect 37426 10376 37738 10432
rect 37794 10376 37799 10432
rect 37365 10374 37799 10376
rect 37365 10371 37431 10374
rect 37733 10371 37799 10374
rect 6420 10368 6736 10369
rect 6420 10304 6426 10368
rect 6490 10304 6506 10368
rect 6570 10304 6586 10368
rect 6650 10304 6666 10368
rect 6730 10304 6736 10368
rect 6420 10303 6736 10304
rect 17368 10368 17684 10369
rect 17368 10304 17374 10368
rect 17438 10304 17454 10368
rect 17518 10304 17534 10368
rect 17598 10304 17614 10368
rect 17678 10304 17684 10368
rect 17368 10303 17684 10304
rect 28316 10368 28632 10369
rect 28316 10304 28322 10368
rect 28386 10304 28402 10368
rect 28466 10304 28482 10368
rect 28546 10304 28562 10368
rect 28626 10304 28632 10368
rect 28316 10303 28632 10304
rect 39264 10368 39580 10369
rect 39264 10304 39270 10368
rect 39334 10304 39350 10368
rect 39414 10304 39430 10368
rect 39494 10304 39510 10368
rect 39574 10304 39580 10368
rect 39264 10303 39580 10304
rect 1577 10298 1643 10301
rect 0 10296 1643 10298
rect 0 10240 1582 10296
rect 1638 10240 1643 10296
rect 0 10238 1643 10240
rect 0 10148 800 10238
rect 1577 10235 1643 10238
rect 40309 10162 40375 10165
rect 41321 10162 41387 10165
rect 40309 10160 41387 10162
rect 40309 10104 40314 10160
rect 40370 10104 41326 10160
rect 41382 10104 41387 10160
rect 40309 10102 41387 10104
rect 40309 10099 40375 10102
rect 41321 10099 41387 10102
rect 14273 10026 14339 10029
rect 18689 10026 18755 10029
rect 14273 10024 18755 10026
rect 14273 9968 14278 10024
rect 14334 9968 18694 10024
rect 18750 9968 18755 10024
rect 14273 9966 18755 9968
rect 14273 9963 14339 9966
rect 18689 9963 18755 9966
rect 40309 10026 40375 10029
rect 41137 10026 41203 10029
rect 40309 10024 41203 10026
rect 40309 9968 40314 10024
rect 40370 9968 41142 10024
rect 41198 9968 41203 10024
rect 40309 9966 41203 9968
rect 40309 9963 40375 9966
rect 41137 9963 41203 9966
rect 40677 9890 40743 9893
rect 41689 9890 41755 9893
rect 40677 9888 41755 9890
rect 40677 9832 40682 9888
rect 40738 9832 41694 9888
rect 41750 9832 41755 9888
rect 40677 9830 41755 9832
rect 40677 9827 40743 9830
rect 41689 9827 41755 9830
rect 11894 9824 12210 9825
rect 11894 9760 11900 9824
rect 11964 9760 11980 9824
rect 12044 9760 12060 9824
rect 12124 9760 12140 9824
rect 12204 9760 12210 9824
rect 11894 9759 12210 9760
rect 22842 9824 23158 9825
rect 22842 9760 22848 9824
rect 22912 9760 22928 9824
rect 22992 9760 23008 9824
rect 23072 9760 23088 9824
rect 23152 9760 23158 9824
rect 22842 9759 23158 9760
rect 33790 9824 34106 9825
rect 33790 9760 33796 9824
rect 33860 9760 33876 9824
rect 33940 9760 33956 9824
rect 34020 9760 34036 9824
rect 34100 9760 34106 9824
rect 33790 9759 34106 9760
rect 44738 9824 45054 9825
rect 44738 9760 44744 9824
rect 44808 9760 44824 9824
rect 44888 9760 44904 9824
rect 44968 9760 44984 9824
rect 45048 9760 45054 9824
rect 44738 9759 45054 9760
rect 39665 9618 39731 9621
rect 40953 9618 41019 9621
rect 39665 9616 41019 9618
rect 39665 9560 39670 9616
rect 39726 9560 40958 9616
rect 41014 9560 41019 9616
rect 39665 9558 41019 9560
rect 39665 9555 39731 9558
rect 40953 9555 41019 9558
rect 6420 9280 6736 9281
rect 6420 9216 6426 9280
rect 6490 9216 6506 9280
rect 6570 9216 6586 9280
rect 6650 9216 6666 9280
rect 6730 9216 6736 9280
rect 6420 9215 6736 9216
rect 17368 9280 17684 9281
rect 17368 9216 17374 9280
rect 17438 9216 17454 9280
rect 17518 9216 17534 9280
rect 17598 9216 17614 9280
rect 17678 9216 17684 9280
rect 17368 9215 17684 9216
rect 28316 9280 28632 9281
rect 28316 9216 28322 9280
rect 28386 9216 28402 9280
rect 28466 9216 28482 9280
rect 28546 9216 28562 9280
rect 28626 9216 28632 9280
rect 28316 9215 28632 9216
rect 39264 9280 39580 9281
rect 39264 9216 39270 9280
rect 39334 9216 39350 9280
rect 39414 9216 39430 9280
rect 39494 9216 39510 9280
rect 39574 9216 39580 9280
rect 39264 9215 39580 9216
rect 39205 9074 39271 9077
rect 40217 9074 40283 9077
rect 39205 9072 40283 9074
rect 39205 9016 39210 9072
rect 39266 9016 40222 9072
rect 40278 9016 40283 9072
rect 39205 9014 40283 9016
rect 39205 9011 39271 9014
rect 40217 9011 40283 9014
rect 44173 8938 44239 8941
rect 45200 8938 46000 9028
rect 44173 8936 46000 8938
rect 44173 8880 44178 8936
rect 44234 8880 46000 8936
rect 44173 8878 46000 8880
rect 44173 8875 44239 8878
rect 45200 8788 46000 8878
rect 11894 8736 12210 8737
rect 11894 8672 11900 8736
rect 11964 8672 11980 8736
rect 12044 8672 12060 8736
rect 12124 8672 12140 8736
rect 12204 8672 12210 8736
rect 11894 8671 12210 8672
rect 22842 8736 23158 8737
rect 22842 8672 22848 8736
rect 22912 8672 22928 8736
rect 22992 8672 23008 8736
rect 23072 8672 23088 8736
rect 23152 8672 23158 8736
rect 22842 8671 23158 8672
rect 33790 8736 34106 8737
rect 33790 8672 33796 8736
rect 33860 8672 33876 8736
rect 33940 8672 33956 8736
rect 34020 8672 34036 8736
rect 34100 8672 34106 8736
rect 33790 8671 34106 8672
rect 44738 8736 45054 8737
rect 44738 8672 44744 8736
rect 44808 8672 44824 8736
rect 44888 8672 44904 8736
rect 44968 8672 44984 8736
rect 45048 8672 45054 8736
rect 44738 8671 45054 8672
rect 32397 8530 32463 8533
rect 36169 8530 36235 8533
rect 32397 8528 36235 8530
rect 32397 8472 32402 8528
rect 32458 8472 36174 8528
rect 36230 8472 36235 8528
rect 32397 8470 36235 8472
rect 32397 8467 32463 8470
rect 36169 8467 36235 8470
rect 0 8258 800 8348
rect 1577 8258 1643 8261
rect 0 8256 1643 8258
rect 0 8200 1582 8256
rect 1638 8200 1643 8256
rect 0 8198 1643 8200
rect 0 8108 800 8198
rect 1577 8195 1643 8198
rect 6420 8192 6736 8193
rect 6420 8128 6426 8192
rect 6490 8128 6506 8192
rect 6570 8128 6586 8192
rect 6650 8128 6666 8192
rect 6730 8128 6736 8192
rect 6420 8127 6736 8128
rect 17368 8192 17684 8193
rect 17368 8128 17374 8192
rect 17438 8128 17454 8192
rect 17518 8128 17534 8192
rect 17598 8128 17614 8192
rect 17678 8128 17684 8192
rect 17368 8127 17684 8128
rect 28316 8192 28632 8193
rect 28316 8128 28322 8192
rect 28386 8128 28402 8192
rect 28466 8128 28482 8192
rect 28546 8128 28562 8192
rect 28626 8128 28632 8192
rect 28316 8127 28632 8128
rect 39264 8192 39580 8193
rect 39264 8128 39270 8192
rect 39334 8128 39350 8192
rect 39414 8128 39430 8192
rect 39494 8128 39510 8192
rect 39574 8128 39580 8192
rect 39264 8127 39580 8128
rect 20437 7850 20503 7853
rect 26049 7850 26115 7853
rect 20437 7848 26115 7850
rect 20437 7792 20442 7848
rect 20498 7792 26054 7848
rect 26110 7792 26115 7848
rect 20437 7790 26115 7792
rect 20437 7787 20503 7790
rect 26049 7787 26115 7790
rect 44173 7850 44239 7853
rect 44173 7848 45202 7850
rect 44173 7792 44178 7848
rect 44234 7792 45202 7848
rect 44173 7790 45202 7792
rect 44173 7787 44239 7790
rect 45142 7668 45202 7790
rect 11894 7648 12210 7649
rect 11894 7584 11900 7648
rect 11964 7584 11980 7648
rect 12044 7584 12060 7648
rect 12124 7584 12140 7648
rect 12204 7584 12210 7648
rect 11894 7583 12210 7584
rect 22842 7648 23158 7649
rect 22842 7584 22848 7648
rect 22912 7584 22928 7648
rect 22992 7584 23008 7648
rect 23072 7584 23088 7648
rect 23152 7584 23158 7648
rect 22842 7583 23158 7584
rect 33790 7648 34106 7649
rect 33790 7584 33796 7648
rect 33860 7584 33876 7648
rect 33940 7584 33956 7648
rect 34020 7584 34036 7648
rect 34100 7584 34106 7648
rect 33790 7583 34106 7584
rect 44738 7648 45054 7649
rect 44738 7584 44744 7648
rect 44808 7584 44824 7648
rect 44888 7584 44904 7648
rect 44968 7584 44984 7648
rect 45048 7584 45054 7648
rect 44738 7583 45054 7584
rect 45142 7518 46000 7668
rect 22369 7442 22435 7445
rect 27705 7442 27771 7445
rect 22369 7440 27771 7442
rect 22369 7384 22374 7440
rect 22430 7384 27710 7440
rect 27766 7384 27771 7440
rect 45200 7428 46000 7518
rect 22369 7382 27771 7384
rect 22369 7379 22435 7382
rect 27705 7379 27771 7382
rect 6420 7104 6736 7105
rect 6420 7040 6426 7104
rect 6490 7040 6506 7104
rect 6570 7040 6586 7104
rect 6650 7040 6666 7104
rect 6730 7040 6736 7104
rect 6420 7039 6736 7040
rect 17368 7104 17684 7105
rect 17368 7040 17374 7104
rect 17438 7040 17454 7104
rect 17518 7040 17534 7104
rect 17598 7040 17614 7104
rect 17678 7040 17684 7104
rect 17368 7039 17684 7040
rect 28316 7104 28632 7105
rect 28316 7040 28322 7104
rect 28386 7040 28402 7104
rect 28466 7040 28482 7104
rect 28546 7040 28562 7104
rect 28626 7040 28632 7104
rect 28316 7039 28632 7040
rect 39264 7104 39580 7105
rect 39264 7040 39270 7104
rect 39334 7040 39350 7104
rect 39414 7040 39430 7104
rect 39494 7040 39510 7104
rect 39574 7040 39580 7104
rect 39264 7039 39580 7040
rect 0 6898 800 6988
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6748 800 6838
rect 1577 6835 1643 6838
rect 27429 6898 27495 6901
rect 33133 6898 33199 6901
rect 27429 6896 33199 6898
rect 27429 6840 27434 6896
rect 27490 6840 33138 6896
rect 33194 6840 33199 6896
rect 27429 6838 33199 6840
rect 27429 6835 27495 6838
rect 33133 6835 33199 6838
rect 11894 6560 12210 6561
rect 11894 6496 11900 6560
rect 11964 6496 11980 6560
rect 12044 6496 12060 6560
rect 12124 6496 12140 6560
rect 12204 6496 12210 6560
rect 11894 6495 12210 6496
rect 22842 6560 23158 6561
rect 22842 6496 22848 6560
rect 22912 6496 22928 6560
rect 22992 6496 23008 6560
rect 23072 6496 23088 6560
rect 23152 6496 23158 6560
rect 22842 6495 23158 6496
rect 33790 6560 34106 6561
rect 33790 6496 33796 6560
rect 33860 6496 33876 6560
rect 33940 6496 33956 6560
rect 34020 6496 34036 6560
rect 34100 6496 34106 6560
rect 33790 6495 34106 6496
rect 44738 6560 45054 6561
rect 44738 6496 44744 6560
rect 44808 6496 44824 6560
rect 44888 6496 44904 6560
rect 44968 6496 44984 6560
rect 45048 6496 45054 6560
rect 44738 6495 45054 6496
rect 6420 6016 6736 6017
rect 6420 5952 6426 6016
rect 6490 5952 6506 6016
rect 6570 5952 6586 6016
rect 6650 5952 6666 6016
rect 6730 5952 6736 6016
rect 6420 5951 6736 5952
rect 17368 6016 17684 6017
rect 17368 5952 17374 6016
rect 17438 5952 17454 6016
rect 17518 5952 17534 6016
rect 17598 5952 17614 6016
rect 17678 5952 17684 6016
rect 17368 5951 17684 5952
rect 28316 6016 28632 6017
rect 28316 5952 28322 6016
rect 28386 5952 28402 6016
rect 28466 5952 28482 6016
rect 28546 5952 28562 6016
rect 28626 5952 28632 6016
rect 28316 5951 28632 5952
rect 39264 6016 39580 6017
rect 39264 5952 39270 6016
rect 39334 5952 39350 6016
rect 39414 5952 39430 6016
rect 39494 5952 39510 6016
rect 39574 5952 39580 6016
rect 39264 5951 39580 5952
rect 8201 5674 8267 5677
rect 12709 5674 12775 5677
rect 8201 5672 12775 5674
rect 8201 5616 8206 5672
rect 8262 5616 12714 5672
rect 12770 5616 12775 5672
rect 8201 5614 12775 5616
rect 8201 5611 8267 5614
rect 12709 5611 12775 5614
rect 20621 5674 20687 5677
rect 26417 5674 26483 5677
rect 20621 5672 26483 5674
rect 20621 5616 20626 5672
rect 20682 5616 26422 5672
rect 26478 5616 26483 5672
rect 20621 5614 26483 5616
rect 20621 5611 20687 5614
rect 26417 5611 26483 5614
rect 27797 5674 27863 5677
rect 28625 5674 28691 5677
rect 27797 5672 28691 5674
rect 27797 5616 27802 5672
rect 27858 5616 28630 5672
rect 28686 5616 28691 5672
rect 27797 5614 28691 5616
rect 27797 5611 27863 5614
rect 28625 5611 28691 5614
rect 45200 5538 46000 5628
rect 11894 5472 12210 5473
rect 11894 5408 11900 5472
rect 11964 5408 11980 5472
rect 12044 5408 12060 5472
rect 12124 5408 12140 5472
rect 12204 5408 12210 5472
rect 11894 5407 12210 5408
rect 22842 5472 23158 5473
rect 22842 5408 22848 5472
rect 22912 5408 22928 5472
rect 22992 5408 23008 5472
rect 23072 5408 23088 5472
rect 23152 5408 23158 5472
rect 22842 5407 23158 5408
rect 33790 5472 34106 5473
rect 33790 5408 33796 5472
rect 33860 5408 33876 5472
rect 33940 5408 33956 5472
rect 34020 5408 34036 5472
rect 34100 5408 34106 5472
rect 33790 5407 34106 5408
rect 44738 5472 45054 5473
rect 44738 5408 44744 5472
rect 44808 5408 44824 5472
rect 44888 5408 44904 5472
rect 44968 5408 44984 5472
rect 45048 5408 45054 5472
rect 44738 5407 45054 5408
rect 45142 5388 46000 5538
rect 44081 5266 44147 5269
rect 45142 5266 45202 5388
rect 44081 5264 45202 5266
rect 44081 5208 44086 5264
rect 44142 5208 45202 5264
rect 44081 5206 45202 5208
rect 44081 5203 44147 5206
rect 0 4858 800 4948
rect 6420 4928 6736 4929
rect 6420 4864 6426 4928
rect 6490 4864 6506 4928
rect 6570 4864 6586 4928
rect 6650 4864 6666 4928
rect 6730 4864 6736 4928
rect 6420 4863 6736 4864
rect 17368 4928 17684 4929
rect 17368 4864 17374 4928
rect 17438 4864 17454 4928
rect 17518 4864 17534 4928
rect 17598 4864 17614 4928
rect 17678 4864 17684 4928
rect 17368 4863 17684 4864
rect 28316 4928 28632 4929
rect 28316 4864 28322 4928
rect 28386 4864 28402 4928
rect 28466 4864 28482 4928
rect 28546 4864 28562 4928
rect 28626 4864 28632 4928
rect 28316 4863 28632 4864
rect 39264 4928 39580 4929
rect 39264 4864 39270 4928
rect 39334 4864 39350 4928
rect 39414 4864 39430 4928
rect 39494 4864 39510 4928
rect 39574 4864 39580 4928
rect 39264 4863 39580 4864
rect 1393 4858 1459 4861
rect 0 4856 1459 4858
rect 0 4800 1398 4856
rect 1454 4800 1459 4856
rect 0 4798 1459 4800
rect 0 4708 800 4798
rect 1393 4795 1459 4798
rect 11894 4384 12210 4385
rect 11894 4320 11900 4384
rect 11964 4320 11980 4384
rect 12044 4320 12060 4384
rect 12124 4320 12140 4384
rect 12204 4320 12210 4384
rect 11894 4319 12210 4320
rect 22842 4384 23158 4385
rect 22842 4320 22848 4384
rect 22912 4320 22928 4384
rect 22992 4320 23008 4384
rect 23072 4320 23088 4384
rect 23152 4320 23158 4384
rect 22842 4319 23158 4320
rect 33790 4384 34106 4385
rect 33790 4320 33796 4384
rect 33860 4320 33876 4384
rect 33940 4320 33956 4384
rect 34020 4320 34036 4384
rect 34100 4320 34106 4384
rect 33790 4319 34106 4320
rect 44738 4384 45054 4385
rect 44738 4320 44744 4384
rect 44808 4320 44824 4384
rect 44888 4320 44904 4384
rect 44968 4320 44984 4384
rect 45048 4320 45054 4384
rect 44738 4319 45054 4320
rect 44081 4178 44147 4181
rect 45200 4178 46000 4268
rect 44081 4176 46000 4178
rect 44081 4120 44086 4176
rect 44142 4120 46000 4176
rect 44081 4118 46000 4120
rect 44081 4115 44147 4118
rect 45200 4028 46000 4118
rect 6420 3840 6736 3841
rect 6420 3776 6426 3840
rect 6490 3776 6506 3840
rect 6570 3776 6586 3840
rect 6650 3776 6666 3840
rect 6730 3776 6736 3840
rect 6420 3775 6736 3776
rect 17368 3840 17684 3841
rect 17368 3776 17374 3840
rect 17438 3776 17454 3840
rect 17518 3776 17534 3840
rect 17598 3776 17614 3840
rect 17678 3776 17684 3840
rect 17368 3775 17684 3776
rect 28316 3840 28632 3841
rect 28316 3776 28322 3840
rect 28386 3776 28402 3840
rect 28466 3776 28482 3840
rect 28546 3776 28562 3840
rect 28626 3776 28632 3840
rect 28316 3775 28632 3776
rect 39264 3840 39580 3841
rect 39264 3776 39270 3840
rect 39334 3776 39350 3840
rect 39414 3776 39430 3840
rect 39494 3776 39510 3840
rect 39574 3776 39580 3840
rect 39264 3775 39580 3776
rect 0 3498 800 3588
rect 1577 3498 1643 3501
rect 0 3496 1643 3498
rect 0 3440 1582 3496
rect 1638 3440 1643 3496
rect 0 3438 1643 3440
rect 0 3348 800 3438
rect 1577 3435 1643 3438
rect 11894 3296 12210 3297
rect 11894 3232 11900 3296
rect 11964 3232 11980 3296
rect 12044 3232 12060 3296
rect 12124 3232 12140 3296
rect 12204 3232 12210 3296
rect 11894 3231 12210 3232
rect 22842 3296 23158 3297
rect 22842 3232 22848 3296
rect 22912 3232 22928 3296
rect 22992 3232 23008 3296
rect 23072 3232 23088 3296
rect 23152 3232 23158 3296
rect 22842 3231 23158 3232
rect 33790 3296 34106 3297
rect 33790 3232 33796 3296
rect 33860 3232 33876 3296
rect 33940 3232 33956 3296
rect 34020 3232 34036 3296
rect 34100 3232 34106 3296
rect 33790 3231 34106 3232
rect 44738 3296 45054 3297
rect 44738 3232 44744 3296
rect 44808 3232 44824 3296
rect 44888 3232 44904 3296
rect 44968 3232 44984 3296
rect 45048 3232 45054 3296
rect 44738 3231 45054 3232
rect 6420 2752 6736 2753
rect 6420 2688 6426 2752
rect 6490 2688 6506 2752
rect 6570 2688 6586 2752
rect 6650 2688 6666 2752
rect 6730 2688 6736 2752
rect 6420 2687 6736 2688
rect 17368 2752 17684 2753
rect 17368 2688 17374 2752
rect 17438 2688 17454 2752
rect 17518 2688 17534 2752
rect 17598 2688 17614 2752
rect 17678 2688 17684 2752
rect 17368 2687 17684 2688
rect 28316 2752 28632 2753
rect 28316 2688 28322 2752
rect 28386 2688 28402 2752
rect 28466 2688 28482 2752
rect 28546 2688 28562 2752
rect 28626 2688 28632 2752
rect 28316 2687 28632 2688
rect 39264 2752 39580 2753
rect 39264 2688 39270 2752
rect 39334 2688 39350 2752
rect 39414 2688 39430 2752
rect 39494 2688 39510 2752
rect 39574 2688 39580 2752
rect 39264 2687 39580 2688
rect 44081 2410 44147 2413
rect 44081 2408 45202 2410
rect 44081 2352 44086 2408
rect 44142 2352 45202 2408
rect 44081 2350 45202 2352
rect 44081 2347 44147 2350
rect 45142 2228 45202 2350
rect 11894 2208 12210 2209
rect 11894 2144 11900 2208
rect 11964 2144 11980 2208
rect 12044 2144 12060 2208
rect 12124 2144 12140 2208
rect 12204 2144 12210 2208
rect 11894 2143 12210 2144
rect 22842 2208 23158 2209
rect 22842 2144 22848 2208
rect 22912 2144 22928 2208
rect 22992 2144 23008 2208
rect 23072 2144 23088 2208
rect 23152 2144 23158 2208
rect 22842 2143 23158 2144
rect 33790 2208 34106 2209
rect 33790 2144 33796 2208
rect 33860 2144 33876 2208
rect 33940 2144 33956 2208
rect 34020 2144 34036 2208
rect 34100 2144 34106 2208
rect 33790 2143 34106 2144
rect 44738 2208 45054 2209
rect 44738 2144 44744 2208
rect 44808 2144 44824 2208
rect 44888 2144 44904 2208
rect 44968 2144 44984 2208
rect 45048 2144 45054 2208
rect 44738 2143 45054 2144
rect 45142 2078 46000 2228
rect 45200 1988 46000 2078
rect 0 1458 800 1548
rect 1577 1458 1643 1461
rect 0 1456 1643 1458
rect 0 1400 1582 1456
rect 1638 1400 1643 1456
rect 0 1398 1643 1400
rect 0 1308 800 1398
rect 1577 1395 1643 1398
rect 44173 778 44239 781
rect 45200 778 46000 868
rect 44173 776 46000 778
rect 44173 720 44178 776
rect 44234 720 46000 776
rect 44173 718 46000 720
rect 44173 715 44239 718
rect 45200 628 46000 718
<< via3 >>
rect 11900 17436 11964 17440
rect 11900 17380 11904 17436
rect 11904 17380 11960 17436
rect 11960 17380 11964 17436
rect 11900 17376 11964 17380
rect 11980 17436 12044 17440
rect 11980 17380 11984 17436
rect 11984 17380 12040 17436
rect 12040 17380 12044 17436
rect 11980 17376 12044 17380
rect 12060 17436 12124 17440
rect 12060 17380 12064 17436
rect 12064 17380 12120 17436
rect 12120 17380 12124 17436
rect 12060 17376 12124 17380
rect 12140 17436 12204 17440
rect 12140 17380 12144 17436
rect 12144 17380 12200 17436
rect 12200 17380 12204 17436
rect 12140 17376 12204 17380
rect 22848 17436 22912 17440
rect 22848 17380 22852 17436
rect 22852 17380 22908 17436
rect 22908 17380 22912 17436
rect 22848 17376 22912 17380
rect 22928 17436 22992 17440
rect 22928 17380 22932 17436
rect 22932 17380 22988 17436
rect 22988 17380 22992 17436
rect 22928 17376 22992 17380
rect 23008 17436 23072 17440
rect 23008 17380 23012 17436
rect 23012 17380 23068 17436
rect 23068 17380 23072 17436
rect 23008 17376 23072 17380
rect 23088 17436 23152 17440
rect 23088 17380 23092 17436
rect 23092 17380 23148 17436
rect 23148 17380 23152 17436
rect 23088 17376 23152 17380
rect 33796 17436 33860 17440
rect 33796 17380 33800 17436
rect 33800 17380 33856 17436
rect 33856 17380 33860 17436
rect 33796 17376 33860 17380
rect 33876 17436 33940 17440
rect 33876 17380 33880 17436
rect 33880 17380 33936 17436
rect 33936 17380 33940 17436
rect 33876 17376 33940 17380
rect 33956 17436 34020 17440
rect 33956 17380 33960 17436
rect 33960 17380 34016 17436
rect 34016 17380 34020 17436
rect 33956 17376 34020 17380
rect 34036 17436 34100 17440
rect 34036 17380 34040 17436
rect 34040 17380 34096 17436
rect 34096 17380 34100 17436
rect 34036 17376 34100 17380
rect 44744 17436 44808 17440
rect 44744 17380 44748 17436
rect 44748 17380 44804 17436
rect 44804 17380 44808 17436
rect 44744 17376 44808 17380
rect 44824 17436 44888 17440
rect 44824 17380 44828 17436
rect 44828 17380 44884 17436
rect 44884 17380 44888 17436
rect 44824 17376 44888 17380
rect 44904 17436 44968 17440
rect 44904 17380 44908 17436
rect 44908 17380 44964 17436
rect 44964 17380 44968 17436
rect 44904 17376 44968 17380
rect 44984 17436 45048 17440
rect 44984 17380 44988 17436
rect 44988 17380 45044 17436
rect 45044 17380 45048 17436
rect 44984 17376 45048 17380
rect 6426 16892 6490 16896
rect 6426 16836 6430 16892
rect 6430 16836 6486 16892
rect 6486 16836 6490 16892
rect 6426 16832 6490 16836
rect 6506 16892 6570 16896
rect 6506 16836 6510 16892
rect 6510 16836 6566 16892
rect 6566 16836 6570 16892
rect 6506 16832 6570 16836
rect 6586 16892 6650 16896
rect 6586 16836 6590 16892
rect 6590 16836 6646 16892
rect 6646 16836 6650 16892
rect 6586 16832 6650 16836
rect 6666 16892 6730 16896
rect 6666 16836 6670 16892
rect 6670 16836 6726 16892
rect 6726 16836 6730 16892
rect 6666 16832 6730 16836
rect 17374 16892 17438 16896
rect 17374 16836 17378 16892
rect 17378 16836 17434 16892
rect 17434 16836 17438 16892
rect 17374 16832 17438 16836
rect 17454 16892 17518 16896
rect 17454 16836 17458 16892
rect 17458 16836 17514 16892
rect 17514 16836 17518 16892
rect 17454 16832 17518 16836
rect 17534 16892 17598 16896
rect 17534 16836 17538 16892
rect 17538 16836 17594 16892
rect 17594 16836 17598 16892
rect 17534 16832 17598 16836
rect 17614 16892 17678 16896
rect 17614 16836 17618 16892
rect 17618 16836 17674 16892
rect 17674 16836 17678 16892
rect 17614 16832 17678 16836
rect 28322 16892 28386 16896
rect 28322 16836 28326 16892
rect 28326 16836 28382 16892
rect 28382 16836 28386 16892
rect 28322 16832 28386 16836
rect 28402 16892 28466 16896
rect 28402 16836 28406 16892
rect 28406 16836 28462 16892
rect 28462 16836 28466 16892
rect 28402 16832 28466 16836
rect 28482 16892 28546 16896
rect 28482 16836 28486 16892
rect 28486 16836 28542 16892
rect 28542 16836 28546 16892
rect 28482 16832 28546 16836
rect 28562 16892 28626 16896
rect 28562 16836 28566 16892
rect 28566 16836 28622 16892
rect 28622 16836 28626 16892
rect 28562 16832 28626 16836
rect 39270 16892 39334 16896
rect 39270 16836 39274 16892
rect 39274 16836 39330 16892
rect 39330 16836 39334 16892
rect 39270 16832 39334 16836
rect 39350 16892 39414 16896
rect 39350 16836 39354 16892
rect 39354 16836 39410 16892
rect 39410 16836 39414 16892
rect 39350 16832 39414 16836
rect 39430 16892 39494 16896
rect 39430 16836 39434 16892
rect 39434 16836 39490 16892
rect 39490 16836 39494 16892
rect 39430 16832 39494 16836
rect 39510 16892 39574 16896
rect 39510 16836 39514 16892
rect 39514 16836 39570 16892
rect 39570 16836 39574 16892
rect 39510 16832 39574 16836
rect 11900 16348 11964 16352
rect 11900 16292 11904 16348
rect 11904 16292 11960 16348
rect 11960 16292 11964 16348
rect 11900 16288 11964 16292
rect 11980 16348 12044 16352
rect 11980 16292 11984 16348
rect 11984 16292 12040 16348
rect 12040 16292 12044 16348
rect 11980 16288 12044 16292
rect 12060 16348 12124 16352
rect 12060 16292 12064 16348
rect 12064 16292 12120 16348
rect 12120 16292 12124 16348
rect 12060 16288 12124 16292
rect 12140 16348 12204 16352
rect 12140 16292 12144 16348
rect 12144 16292 12200 16348
rect 12200 16292 12204 16348
rect 12140 16288 12204 16292
rect 22848 16348 22912 16352
rect 22848 16292 22852 16348
rect 22852 16292 22908 16348
rect 22908 16292 22912 16348
rect 22848 16288 22912 16292
rect 22928 16348 22992 16352
rect 22928 16292 22932 16348
rect 22932 16292 22988 16348
rect 22988 16292 22992 16348
rect 22928 16288 22992 16292
rect 23008 16348 23072 16352
rect 23008 16292 23012 16348
rect 23012 16292 23068 16348
rect 23068 16292 23072 16348
rect 23008 16288 23072 16292
rect 23088 16348 23152 16352
rect 23088 16292 23092 16348
rect 23092 16292 23148 16348
rect 23148 16292 23152 16348
rect 23088 16288 23152 16292
rect 33796 16348 33860 16352
rect 33796 16292 33800 16348
rect 33800 16292 33856 16348
rect 33856 16292 33860 16348
rect 33796 16288 33860 16292
rect 33876 16348 33940 16352
rect 33876 16292 33880 16348
rect 33880 16292 33936 16348
rect 33936 16292 33940 16348
rect 33876 16288 33940 16292
rect 33956 16348 34020 16352
rect 33956 16292 33960 16348
rect 33960 16292 34016 16348
rect 34016 16292 34020 16348
rect 33956 16288 34020 16292
rect 34036 16348 34100 16352
rect 34036 16292 34040 16348
rect 34040 16292 34096 16348
rect 34096 16292 34100 16348
rect 34036 16288 34100 16292
rect 44744 16348 44808 16352
rect 44744 16292 44748 16348
rect 44748 16292 44804 16348
rect 44804 16292 44808 16348
rect 44744 16288 44808 16292
rect 44824 16348 44888 16352
rect 44824 16292 44828 16348
rect 44828 16292 44884 16348
rect 44884 16292 44888 16348
rect 44824 16288 44888 16292
rect 44904 16348 44968 16352
rect 44904 16292 44908 16348
rect 44908 16292 44964 16348
rect 44964 16292 44968 16348
rect 44904 16288 44968 16292
rect 44984 16348 45048 16352
rect 44984 16292 44988 16348
rect 44988 16292 45044 16348
rect 45044 16292 45048 16348
rect 44984 16288 45048 16292
rect 6426 15804 6490 15808
rect 6426 15748 6430 15804
rect 6430 15748 6486 15804
rect 6486 15748 6490 15804
rect 6426 15744 6490 15748
rect 6506 15804 6570 15808
rect 6506 15748 6510 15804
rect 6510 15748 6566 15804
rect 6566 15748 6570 15804
rect 6506 15744 6570 15748
rect 6586 15804 6650 15808
rect 6586 15748 6590 15804
rect 6590 15748 6646 15804
rect 6646 15748 6650 15804
rect 6586 15744 6650 15748
rect 6666 15804 6730 15808
rect 6666 15748 6670 15804
rect 6670 15748 6726 15804
rect 6726 15748 6730 15804
rect 6666 15744 6730 15748
rect 17374 15804 17438 15808
rect 17374 15748 17378 15804
rect 17378 15748 17434 15804
rect 17434 15748 17438 15804
rect 17374 15744 17438 15748
rect 17454 15804 17518 15808
rect 17454 15748 17458 15804
rect 17458 15748 17514 15804
rect 17514 15748 17518 15804
rect 17454 15744 17518 15748
rect 17534 15804 17598 15808
rect 17534 15748 17538 15804
rect 17538 15748 17594 15804
rect 17594 15748 17598 15804
rect 17534 15744 17598 15748
rect 17614 15804 17678 15808
rect 17614 15748 17618 15804
rect 17618 15748 17674 15804
rect 17674 15748 17678 15804
rect 17614 15744 17678 15748
rect 28322 15804 28386 15808
rect 28322 15748 28326 15804
rect 28326 15748 28382 15804
rect 28382 15748 28386 15804
rect 28322 15744 28386 15748
rect 28402 15804 28466 15808
rect 28402 15748 28406 15804
rect 28406 15748 28462 15804
rect 28462 15748 28466 15804
rect 28402 15744 28466 15748
rect 28482 15804 28546 15808
rect 28482 15748 28486 15804
rect 28486 15748 28542 15804
rect 28542 15748 28546 15804
rect 28482 15744 28546 15748
rect 28562 15804 28626 15808
rect 28562 15748 28566 15804
rect 28566 15748 28622 15804
rect 28622 15748 28626 15804
rect 28562 15744 28626 15748
rect 39270 15804 39334 15808
rect 39270 15748 39274 15804
rect 39274 15748 39330 15804
rect 39330 15748 39334 15804
rect 39270 15744 39334 15748
rect 39350 15804 39414 15808
rect 39350 15748 39354 15804
rect 39354 15748 39410 15804
rect 39410 15748 39414 15804
rect 39350 15744 39414 15748
rect 39430 15804 39494 15808
rect 39430 15748 39434 15804
rect 39434 15748 39490 15804
rect 39490 15748 39494 15804
rect 39430 15744 39494 15748
rect 39510 15804 39574 15808
rect 39510 15748 39514 15804
rect 39514 15748 39570 15804
rect 39570 15748 39574 15804
rect 39510 15744 39574 15748
rect 11900 15260 11964 15264
rect 11900 15204 11904 15260
rect 11904 15204 11960 15260
rect 11960 15204 11964 15260
rect 11900 15200 11964 15204
rect 11980 15260 12044 15264
rect 11980 15204 11984 15260
rect 11984 15204 12040 15260
rect 12040 15204 12044 15260
rect 11980 15200 12044 15204
rect 12060 15260 12124 15264
rect 12060 15204 12064 15260
rect 12064 15204 12120 15260
rect 12120 15204 12124 15260
rect 12060 15200 12124 15204
rect 12140 15260 12204 15264
rect 12140 15204 12144 15260
rect 12144 15204 12200 15260
rect 12200 15204 12204 15260
rect 12140 15200 12204 15204
rect 22848 15260 22912 15264
rect 22848 15204 22852 15260
rect 22852 15204 22908 15260
rect 22908 15204 22912 15260
rect 22848 15200 22912 15204
rect 22928 15260 22992 15264
rect 22928 15204 22932 15260
rect 22932 15204 22988 15260
rect 22988 15204 22992 15260
rect 22928 15200 22992 15204
rect 23008 15260 23072 15264
rect 23008 15204 23012 15260
rect 23012 15204 23068 15260
rect 23068 15204 23072 15260
rect 23008 15200 23072 15204
rect 23088 15260 23152 15264
rect 23088 15204 23092 15260
rect 23092 15204 23148 15260
rect 23148 15204 23152 15260
rect 23088 15200 23152 15204
rect 33796 15260 33860 15264
rect 33796 15204 33800 15260
rect 33800 15204 33856 15260
rect 33856 15204 33860 15260
rect 33796 15200 33860 15204
rect 33876 15260 33940 15264
rect 33876 15204 33880 15260
rect 33880 15204 33936 15260
rect 33936 15204 33940 15260
rect 33876 15200 33940 15204
rect 33956 15260 34020 15264
rect 33956 15204 33960 15260
rect 33960 15204 34016 15260
rect 34016 15204 34020 15260
rect 33956 15200 34020 15204
rect 34036 15260 34100 15264
rect 34036 15204 34040 15260
rect 34040 15204 34096 15260
rect 34096 15204 34100 15260
rect 34036 15200 34100 15204
rect 44744 15260 44808 15264
rect 44744 15204 44748 15260
rect 44748 15204 44804 15260
rect 44804 15204 44808 15260
rect 44744 15200 44808 15204
rect 44824 15260 44888 15264
rect 44824 15204 44828 15260
rect 44828 15204 44884 15260
rect 44884 15204 44888 15260
rect 44824 15200 44888 15204
rect 44904 15260 44968 15264
rect 44904 15204 44908 15260
rect 44908 15204 44964 15260
rect 44964 15204 44968 15260
rect 44904 15200 44968 15204
rect 44984 15260 45048 15264
rect 44984 15204 44988 15260
rect 44988 15204 45044 15260
rect 45044 15204 45048 15260
rect 44984 15200 45048 15204
rect 6426 14716 6490 14720
rect 6426 14660 6430 14716
rect 6430 14660 6486 14716
rect 6486 14660 6490 14716
rect 6426 14656 6490 14660
rect 6506 14716 6570 14720
rect 6506 14660 6510 14716
rect 6510 14660 6566 14716
rect 6566 14660 6570 14716
rect 6506 14656 6570 14660
rect 6586 14716 6650 14720
rect 6586 14660 6590 14716
rect 6590 14660 6646 14716
rect 6646 14660 6650 14716
rect 6586 14656 6650 14660
rect 6666 14716 6730 14720
rect 6666 14660 6670 14716
rect 6670 14660 6726 14716
rect 6726 14660 6730 14716
rect 6666 14656 6730 14660
rect 17374 14716 17438 14720
rect 17374 14660 17378 14716
rect 17378 14660 17434 14716
rect 17434 14660 17438 14716
rect 17374 14656 17438 14660
rect 17454 14716 17518 14720
rect 17454 14660 17458 14716
rect 17458 14660 17514 14716
rect 17514 14660 17518 14716
rect 17454 14656 17518 14660
rect 17534 14716 17598 14720
rect 17534 14660 17538 14716
rect 17538 14660 17594 14716
rect 17594 14660 17598 14716
rect 17534 14656 17598 14660
rect 17614 14716 17678 14720
rect 17614 14660 17618 14716
rect 17618 14660 17674 14716
rect 17674 14660 17678 14716
rect 17614 14656 17678 14660
rect 28322 14716 28386 14720
rect 28322 14660 28326 14716
rect 28326 14660 28382 14716
rect 28382 14660 28386 14716
rect 28322 14656 28386 14660
rect 28402 14716 28466 14720
rect 28402 14660 28406 14716
rect 28406 14660 28462 14716
rect 28462 14660 28466 14716
rect 28402 14656 28466 14660
rect 28482 14716 28546 14720
rect 28482 14660 28486 14716
rect 28486 14660 28542 14716
rect 28542 14660 28546 14716
rect 28482 14656 28546 14660
rect 28562 14716 28626 14720
rect 28562 14660 28566 14716
rect 28566 14660 28622 14716
rect 28622 14660 28626 14716
rect 28562 14656 28626 14660
rect 39270 14716 39334 14720
rect 39270 14660 39274 14716
rect 39274 14660 39330 14716
rect 39330 14660 39334 14716
rect 39270 14656 39334 14660
rect 39350 14716 39414 14720
rect 39350 14660 39354 14716
rect 39354 14660 39410 14716
rect 39410 14660 39414 14716
rect 39350 14656 39414 14660
rect 39430 14716 39494 14720
rect 39430 14660 39434 14716
rect 39434 14660 39490 14716
rect 39490 14660 39494 14716
rect 39430 14656 39494 14660
rect 39510 14716 39574 14720
rect 39510 14660 39514 14716
rect 39514 14660 39570 14716
rect 39570 14660 39574 14716
rect 39510 14656 39574 14660
rect 11900 14172 11964 14176
rect 11900 14116 11904 14172
rect 11904 14116 11960 14172
rect 11960 14116 11964 14172
rect 11900 14112 11964 14116
rect 11980 14172 12044 14176
rect 11980 14116 11984 14172
rect 11984 14116 12040 14172
rect 12040 14116 12044 14172
rect 11980 14112 12044 14116
rect 12060 14172 12124 14176
rect 12060 14116 12064 14172
rect 12064 14116 12120 14172
rect 12120 14116 12124 14172
rect 12060 14112 12124 14116
rect 12140 14172 12204 14176
rect 12140 14116 12144 14172
rect 12144 14116 12200 14172
rect 12200 14116 12204 14172
rect 12140 14112 12204 14116
rect 22848 14172 22912 14176
rect 22848 14116 22852 14172
rect 22852 14116 22908 14172
rect 22908 14116 22912 14172
rect 22848 14112 22912 14116
rect 22928 14172 22992 14176
rect 22928 14116 22932 14172
rect 22932 14116 22988 14172
rect 22988 14116 22992 14172
rect 22928 14112 22992 14116
rect 23008 14172 23072 14176
rect 23008 14116 23012 14172
rect 23012 14116 23068 14172
rect 23068 14116 23072 14172
rect 23008 14112 23072 14116
rect 23088 14172 23152 14176
rect 23088 14116 23092 14172
rect 23092 14116 23148 14172
rect 23148 14116 23152 14172
rect 23088 14112 23152 14116
rect 33796 14172 33860 14176
rect 33796 14116 33800 14172
rect 33800 14116 33856 14172
rect 33856 14116 33860 14172
rect 33796 14112 33860 14116
rect 33876 14172 33940 14176
rect 33876 14116 33880 14172
rect 33880 14116 33936 14172
rect 33936 14116 33940 14172
rect 33876 14112 33940 14116
rect 33956 14172 34020 14176
rect 33956 14116 33960 14172
rect 33960 14116 34016 14172
rect 34016 14116 34020 14172
rect 33956 14112 34020 14116
rect 34036 14172 34100 14176
rect 34036 14116 34040 14172
rect 34040 14116 34096 14172
rect 34096 14116 34100 14172
rect 34036 14112 34100 14116
rect 44744 14172 44808 14176
rect 44744 14116 44748 14172
rect 44748 14116 44804 14172
rect 44804 14116 44808 14172
rect 44744 14112 44808 14116
rect 44824 14172 44888 14176
rect 44824 14116 44828 14172
rect 44828 14116 44884 14172
rect 44884 14116 44888 14172
rect 44824 14112 44888 14116
rect 44904 14172 44968 14176
rect 44904 14116 44908 14172
rect 44908 14116 44964 14172
rect 44964 14116 44968 14172
rect 44904 14112 44968 14116
rect 44984 14172 45048 14176
rect 44984 14116 44988 14172
rect 44988 14116 45044 14172
rect 45044 14116 45048 14172
rect 44984 14112 45048 14116
rect 6426 13628 6490 13632
rect 6426 13572 6430 13628
rect 6430 13572 6486 13628
rect 6486 13572 6490 13628
rect 6426 13568 6490 13572
rect 6506 13628 6570 13632
rect 6506 13572 6510 13628
rect 6510 13572 6566 13628
rect 6566 13572 6570 13628
rect 6506 13568 6570 13572
rect 6586 13628 6650 13632
rect 6586 13572 6590 13628
rect 6590 13572 6646 13628
rect 6646 13572 6650 13628
rect 6586 13568 6650 13572
rect 6666 13628 6730 13632
rect 6666 13572 6670 13628
rect 6670 13572 6726 13628
rect 6726 13572 6730 13628
rect 6666 13568 6730 13572
rect 17374 13628 17438 13632
rect 17374 13572 17378 13628
rect 17378 13572 17434 13628
rect 17434 13572 17438 13628
rect 17374 13568 17438 13572
rect 17454 13628 17518 13632
rect 17454 13572 17458 13628
rect 17458 13572 17514 13628
rect 17514 13572 17518 13628
rect 17454 13568 17518 13572
rect 17534 13628 17598 13632
rect 17534 13572 17538 13628
rect 17538 13572 17594 13628
rect 17594 13572 17598 13628
rect 17534 13568 17598 13572
rect 17614 13628 17678 13632
rect 17614 13572 17618 13628
rect 17618 13572 17674 13628
rect 17674 13572 17678 13628
rect 17614 13568 17678 13572
rect 28322 13628 28386 13632
rect 28322 13572 28326 13628
rect 28326 13572 28382 13628
rect 28382 13572 28386 13628
rect 28322 13568 28386 13572
rect 28402 13628 28466 13632
rect 28402 13572 28406 13628
rect 28406 13572 28462 13628
rect 28462 13572 28466 13628
rect 28402 13568 28466 13572
rect 28482 13628 28546 13632
rect 28482 13572 28486 13628
rect 28486 13572 28542 13628
rect 28542 13572 28546 13628
rect 28482 13568 28546 13572
rect 28562 13628 28626 13632
rect 28562 13572 28566 13628
rect 28566 13572 28622 13628
rect 28622 13572 28626 13628
rect 28562 13568 28626 13572
rect 39270 13628 39334 13632
rect 39270 13572 39274 13628
rect 39274 13572 39330 13628
rect 39330 13572 39334 13628
rect 39270 13568 39334 13572
rect 39350 13628 39414 13632
rect 39350 13572 39354 13628
rect 39354 13572 39410 13628
rect 39410 13572 39414 13628
rect 39350 13568 39414 13572
rect 39430 13628 39494 13632
rect 39430 13572 39434 13628
rect 39434 13572 39490 13628
rect 39490 13572 39494 13628
rect 39430 13568 39494 13572
rect 39510 13628 39574 13632
rect 39510 13572 39514 13628
rect 39514 13572 39570 13628
rect 39570 13572 39574 13628
rect 39510 13568 39574 13572
rect 11900 13084 11964 13088
rect 11900 13028 11904 13084
rect 11904 13028 11960 13084
rect 11960 13028 11964 13084
rect 11900 13024 11964 13028
rect 11980 13084 12044 13088
rect 11980 13028 11984 13084
rect 11984 13028 12040 13084
rect 12040 13028 12044 13084
rect 11980 13024 12044 13028
rect 12060 13084 12124 13088
rect 12060 13028 12064 13084
rect 12064 13028 12120 13084
rect 12120 13028 12124 13084
rect 12060 13024 12124 13028
rect 12140 13084 12204 13088
rect 12140 13028 12144 13084
rect 12144 13028 12200 13084
rect 12200 13028 12204 13084
rect 12140 13024 12204 13028
rect 22848 13084 22912 13088
rect 22848 13028 22852 13084
rect 22852 13028 22908 13084
rect 22908 13028 22912 13084
rect 22848 13024 22912 13028
rect 22928 13084 22992 13088
rect 22928 13028 22932 13084
rect 22932 13028 22988 13084
rect 22988 13028 22992 13084
rect 22928 13024 22992 13028
rect 23008 13084 23072 13088
rect 23008 13028 23012 13084
rect 23012 13028 23068 13084
rect 23068 13028 23072 13084
rect 23008 13024 23072 13028
rect 23088 13084 23152 13088
rect 23088 13028 23092 13084
rect 23092 13028 23148 13084
rect 23148 13028 23152 13084
rect 23088 13024 23152 13028
rect 33796 13084 33860 13088
rect 33796 13028 33800 13084
rect 33800 13028 33856 13084
rect 33856 13028 33860 13084
rect 33796 13024 33860 13028
rect 33876 13084 33940 13088
rect 33876 13028 33880 13084
rect 33880 13028 33936 13084
rect 33936 13028 33940 13084
rect 33876 13024 33940 13028
rect 33956 13084 34020 13088
rect 33956 13028 33960 13084
rect 33960 13028 34016 13084
rect 34016 13028 34020 13084
rect 33956 13024 34020 13028
rect 34036 13084 34100 13088
rect 34036 13028 34040 13084
rect 34040 13028 34096 13084
rect 34096 13028 34100 13084
rect 34036 13024 34100 13028
rect 44744 13084 44808 13088
rect 44744 13028 44748 13084
rect 44748 13028 44804 13084
rect 44804 13028 44808 13084
rect 44744 13024 44808 13028
rect 44824 13084 44888 13088
rect 44824 13028 44828 13084
rect 44828 13028 44884 13084
rect 44884 13028 44888 13084
rect 44824 13024 44888 13028
rect 44904 13084 44968 13088
rect 44904 13028 44908 13084
rect 44908 13028 44964 13084
rect 44964 13028 44968 13084
rect 44904 13024 44968 13028
rect 44984 13084 45048 13088
rect 44984 13028 44988 13084
rect 44988 13028 45044 13084
rect 45044 13028 45048 13084
rect 44984 13024 45048 13028
rect 6426 12540 6490 12544
rect 6426 12484 6430 12540
rect 6430 12484 6486 12540
rect 6486 12484 6490 12540
rect 6426 12480 6490 12484
rect 6506 12540 6570 12544
rect 6506 12484 6510 12540
rect 6510 12484 6566 12540
rect 6566 12484 6570 12540
rect 6506 12480 6570 12484
rect 6586 12540 6650 12544
rect 6586 12484 6590 12540
rect 6590 12484 6646 12540
rect 6646 12484 6650 12540
rect 6586 12480 6650 12484
rect 6666 12540 6730 12544
rect 6666 12484 6670 12540
rect 6670 12484 6726 12540
rect 6726 12484 6730 12540
rect 6666 12480 6730 12484
rect 17374 12540 17438 12544
rect 17374 12484 17378 12540
rect 17378 12484 17434 12540
rect 17434 12484 17438 12540
rect 17374 12480 17438 12484
rect 17454 12540 17518 12544
rect 17454 12484 17458 12540
rect 17458 12484 17514 12540
rect 17514 12484 17518 12540
rect 17454 12480 17518 12484
rect 17534 12540 17598 12544
rect 17534 12484 17538 12540
rect 17538 12484 17594 12540
rect 17594 12484 17598 12540
rect 17534 12480 17598 12484
rect 17614 12540 17678 12544
rect 17614 12484 17618 12540
rect 17618 12484 17674 12540
rect 17674 12484 17678 12540
rect 17614 12480 17678 12484
rect 28322 12540 28386 12544
rect 28322 12484 28326 12540
rect 28326 12484 28382 12540
rect 28382 12484 28386 12540
rect 28322 12480 28386 12484
rect 28402 12540 28466 12544
rect 28402 12484 28406 12540
rect 28406 12484 28462 12540
rect 28462 12484 28466 12540
rect 28402 12480 28466 12484
rect 28482 12540 28546 12544
rect 28482 12484 28486 12540
rect 28486 12484 28542 12540
rect 28542 12484 28546 12540
rect 28482 12480 28546 12484
rect 28562 12540 28626 12544
rect 28562 12484 28566 12540
rect 28566 12484 28622 12540
rect 28622 12484 28626 12540
rect 28562 12480 28626 12484
rect 39270 12540 39334 12544
rect 39270 12484 39274 12540
rect 39274 12484 39330 12540
rect 39330 12484 39334 12540
rect 39270 12480 39334 12484
rect 39350 12540 39414 12544
rect 39350 12484 39354 12540
rect 39354 12484 39410 12540
rect 39410 12484 39414 12540
rect 39350 12480 39414 12484
rect 39430 12540 39494 12544
rect 39430 12484 39434 12540
rect 39434 12484 39490 12540
rect 39490 12484 39494 12540
rect 39430 12480 39494 12484
rect 39510 12540 39574 12544
rect 39510 12484 39514 12540
rect 39514 12484 39570 12540
rect 39570 12484 39574 12540
rect 39510 12480 39574 12484
rect 11900 11996 11964 12000
rect 11900 11940 11904 11996
rect 11904 11940 11960 11996
rect 11960 11940 11964 11996
rect 11900 11936 11964 11940
rect 11980 11996 12044 12000
rect 11980 11940 11984 11996
rect 11984 11940 12040 11996
rect 12040 11940 12044 11996
rect 11980 11936 12044 11940
rect 12060 11996 12124 12000
rect 12060 11940 12064 11996
rect 12064 11940 12120 11996
rect 12120 11940 12124 11996
rect 12060 11936 12124 11940
rect 12140 11996 12204 12000
rect 12140 11940 12144 11996
rect 12144 11940 12200 11996
rect 12200 11940 12204 11996
rect 12140 11936 12204 11940
rect 22848 11996 22912 12000
rect 22848 11940 22852 11996
rect 22852 11940 22908 11996
rect 22908 11940 22912 11996
rect 22848 11936 22912 11940
rect 22928 11996 22992 12000
rect 22928 11940 22932 11996
rect 22932 11940 22988 11996
rect 22988 11940 22992 11996
rect 22928 11936 22992 11940
rect 23008 11996 23072 12000
rect 23008 11940 23012 11996
rect 23012 11940 23068 11996
rect 23068 11940 23072 11996
rect 23008 11936 23072 11940
rect 23088 11996 23152 12000
rect 23088 11940 23092 11996
rect 23092 11940 23148 11996
rect 23148 11940 23152 11996
rect 23088 11936 23152 11940
rect 33796 11996 33860 12000
rect 33796 11940 33800 11996
rect 33800 11940 33856 11996
rect 33856 11940 33860 11996
rect 33796 11936 33860 11940
rect 33876 11996 33940 12000
rect 33876 11940 33880 11996
rect 33880 11940 33936 11996
rect 33936 11940 33940 11996
rect 33876 11936 33940 11940
rect 33956 11996 34020 12000
rect 33956 11940 33960 11996
rect 33960 11940 34016 11996
rect 34016 11940 34020 11996
rect 33956 11936 34020 11940
rect 34036 11996 34100 12000
rect 34036 11940 34040 11996
rect 34040 11940 34096 11996
rect 34096 11940 34100 11996
rect 34036 11936 34100 11940
rect 44744 11996 44808 12000
rect 44744 11940 44748 11996
rect 44748 11940 44804 11996
rect 44804 11940 44808 11996
rect 44744 11936 44808 11940
rect 44824 11996 44888 12000
rect 44824 11940 44828 11996
rect 44828 11940 44884 11996
rect 44884 11940 44888 11996
rect 44824 11936 44888 11940
rect 44904 11996 44968 12000
rect 44904 11940 44908 11996
rect 44908 11940 44964 11996
rect 44964 11940 44968 11996
rect 44904 11936 44968 11940
rect 44984 11996 45048 12000
rect 44984 11940 44988 11996
rect 44988 11940 45044 11996
rect 45044 11940 45048 11996
rect 44984 11936 45048 11940
rect 6426 11452 6490 11456
rect 6426 11396 6430 11452
rect 6430 11396 6486 11452
rect 6486 11396 6490 11452
rect 6426 11392 6490 11396
rect 6506 11452 6570 11456
rect 6506 11396 6510 11452
rect 6510 11396 6566 11452
rect 6566 11396 6570 11452
rect 6506 11392 6570 11396
rect 6586 11452 6650 11456
rect 6586 11396 6590 11452
rect 6590 11396 6646 11452
rect 6646 11396 6650 11452
rect 6586 11392 6650 11396
rect 6666 11452 6730 11456
rect 6666 11396 6670 11452
rect 6670 11396 6726 11452
rect 6726 11396 6730 11452
rect 6666 11392 6730 11396
rect 17374 11452 17438 11456
rect 17374 11396 17378 11452
rect 17378 11396 17434 11452
rect 17434 11396 17438 11452
rect 17374 11392 17438 11396
rect 17454 11452 17518 11456
rect 17454 11396 17458 11452
rect 17458 11396 17514 11452
rect 17514 11396 17518 11452
rect 17454 11392 17518 11396
rect 17534 11452 17598 11456
rect 17534 11396 17538 11452
rect 17538 11396 17594 11452
rect 17594 11396 17598 11452
rect 17534 11392 17598 11396
rect 17614 11452 17678 11456
rect 17614 11396 17618 11452
rect 17618 11396 17674 11452
rect 17674 11396 17678 11452
rect 17614 11392 17678 11396
rect 28322 11452 28386 11456
rect 28322 11396 28326 11452
rect 28326 11396 28382 11452
rect 28382 11396 28386 11452
rect 28322 11392 28386 11396
rect 28402 11452 28466 11456
rect 28402 11396 28406 11452
rect 28406 11396 28462 11452
rect 28462 11396 28466 11452
rect 28402 11392 28466 11396
rect 28482 11452 28546 11456
rect 28482 11396 28486 11452
rect 28486 11396 28542 11452
rect 28542 11396 28546 11452
rect 28482 11392 28546 11396
rect 28562 11452 28626 11456
rect 28562 11396 28566 11452
rect 28566 11396 28622 11452
rect 28622 11396 28626 11452
rect 28562 11392 28626 11396
rect 39270 11452 39334 11456
rect 39270 11396 39274 11452
rect 39274 11396 39330 11452
rect 39330 11396 39334 11452
rect 39270 11392 39334 11396
rect 39350 11452 39414 11456
rect 39350 11396 39354 11452
rect 39354 11396 39410 11452
rect 39410 11396 39414 11452
rect 39350 11392 39414 11396
rect 39430 11452 39494 11456
rect 39430 11396 39434 11452
rect 39434 11396 39490 11452
rect 39490 11396 39494 11452
rect 39430 11392 39494 11396
rect 39510 11452 39574 11456
rect 39510 11396 39514 11452
rect 39514 11396 39570 11452
rect 39570 11396 39574 11452
rect 39510 11392 39574 11396
rect 11900 10908 11964 10912
rect 11900 10852 11904 10908
rect 11904 10852 11960 10908
rect 11960 10852 11964 10908
rect 11900 10848 11964 10852
rect 11980 10908 12044 10912
rect 11980 10852 11984 10908
rect 11984 10852 12040 10908
rect 12040 10852 12044 10908
rect 11980 10848 12044 10852
rect 12060 10908 12124 10912
rect 12060 10852 12064 10908
rect 12064 10852 12120 10908
rect 12120 10852 12124 10908
rect 12060 10848 12124 10852
rect 12140 10908 12204 10912
rect 12140 10852 12144 10908
rect 12144 10852 12200 10908
rect 12200 10852 12204 10908
rect 12140 10848 12204 10852
rect 22848 10908 22912 10912
rect 22848 10852 22852 10908
rect 22852 10852 22908 10908
rect 22908 10852 22912 10908
rect 22848 10848 22912 10852
rect 22928 10908 22992 10912
rect 22928 10852 22932 10908
rect 22932 10852 22988 10908
rect 22988 10852 22992 10908
rect 22928 10848 22992 10852
rect 23008 10908 23072 10912
rect 23008 10852 23012 10908
rect 23012 10852 23068 10908
rect 23068 10852 23072 10908
rect 23008 10848 23072 10852
rect 23088 10908 23152 10912
rect 23088 10852 23092 10908
rect 23092 10852 23148 10908
rect 23148 10852 23152 10908
rect 23088 10848 23152 10852
rect 33796 10908 33860 10912
rect 33796 10852 33800 10908
rect 33800 10852 33856 10908
rect 33856 10852 33860 10908
rect 33796 10848 33860 10852
rect 33876 10908 33940 10912
rect 33876 10852 33880 10908
rect 33880 10852 33936 10908
rect 33936 10852 33940 10908
rect 33876 10848 33940 10852
rect 33956 10908 34020 10912
rect 33956 10852 33960 10908
rect 33960 10852 34016 10908
rect 34016 10852 34020 10908
rect 33956 10848 34020 10852
rect 34036 10908 34100 10912
rect 34036 10852 34040 10908
rect 34040 10852 34096 10908
rect 34096 10852 34100 10908
rect 34036 10848 34100 10852
rect 44744 10908 44808 10912
rect 44744 10852 44748 10908
rect 44748 10852 44804 10908
rect 44804 10852 44808 10908
rect 44744 10848 44808 10852
rect 44824 10908 44888 10912
rect 44824 10852 44828 10908
rect 44828 10852 44884 10908
rect 44884 10852 44888 10908
rect 44824 10848 44888 10852
rect 44904 10908 44968 10912
rect 44904 10852 44908 10908
rect 44908 10852 44964 10908
rect 44964 10852 44968 10908
rect 44904 10848 44968 10852
rect 44984 10908 45048 10912
rect 44984 10852 44988 10908
rect 44988 10852 45044 10908
rect 45044 10852 45048 10908
rect 44984 10848 45048 10852
rect 6426 10364 6490 10368
rect 6426 10308 6430 10364
rect 6430 10308 6486 10364
rect 6486 10308 6490 10364
rect 6426 10304 6490 10308
rect 6506 10364 6570 10368
rect 6506 10308 6510 10364
rect 6510 10308 6566 10364
rect 6566 10308 6570 10364
rect 6506 10304 6570 10308
rect 6586 10364 6650 10368
rect 6586 10308 6590 10364
rect 6590 10308 6646 10364
rect 6646 10308 6650 10364
rect 6586 10304 6650 10308
rect 6666 10364 6730 10368
rect 6666 10308 6670 10364
rect 6670 10308 6726 10364
rect 6726 10308 6730 10364
rect 6666 10304 6730 10308
rect 17374 10364 17438 10368
rect 17374 10308 17378 10364
rect 17378 10308 17434 10364
rect 17434 10308 17438 10364
rect 17374 10304 17438 10308
rect 17454 10364 17518 10368
rect 17454 10308 17458 10364
rect 17458 10308 17514 10364
rect 17514 10308 17518 10364
rect 17454 10304 17518 10308
rect 17534 10364 17598 10368
rect 17534 10308 17538 10364
rect 17538 10308 17594 10364
rect 17594 10308 17598 10364
rect 17534 10304 17598 10308
rect 17614 10364 17678 10368
rect 17614 10308 17618 10364
rect 17618 10308 17674 10364
rect 17674 10308 17678 10364
rect 17614 10304 17678 10308
rect 28322 10364 28386 10368
rect 28322 10308 28326 10364
rect 28326 10308 28382 10364
rect 28382 10308 28386 10364
rect 28322 10304 28386 10308
rect 28402 10364 28466 10368
rect 28402 10308 28406 10364
rect 28406 10308 28462 10364
rect 28462 10308 28466 10364
rect 28402 10304 28466 10308
rect 28482 10364 28546 10368
rect 28482 10308 28486 10364
rect 28486 10308 28542 10364
rect 28542 10308 28546 10364
rect 28482 10304 28546 10308
rect 28562 10364 28626 10368
rect 28562 10308 28566 10364
rect 28566 10308 28622 10364
rect 28622 10308 28626 10364
rect 28562 10304 28626 10308
rect 39270 10364 39334 10368
rect 39270 10308 39274 10364
rect 39274 10308 39330 10364
rect 39330 10308 39334 10364
rect 39270 10304 39334 10308
rect 39350 10364 39414 10368
rect 39350 10308 39354 10364
rect 39354 10308 39410 10364
rect 39410 10308 39414 10364
rect 39350 10304 39414 10308
rect 39430 10364 39494 10368
rect 39430 10308 39434 10364
rect 39434 10308 39490 10364
rect 39490 10308 39494 10364
rect 39430 10304 39494 10308
rect 39510 10364 39574 10368
rect 39510 10308 39514 10364
rect 39514 10308 39570 10364
rect 39570 10308 39574 10364
rect 39510 10304 39574 10308
rect 11900 9820 11964 9824
rect 11900 9764 11904 9820
rect 11904 9764 11960 9820
rect 11960 9764 11964 9820
rect 11900 9760 11964 9764
rect 11980 9820 12044 9824
rect 11980 9764 11984 9820
rect 11984 9764 12040 9820
rect 12040 9764 12044 9820
rect 11980 9760 12044 9764
rect 12060 9820 12124 9824
rect 12060 9764 12064 9820
rect 12064 9764 12120 9820
rect 12120 9764 12124 9820
rect 12060 9760 12124 9764
rect 12140 9820 12204 9824
rect 12140 9764 12144 9820
rect 12144 9764 12200 9820
rect 12200 9764 12204 9820
rect 12140 9760 12204 9764
rect 22848 9820 22912 9824
rect 22848 9764 22852 9820
rect 22852 9764 22908 9820
rect 22908 9764 22912 9820
rect 22848 9760 22912 9764
rect 22928 9820 22992 9824
rect 22928 9764 22932 9820
rect 22932 9764 22988 9820
rect 22988 9764 22992 9820
rect 22928 9760 22992 9764
rect 23008 9820 23072 9824
rect 23008 9764 23012 9820
rect 23012 9764 23068 9820
rect 23068 9764 23072 9820
rect 23008 9760 23072 9764
rect 23088 9820 23152 9824
rect 23088 9764 23092 9820
rect 23092 9764 23148 9820
rect 23148 9764 23152 9820
rect 23088 9760 23152 9764
rect 33796 9820 33860 9824
rect 33796 9764 33800 9820
rect 33800 9764 33856 9820
rect 33856 9764 33860 9820
rect 33796 9760 33860 9764
rect 33876 9820 33940 9824
rect 33876 9764 33880 9820
rect 33880 9764 33936 9820
rect 33936 9764 33940 9820
rect 33876 9760 33940 9764
rect 33956 9820 34020 9824
rect 33956 9764 33960 9820
rect 33960 9764 34016 9820
rect 34016 9764 34020 9820
rect 33956 9760 34020 9764
rect 34036 9820 34100 9824
rect 34036 9764 34040 9820
rect 34040 9764 34096 9820
rect 34096 9764 34100 9820
rect 34036 9760 34100 9764
rect 44744 9820 44808 9824
rect 44744 9764 44748 9820
rect 44748 9764 44804 9820
rect 44804 9764 44808 9820
rect 44744 9760 44808 9764
rect 44824 9820 44888 9824
rect 44824 9764 44828 9820
rect 44828 9764 44884 9820
rect 44884 9764 44888 9820
rect 44824 9760 44888 9764
rect 44904 9820 44968 9824
rect 44904 9764 44908 9820
rect 44908 9764 44964 9820
rect 44964 9764 44968 9820
rect 44904 9760 44968 9764
rect 44984 9820 45048 9824
rect 44984 9764 44988 9820
rect 44988 9764 45044 9820
rect 45044 9764 45048 9820
rect 44984 9760 45048 9764
rect 6426 9276 6490 9280
rect 6426 9220 6430 9276
rect 6430 9220 6486 9276
rect 6486 9220 6490 9276
rect 6426 9216 6490 9220
rect 6506 9276 6570 9280
rect 6506 9220 6510 9276
rect 6510 9220 6566 9276
rect 6566 9220 6570 9276
rect 6506 9216 6570 9220
rect 6586 9276 6650 9280
rect 6586 9220 6590 9276
rect 6590 9220 6646 9276
rect 6646 9220 6650 9276
rect 6586 9216 6650 9220
rect 6666 9276 6730 9280
rect 6666 9220 6670 9276
rect 6670 9220 6726 9276
rect 6726 9220 6730 9276
rect 6666 9216 6730 9220
rect 17374 9276 17438 9280
rect 17374 9220 17378 9276
rect 17378 9220 17434 9276
rect 17434 9220 17438 9276
rect 17374 9216 17438 9220
rect 17454 9276 17518 9280
rect 17454 9220 17458 9276
rect 17458 9220 17514 9276
rect 17514 9220 17518 9276
rect 17454 9216 17518 9220
rect 17534 9276 17598 9280
rect 17534 9220 17538 9276
rect 17538 9220 17594 9276
rect 17594 9220 17598 9276
rect 17534 9216 17598 9220
rect 17614 9276 17678 9280
rect 17614 9220 17618 9276
rect 17618 9220 17674 9276
rect 17674 9220 17678 9276
rect 17614 9216 17678 9220
rect 28322 9276 28386 9280
rect 28322 9220 28326 9276
rect 28326 9220 28382 9276
rect 28382 9220 28386 9276
rect 28322 9216 28386 9220
rect 28402 9276 28466 9280
rect 28402 9220 28406 9276
rect 28406 9220 28462 9276
rect 28462 9220 28466 9276
rect 28402 9216 28466 9220
rect 28482 9276 28546 9280
rect 28482 9220 28486 9276
rect 28486 9220 28542 9276
rect 28542 9220 28546 9276
rect 28482 9216 28546 9220
rect 28562 9276 28626 9280
rect 28562 9220 28566 9276
rect 28566 9220 28622 9276
rect 28622 9220 28626 9276
rect 28562 9216 28626 9220
rect 39270 9276 39334 9280
rect 39270 9220 39274 9276
rect 39274 9220 39330 9276
rect 39330 9220 39334 9276
rect 39270 9216 39334 9220
rect 39350 9276 39414 9280
rect 39350 9220 39354 9276
rect 39354 9220 39410 9276
rect 39410 9220 39414 9276
rect 39350 9216 39414 9220
rect 39430 9276 39494 9280
rect 39430 9220 39434 9276
rect 39434 9220 39490 9276
rect 39490 9220 39494 9276
rect 39430 9216 39494 9220
rect 39510 9276 39574 9280
rect 39510 9220 39514 9276
rect 39514 9220 39570 9276
rect 39570 9220 39574 9276
rect 39510 9216 39574 9220
rect 11900 8732 11964 8736
rect 11900 8676 11904 8732
rect 11904 8676 11960 8732
rect 11960 8676 11964 8732
rect 11900 8672 11964 8676
rect 11980 8732 12044 8736
rect 11980 8676 11984 8732
rect 11984 8676 12040 8732
rect 12040 8676 12044 8732
rect 11980 8672 12044 8676
rect 12060 8732 12124 8736
rect 12060 8676 12064 8732
rect 12064 8676 12120 8732
rect 12120 8676 12124 8732
rect 12060 8672 12124 8676
rect 12140 8732 12204 8736
rect 12140 8676 12144 8732
rect 12144 8676 12200 8732
rect 12200 8676 12204 8732
rect 12140 8672 12204 8676
rect 22848 8732 22912 8736
rect 22848 8676 22852 8732
rect 22852 8676 22908 8732
rect 22908 8676 22912 8732
rect 22848 8672 22912 8676
rect 22928 8732 22992 8736
rect 22928 8676 22932 8732
rect 22932 8676 22988 8732
rect 22988 8676 22992 8732
rect 22928 8672 22992 8676
rect 23008 8732 23072 8736
rect 23008 8676 23012 8732
rect 23012 8676 23068 8732
rect 23068 8676 23072 8732
rect 23008 8672 23072 8676
rect 23088 8732 23152 8736
rect 23088 8676 23092 8732
rect 23092 8676 23148 8732
rect 23148 8676 23152 8732
rect 23088 8672 23152 8676
rect 33796 8732 33860 8736
rect 33796 8676 33800 8732
rect 33800 8676 33856 8732
rect 33856 8676 33860 8732
rect 33796 8672 33860 8676
rect 33876 8732 33940 8736
rect 33876 8676 33880 8732
rect 33880 8676 33936 8732
rect 33936 8676 33940 8732
rect 33876 8672 33940 8676
rect 33956 8732 34020 8736
rect 33956 8676 33960 8732
rect 33960 8676 34016 8732
rect 34016 8676 34020 8732
rect 33956 8672 34020 8676
rect 34036 8732 34100 8736
rect 34036 8676 34040 8732
rect 34040 8676 34096 8732
rect 34096 8676 34100 8732
rect 34036 8672 34100 8676
rect 44744 8732 44808 8736
rect 44744 8676 44748 8732
rect 44748 8676 44804 8732
rect 44804 8676 44808 8732
rect 44744 8672 44808 8676
rect 44824 8732 44888 8736
rect 44824 8676 44828 8732
rect 44828 8676 44884 8732
rect 44884 8676 44888 8732
rect 44824 8672 44888 8676
rect 44904 8732 44968 8736
rect 44904 8676 44908 8732
rect 44908 8676 44964 8732
rect 44964 8676 44968 8732
rect 44904 8672 44968 8676
rect 44984 8732 45048 8736
rect 44984 8676 44988 8732
rect 44988 8676 45044 8732
rect 45044 8676 45048 8732
rect 44984 8672 45048 8676
rect 6426 8188 6490 8192
rect 6426 8132 6430 8188
rect 6430 8132 6486 8188
rect 6486 8132 6490 8188
rect 6426 8128 6490 8132
rect 6506 8188 6570 8192
rect 6506 8132 6510 8188
rect 6510 8132 6566 8188
rect 6566 8132 6570 8188
rect 6506 8128 6570 8132
rect 6586 8188 6650 8192
rect 6586 8132 6590 8188
rect 6590 8132 6646 8188
rect 6646 8132 6650 8188
rect 6586 8128 6650 8132
rect 6666 8188 6730 8192
rect 6666 8132 6670 8188
rect 6670 8132 6726 8188
rect 6726 8132 6730 8188
rect 6666 8128 6730 8132
rect 17374 8188 17438 8192
rect 17374 8132 17378 8188
rect 17378 8132 17434 8188
rect 17434 8132 17438 8188
rect 17374 8128 17438 8132
rect 17454 8188 17518 8192
rect 17454 8132 17458 8188
rect 17458 8132 17514 8188
rect 17514 8132 17518 8188
rect 17454 8128 17518 8132
rect 17534 8188 17598 8192
rect 17534 8132 17538 8188
rect 17538 8132 17594 8188
rect 17594 8132 17598 8188
rect 17534 8128 17598 8132
rect 17614 8188 17678 8192
rect 17614 8132 17618 8188
rect 17618 8132 17674 8188
rect 17674 8132 17678 8188
rect 17614 8128 17678 8132
rect 28322 8188 28386 8192
rect 28322 8132 28326 8188
rect 28326 8132 28382 8188
rect 28382 8132 28386 8188
rect 28322 8128 28386 8132
rect 28402 8188 28466 8192
rect 28402 8132 28406 8188
rect 28406 8132 28462 8188
rect 28462 8132 28466 8188
rect 28402 8128 28466 8132
rect 28482 8188 28546 8192
rect 28482 8132 28486 8188
rect 28486 8132 28542 8188
rect 28542 8132 28546 8188
rect 28482 8128 28546 8132
rect 28562 8188 28626 8192
rect 28562 8132 28566 8188
rect 28566 8132 28622 8188
rect 28622 8132 28626 8188
rect 28562 8128 28626 8132
rect 39270 8188 39334 8192
rect 39270 8132 39274 8188
rect 39274 8132 39330 8188
rect 39330 8132 39334 8188
rect 39270 8128 39334 8132
rect 39350 8188 39414 8192
rect 39350 8132 39354 8188
rect 39354 8132 39410 8188
rect 39410 8132 39414 8188
rect 39350 8128 39414 8132
rect 39430 8188 39494 8192
rect 39430 8132 39434 8188
rect 39434 8132 39490 8188
rect 39490 8132 39494 8188
rect 39430 8128 39494 8132
rect 39510 8188 39574 8192
rect 39510 8132 39514 8188
rect 39514 8132 39570 8188
rect 39570 8132 39574 8188
rect 39510 8128 39574 8132
rect 11900 7644 11964 7648
rect 11900 7588 11904 7644
rect 11904 7588 11960 7644
rect 11960 7588 11964 7644
rect 11900 7584 11964 7588
rect 11980 7644 12044 7648
rect 11980 7588 11984 7644
rect 11984 7588 12040 7644
rect 12040 7588 12044 7644
rect 11980 7584 12044 7588
rect 12060 7644 12124 7648
rect 12060 7588 12064 7644
rect 12064 7588 12120 7644
rect 12120 7588 12124 7644
rect 12060 7584 12124 7588
rect 12140 7644 12204 7648
rect 12140 7588 12144 7644
rect 12144 7588 12200 7644
rect 12200 7588 12204 7644
rect 12140 7584 12204 7588
rect 22848 7644 22912 7648
rect 22848 7588 22852 7644
rect 22852 7588 22908 7644
rect 22908 7588 22912 7644
rect 22848 7584 22912 7588
rect 22928 7644 22992 7648
rect 22928 7588 22932 7644
rect 22932 7588 22988 7644
rect 22988 7588 22992 7644
rect 22928 7584 22992 7588
rect 23008 7644 23072 7648
rect 23008 7588 23012 7644
rect 23012 7588 23068 7644
rect 23068 7588 23072 7644
rect 23008 7584 23072 7588
rect 23088 7644 23152 7648
rect 23088 7588 23092 7644
rect 23092 7588 23148 7644
rect 23148 7588 23152 7644
rect 23088 7584 23152 7588
rect 33796 7644 33860 7648
rect 33796 7588 33800 7644
rect 33800 7588 33856 7644
rect 33856 7588 33860 7644
rect 33796 7584 33860 7588
rect 33876 7644 33940 7648
rect 33876 7588 33880 7644
rect 33880 7588 33936 7644
rect 33936 7588 33940 7644
rect 33876 7584 33940 7588
rect 33956 7644 34020 7648
rect 33956 7588 33960 7644
rect 33960 7588 34016 7644
rect 34016 7588 34020 7644
rect 33956 7584 34020 7588
rect 34036 7644 34100 7648
rect 34036 7588 34040 7644
rect 34040 7588 34096 7644
rect 34096 7588 34100 7644
rect 34036 7584 34100 7588
rect 44744 7644 44808 7648
rect 44744 7588 44748 7644
rect 44748 7588 44804 7644
rect 44804 7588 44808 7644
rect 44744 7584 44808 7588
rect 44824 7644 44888 7648
rect 44824 7588 44828 7644
rect 44828 7588 44884 7644
rect 44884 7588 44888 7644
rect 44824 7584 44888 7588
rect 44904 7644 44968 7648
rect 44904 7588 44908 7644
rect 44908 7588 44964 7644
rect 44964 7588 44968 7644
rect 44904 7584 44968 7588
rect 44984 7644 45048 7648
rect 44984 7588 44988 7644
rect 44988 7588 45044 7644
rect 45044 7588 45048 7644
rect 44984 7584 45048 7588
rect 6426 7100 6490 7104
rect 6426 7044 6430 7100
rect 6430 7044 6486 7100
rect 6486 7044 6490 7100
rect 6426 7040 6490 7044
rect 6506 7100 6570 7104
rect 6506 7044 6510 7100
rect 6510 7044 6566 7100
rect 6566 7044 6570 7100
rect 6506 7040 6570 7044
rect 6586 7100 6650 7104
rect 6586 7044 6590 7100
rect 6590 7044 6646 7100
rect 6646 7044 6650 7100
rect 6586 7040 6650 7044
rect 6666 7100 6730 7104
rect 6666 7044 6670 7100
rect 6670 7044 6726 7100
rect 6726 7044 6730 7100
rect 6666 7040 6730 7044
rect 17374 7100 17438 7104
rect 17374 7044 17378 7100
rect 17378 7044 17434 7100
rect 17434 7044 17438 7100
rect 17374 7040 17438 7044
rect 17454 7100 17518 7104
rect 17454 7044 17458 7100
rect 17458 7044 17514 7100
rect 17514 7044 17518 7100
rect 17454 7040 17518 7044
rect 17534 7100 17598 7104
rect 17534 7044 17538 7100
rect 17538 7044 17594 7100
rect 17594 7044 17598 7100
rect 17534 7040 17598 7044
rect 17614 7100 17678 7104
rect 17614 7044 17618 7100
rect 17618 7044 17674 7100
rect 17674 7044 17678 7100
rect 17614 7040 17678 7044
rect 28322 7100 28386 7104
rect 28322 7044 28326 7100
rect 28326 7044 28382 7100
rect 28382 7044 28386 7100
rect 28322 7040 28386 7044
rect 28402 7100 28466 7104
rect 28402 7044 28406 7100
rect 28406 7044 28462 7100
rect 28462 7044 28466 7100
rect 28402 7040 28466 7044
rect 28482 7100 28546 7104
rect 28482 7044 28486 7100
rect 28486 7044 28542 7100
rect 28542 7044 28546 7100
rect 28482 7040 28546 7044
rect 28562 7100 28626 7104
rect 28562 7044 28566 7100
rect 28566 7044 28622 7100
rect 28622 7044 28626 7100
rect 28562 7040 28626 7044
rect 39270 7100 39334 7104
rect 39270 7044 39274 7100
rect 39274 7044 39330 7100
rect 39330 7044 39334 7100
rect 39270 7040 39334 7044
rect 39350 7100 39414 7104
rect 39350 7044 39354 7100
rect 39354 7044 39410 7100
rect 39410 7044 39414 7100
rect 39350 7040 39414 7044
rect 39430 7100 39494 7104
rect 39430 7044 39434 7100
rect 39434 7044 39490 7100
rect 39490 7044 39494 7100
rect 39430 7040 39494 7044
rect 39510 7100 39574 7104
rect 39510 7044 39514 7100
rect 39514 7044 39570 7100
rect 39570 7044 39574 7100
rect 39510 7040 39574 7044
rect 11900 6556 11964 6560
rect 11900 6500 11904 6556
rect 11904 6500 11960 6556
rect 11960 6500 11964 6556
rect 11900 6496 11964 6500
rect 11980 6556 12044 6560
rect 11980 6500 11984 6556
rect 11984 6500 12040 6556
rect 12040 6500 12044 6556
rect 11980 6496 12044 6500
rect 12060 6556 12124 6560
rect 12060 6500 12064 6556
rect 12064 6500 12120 6556
rect 12120 6500 12124 6556
rect 12060 6496 12124 6500
rect 12140 6556 12204 6560
rect 12140 6500 12144 6556
rect 12144 6500 12200 6556
rect 12200 6500 12204 6556
rect 12140 6496 12204 6500
rect 22848 6556 22912 6560
rect 22848 6500 22852 6556
rect 22852 6500 22908 6556
rect 22908 6500 22912 6556
rect 22848 6496 22912 6500
rect 22928 6556 22992 6560
rect 22928 6500 22932 6556
rect 22932 6500 22988 6556
rect 22988 6500 22992 6556
rect 22928 6496 22992 6500
rect 23008 6556 23072 6560
rect 23008 6500 23012 6556
rect 23012 6500 23068 6556
rect 23068 6500 23072 6556
rect 23008 6496 23072 6500
rect 23088 6556 23152 6560
rect 23088 6500 23092 6556
rect 23092 6500 23148 6556
rect 23148 6500 23152 6556
rect 23088 6496 23152 6500
rect 33796 6556 33860 6560
rect 33796 6500 33800 6556
rect 33800 6500 33856 6556
rect 33856 6500 33860 6556
rect 33796 6496 33860 6500
rect 33876 6556 33940 6560
rect 33876 6500 33880 6556
rect 33880 6500 33936 6556
rect 33936 6500 33940 6556
rect 33876 6496 33940 6500
rect 33956 6556 34020 6560
rect 33956 6500 33960 6556
rect 33960 6500 34016 6556
rect 34016 6500 34020 6556
rect 33956 6496 34020 6500
rect 34036 6556 34100 6560
rect 34036 6500 34040 6556
rect 34040 6500 34096 6556
rect 34096 6500 34100 6556
rect 34036 6496 34100 6500
rect 44744 6556 44808 6560
rect 44744 6500 44748 6556
rect 44748 6500 44804 6556
rect 44804 6500 44808 6556
rect 44744 6496 44808 6500
rect 44824 6556 44888 6560
rect 44824 6500 44828 6556
rect 44828 6500 44884 6556
rect 44884 6500 44888 6556
rect 44824 6496 44888 6500
rect 44904 6556 44968 6560
rect 44904 6500 44908 6556
rect 44908 6500 44964 6556
rect 44964 6500 44968 6556
rect 44904 6496 44968 6500
rect 44984 6556 45048 6560
rect 44984 6500 44988 6556
rect 44988 6500 45044 6556
rect 45044 6500 45048 6556
rect 44984 6496 45048 6500
rect 6426 6012 6490 6016
rect 6426 5956 6430 6012
rect 6430 5956 6486 6012
rect 6486 5956 6490 6012
rect 6426 5952 6490 5956
rect 6506 6012 6570 6016
rect 6506 5956 6510 6012
rect 6510 5956 6566 6012
rect 6566 5956 6570 6012
rect 6506 5952 6570 5956
rect 6586 6012 6650 6016
rect 6586 5956 6590 6012
rect 6590 5956 6646 6012
rect 6646 5956 6650 6012
rect 6586 5952 6650 5956
rect 6666 6012 6730 6016
rect 6666 5956 6670 6012
rect 6670 5956 6726 6012
rect 6726 5956 6730 6012
rect 6666 5952 6730 5956
rect 17374 6012 17438 6016
rect 17374 5956 17378 6012
rect 17378 5956 17434 6012
rect 17434 5956 17438 6012
rect 17374 5952 17438 5956
rect 17454 6012 17518 6016
rect 17454 5956 17458 6012
rect 17458 5956 17514 6012
rect 17514 5956 17518 6012
rect 17454 5952 17518 5956
rect 17534 6012 17598 6016
rect 17534 5956 17538 6012
rect 17538 5956 17594 6012
rect 17594 5956 17598 6012
rect 17534 5952 17598 5956
rect 17614 6012 17678 6016
rect 17614 5956 17618 6012
rect 17618 5956 17674 6012
rect 17674 5956 17678 6012
rect 17614 5952 17678 5956
rect 28322 6012 28386 6016
rect 28322 5956 28326 6012
rect 28326 5956 28382 6012
rect 28382 5956 28386 6012
rect 28322 5952 28386 5956
rect 28402 6012 28466 6016
rect 28402 5956 28406 6012
rect 28406 5956 28462 6012
rect 28462 5956 28466 6012
rect 28402 5952 28466 5956
rect 28482 6012 28546 6016
rect 28482 5956 28486 6012
rect 28486 5956 28542 6012
rect 28542 5956 28546 6012
rect 28482 5952 28546 5956
rect 28562 6012 28626 6016
rect 28562 5956 28566 6012
rect 28566 5956 28622 6012
rect 28622 5956 28626 6012
rect 28562 5952 28626 5956
rect 39270 6012 39334 6016
rect 39270 5956 39274 6012
rect 39274 5956 39330 6012
rect 39330 5956 39334 6012
rect 39270 5952 39334 5956
rect 39350 6012 39414 6016
rect 39350 5956 39354 6012
rect 39354 5956 39410 6012
rect 39410 5956 39414 6012
rect 39350 5952 39414 5956
rect 39430 6012 39494 6016
rect 39430 5956 39434 6012
rect 39434 5956 39490 6012
rect 39490 5956 39494 6012
rect 39430 5952 39494 5956
rect 39510 6012 39574 6016
rect 39510 5956 39514 6012
rect 39514 5956 39570 6012
rect 39570 5956 39574 6012
rect 39510 5952 39574 5956
rect 11900 5468 11964 5472
rect 11900 5412 11904 5468
rect 11904 5412 11960 5468
rect 11960 5412 11964 5468
rect 11900 5408 11964 5412
rect 11980 5468 12044 5472
rect 11980 5412 11984 5468
rect 11984 5412 12040 5468
rect 12040 5412 12044 5468
rect 11980 5408 12044 5412
rect 12060 5468 12124 5472
rect 12060 5412 12064 5468
rect 12064 5412 12120 5468
rect 12120 5412 12124 5468
rect 12060 5408 12124 5412
rect 12140 5468 12204 5472
rect 12140 5412 12144 5468
rect 12144 5412 12200 5468
rect 12200 5412 12204 5468
rect 12140 5408 12204 5412
rect 22848 5468 22912 5472
rect 22848 5412 22852 5468
rect 22852 5412 22908 5468
rect 22908 5412 22912 5468
rect 22848 5408 22912 5412
rect 22928 5468 22992 5472
rect 22928 5412 22932 5468
rect 22932 5412 22988 5468
rect 22988 5412 22992 5468
rect 22928 5408 22992 5412
rect 23008 5468 23072 5472
rect 23008 5412 23012 5468
rect 23012 5412 23068 5468
rect 23068 5412 23072 5468
rect 23008 5408 23072 5412
rect 23088 5468 23152 5472
rect 23088 5412 23092 5468
rect 23092 5412 23148 5468
rect 23148 5412 23152 5468
rect 23088 5408 23152 5412
rect 33796 5468 33860 5472
rect 33796 5412 33800 5468
rect 33800 5412 33856 5468
rect 33856 5412 33860 5468
rect 33796 5408 33860 5412
rect 33876 5468 33940 5472
rect 33876 5412 33880 5468
rect 33880 5412 33936 5468
rect 33936 5412 33940 5468
rect 33876 5408 33940 5412
rect 33956 5468 34020 5472
rect 33956 5412 33960 5468
rect 33960 5412 34016 5468
rect 34016 5412 34020 5468
rect 33956 5408 34020 5412
rect 34036 5468 34100 5472
rect 34036 5412 34040 5468
rect 34040 5412 34096 5468
rect 34096 5412 34100 5468
rect 34036 5408 34100 5412
rect 44744 5468 44808 5472
rect 44744 5412 44748 5468
rect 44748 5412 44804 5468
rect 44804 5412 44808 5468
rect 44744 5408 44808 5412
rect 44824 5468 44888 5472
rect 44824 5412 44828 5468
rect 44828 5412 44884 5468
rect 44884 5412 44888 5468
rect 44824 5408 44888 5412
rect 44904 5468 44968 5472
rect 44904 5412 44908 5468
rect 44908 5412 44964 5468
rect 44964 5412 44968 5468
rect 44904 5408 44968 5412
rect 44984 5468 45048 5472
rect 44984 5412 44988 5468
rect 44988 5412 45044 5468
rect 45044 5412 45048 5468
rect 44984 5408 45048 5412
rect 6426 4924 6490 4928
rect 6426 4868 6430 4924
rect 6430 4868 6486 4924
rect 6486 4868 6490 4924
rect 6426 4864 6490 4868
rect 6506 4924 6570 4928
rect 6506 4868 6510 4924
rect 6510 4868 6566 4924
rect 6566 4868 6570 4924
rect 6506 4864 6570 4868
rect 6586 4924 6650 4928
rect 6586 4868 6590 4924
rect 6590 4868 6646 4924
rect 6646 4868 6650 4924
rect 6586 4864 6650 4868
rect 6666 4924 6730 4928
rect 6666 4868 6670 4924
rect 6670 4868 6726 4924
rect 6726 4868 6730 4924
rect 6666 4864 6730 4868
rect 17374 4924 17438 4928
rect 17374 4868 17378 4924
rect 17378 4868 17434 4924
rect 17434 4868 17438 4924
rect 17374 4864 17438 4868
rect 17454 4924 17518 4928
rect 17454 4868 17458 4924
rect 17458 4868 17514 4924
rect 17514 4868 17518 4924
rect 17454 4864 17518 4868
rect 17534 4924 17598 4928
rect 17534 4868 17538 4924
rect 17538 4868 17594 4924
rect 17594 4868 17598 4924
rect 17534 4864 17598 4868
rect 17614 4924 17678 4928
rect 17614 4868 17618 4924
rect 17618 4868 17674 4924
rect 17674 4868 17678 4924
rect 17614 4864 17678 4868
rect 28322 4924 28386 4928
rect 28322 4868 28326 4924
rect 28326 4868 28382 4924
rect 28382 4868 28386 4924
rect 28322 4864 28386 4868
rect 28402 4924 28466 4928
rect 28402 4868 28406 4924
rect 28406 4868 28462 4924
rect 28462 4868 28466 4924
rect 28402 4864 28466 4868
rect 28482 4924 28546 4928
rect 28482 4868 28486 4924
rect 28486 4868 28542 4924
rect 28542 4868 28546 4924
rect 28482 4864 28546 4868
rect 28562 4924 28626 4928
rect 28562 4868 28566 4924
rect 28566 4868 28622 4924
rect 28622 4868 28626 4924
rect 28562 4864 28626 4868
rect 39270 4924 39334 4928
rect 39270 4868 39274 4924
rect 39274 4868 39330 4924
rect 39330 4868 39334 4924
rect 39270 4864 39334 4868
rect 39350 4924 39414 4928
rect 39350 4868 39354 4924
rect 39354 4868 39410 4924
rect 39410 4868 39414 4924
rect 39350 4864 39414 4868
rect 39430 4924 39494 4928
rect 39430 4868 39434 4924
rect 39434 4868 39490 4924
rect 39490 4868 39494 4924
rect 39430 4864 39494 4868
rect 39510 4924 39574 4928
rect 39510 4868 39514 4924
rect 39514 4868 39570 4924
rect 39570 4868 39574 4924
rect 39510 4864 39574 4868
rect 11900 4380 11964 4384
rect 11900 4324 11904 4380
rect 11904 4324 11960 4380
rect 11960 4324 11964 4380
rect 11900 4320 11964 4324
rect 11980 4380 12044 4384
rect 11980 4324 11984 4380
rect 11984 4324 12040 4380
rect 12040 4324 12044 4380
rect 11980 4320 12044 4324
rect 12060 4380 12124 4384
rect 12060 4324 12064 4380
rect 12064 4324 12120 4380
rect 12120 4324 12124 4380
rect 12060 4320 12124 4324
rect 12140 4380 12204 4384
rect 12140 4324 12144 4380
rect 12144 4324 12200 4380
rect 12200 4324 12204 4380
rect 12140 4320 12204 4324
rect 22848 4380 22912 4384
rect 22848 4324 22852 4380
rect 22852 4324 22908 4380
rect 22908 4324 22912 4380
rect 22848 4320 22912 4324
rect 22928 4380 22992 4384
rect 22928 4324 22932 4380
rect 22932 4324 22988 4380
rect 22988 4324 22992 4380
rect 22928 4320 22992 4324
rect 23008 4380 23072 4384
rect 23008 4324 23012 4380
rect 23012 4324 23068 4380
rect 23068 4324 23072 4380
rect 23008 4320 23072 4324
rect 23088 4380 23152 4384
rect 23088 4324 23092 4380
rect 23092 4324 23148 4380
rect 23148 4324 23152 4380
rect 23088 4320 23152 4324
rect 33796 4380 33860 4384
rect 33796 4324 33800 4380
rect 33800 4324 33856 4380
rect 33856 4324 33860 4380
rect 33796 4320 33860 4324
rect 33876 4380 33940 4384
rect 33876 4324 33880 4380
rect 33880 4324 33936 4380
rect 33936 4324 33940 4380
rect 33876 4320 33940 4324
rect 33956 4380 34020 4384
rect 33956 4324 33960 4380
rect 33960 4324 34016 4380
rect 34016 4324 34020 4380
rect 33956 4320 34020 4324
rect 34036 4380 34100 4384
rect 34036 4324 34040 4380
rect 34040 4324 34096 4380
rect 34096 4324 34100 4380
rect 34036 4320 34100 4324
rect 44744 4380 44808 4384
rect 44744 4324 44748 4380
rect 44748 4324 44804 4380
rect 44804 4324 44808 4380
rect 44744 4320 44808 4324
rect 44824 4380 44888 4384
rect 44824 4324 44828 4380
rect 44828 4324 44884 4380
rect 44884 4324 44888 4380
rect 44824 4320 44888 4324
rect 44904 4380 44968 4384
rect 44904 4324 44908 4380
rect 44908 4324 44964 4380
rect 44964 4324 44968 4380
rect 44904 4320 44968 4324
rect 44984 4380 45048 4384
rect 44984 4324 44988 4380
rect 44988 4324 45044 4380
rect 45044 4324 45048 4380
rect 44984 4320 45048 4324
rect 6426 3836 6490 3840
rect 6426 3780 6430 3836
rect 6430 3780 6486 3836
rect 6486 3780 6490 3836
rect 6426 3776 6490 3780
rect 6506 3836 6570 3840
rect 6506 3780 6510 3836
rect 6510 3780 6566 3836
rect 6566 3780 6570 3836
rect 6506 3776 6570 3780
rect 6586 3836 6650 3840
rect 6586 3780 6590 3836
rect 6590 3780 6646 3836
rect 6646 3780 6650 3836
rect 6586 3776 6650 3780
rect 6666 3836 6730 3840
rect 6666 3780 6670 3836
rect 6670 3780 6726 3836
rect 6726 3780 6730 3836
rect 6666 3776 6730 3780
rect 17374 3836 17438 3840
rect 17374 3780 17378 3836
rect 17378 3780 17434 3836
rect 17434 3780 17438 3836
rect 17374 3776 17438 3780
rect 17454 3836 17518 3840
rect 17454 3780 17458 3836
rect 17458 3780 17514 3836
rect 17514 3780 17518 3836
rect 17454 3776 17518 3780
rect 17534 3836 17598 3840
rect 17534 3780 17538 3836
rect 17538 3780 17594 3836
rect 17594 3780 17598 3836
rect 17534 3776 17598 3780
rect 17614 3836 17678 3840
rect 17614 3780 17618 3836
rect 17618 3780 17674 3836
rect 17674 3780 17678 3836
rect 17614 3776 17678 3780
rect 28322 3836 28386 3840
rect 28322 3780 28326 3836
rect 28326 3780 28382 3836
rect 28382 3780 28386 3836
rect 28322 3776 28386 3780
rect 28402 3836 28466 3840
rect 28402 3780 28406 3836
rect 28406 3780 28462 3836
rect 28462 3780 28466 3836
rect 28402 3776 28466 3780
rect 28482 3836 28546 3840
rect 28482 3780 28486 3836
rect 28486 3780 28542 3836
rect 28542 3780 28546 3836
rect 28482 3776 28546 3780
rect 28562 3836 28626 3840
rect 28562 3780 28566 3836
rect 28566 3780 28622 3836
rect 28622 3780 28626 3836
rect 28562 3776 28626 3780
rect 39270 3836 39334 3840
rect 39270 3780 39274 3836
rect 39274 3780 39330 3836
rect 39330 3780 39334 3836
rect 39270 3776 39334 3780
rect 39350 3836 39414 3840
rect 39350 3780 39354 3836
rect 39354 3780 39410 3836
rect 39410 3780 39414 3836
rect 39350 3776 39414 3780
rect 39430 3836 39494 3840
rect 39430 3780 39434 3836
rect 39434 3780 39490 3836
rect 39490 3780 39494 3836
rect 39430 3776 39494 3780
rect 39510 3836 39574 3840
rect 39510 3780 39514 3836
rect 39514 3780 39570 3836
rect 39570 3780 39574 3836
rect 39510 3776 39574 3780
rect 11900 3292 11964 3296
rect 11900 3236 11904 3292
rect 11904 3236 11960 3292
rect 11960 3236 11964 3292
rect 11900 3232 11964 3236
rect 11980 3292 12044 3296
rect 11980 3236 11984 3292
rect 11984 3236 12040 3292
rect 12040 3236 12044 3292
rect 11980 3232 12044 3236
rect 12060 3292 12124 3296
rect 12060 3236 12064 3292
rect 12064 3236 12120 3292
rect 12120 3236 12124 3292
rect 12060 3232 12124 3236
rect 12140 3292 12204 3296
rect 12140 3236 12144 3292
rect 12144 3236 12200 3292
rect 12200 3236 12204 3292
rect 12140 3232 12204 3236
rect 22848 3292 22912 3296
rect 22848 3236 22852 3292
rect 22852 3236 22908 3292
rect 22908 3236 22912 3292
rect 22848 3232 22912 3236
rect 22928 3292 22992 3296
rect 22928 3236 22932 3292
rect 22932 3236 22988 3292
rect 22988 3236 22992 3292
rect 22928 3232 22992 3236
rect 23008 3292 23072 3296
rect 23008 3236 23012 3292
rect 23012 3236 23068 3292
rect 23068 3236 23072 3292
rect 23008 3232 23072 3236
rect 23088 3292 23152 3296
rect 23088 3236 23092 3292
rect 23092 3236 23148 3292
rect 23148 3236 23152 3292
rect 23088 3232 23152 3236
rect 33796 3292 33860 3296
rect 33796 3236 33800 3292
rect 33800 3236 33856 3292
rect 33856 3236 33860 3292
rect 33796 3232 33860 3236
rect 33876 3292 33940 3296
rect 33876 3236 33880 3292
rect 33880 3236 33936 3292
rect 33936 3236 33940 3292
rect 33876 3232 33940 3236
rect 33956 3292 34020 3296
rect 33956 3236 33960 3292
rect 33960 3236 34016 3292
rect 34016 3236 34020 3292
rect 33956 3232 34020 3236
rect 34036 3292 34100 3296
rect 34036 3236 34040 3292
rect 34040 3236 34096 3292
rect 34096 3236 34100 3292
rect 34036 3232 34100 3236
rect 44744 3292 44808 3296
rect 44744 3236 44748 3292
rect 44748 3236 44804 3292
rect 44804 3236 44808 3292
rect 44744 3232 44808 3236
rect 44824 3292 44888 3296
rect 44824 3236 44828 3292
rect 44828 3236 44884 3292
rect 44884 3236 44888 3292
rect 44824 3232 44888 3236
rect 44904 3292 44968 3296
rect 44904 3236 44908 3292
rect 44908 3236 44964 3292
rect 44964 3236 44968 3292
rect 44904 3232 44968 3236
rect 44984 3292 45048 3296
rect 44984 3236 44988 3292
rect 44988 3236 45044 3292
rect 45044 3236 45048 3292
rect 44984 3232 45048 3236
rect 6426 2748 6490 2752
rect 6426 2692 6430 2748
rect 6430 2692 6486 2748
rect 6486 2692 6490 2748
rect 6426 2688 6490 2692
rect 6506 2748 6570 2752
rect 6506 2692 6510 2748
rect 6510 2692 6566 2748
rect 6566 2692 6570 2748
rect 6506 2688 6570 2692
rect 6586 2748 6650 2752
rect 6586 2692 6590 2748
rect 6590 2692 6646 2748
rect 6646 2692 6650 2748
rect 6586 2688 6650 2692
rect 6666 2748 6730 2752
rect 6666 2692 6670 2748
rect 6670 2692 6726 2748
rect 6726 2692 6730 2748
rect 6666 2688 6730 2692
rect 17374 2748 17438 2752
rect 17374 2692 17378 2748
rect 17378 2692 17434 2748
rect 17434 2692 17438 2748
rect 17374 2688 17438 2692
rect 17454 2748 17518 2752
rect 17454 2692 17458 2748
rect 17458 2692 17514 2748
rect 17514 2692 17518 2748
rect 17454 2688 17518 2692
rect 17534 2748 17598 2752
rect 17534 2692 17538 2748
rect 17538 2692 17594 2748
rect 17594 2692 17598 2748
rect 17534 2688 17598 2692
rect 17614 2748 17678 2752
rect 17614 2692 17618 2748
rect 17618 2692 17674 2748
rect 17674 2692 17678 2748
rect 17614 2688 17678 2692
rect 28322 2748 28386 2752
rect 28322 2692 28326 2748
rect 28326 2692 28382 2748
rect 28382 2692 28386 2748
rect 28322 2688 28386 2692
rect 28402 2748 28466 2752
rect 28402 2692 28406 2748
rect 28406 2692 28462 2748
rect 28462 2692 28466 2748
rect 28402 2688 28466 2692
rect 28482 2748 28546 2752
rect 28482 2692 28486 2748
rect 28486 2692 28542 2748
rect 28542 2692 28546 2748
rect 28482 2688 28546 2692
rect 28562 2748 28626 2752
rect 28562 2692 28566 2748
rect 28566 2692 28622 2748
rect 28622 2692 28626 2748
rect 28562 2688 28626 2692
rect 39270 2748 39334 2752
rect 39270 2692 39274 2748
rect 39274 2692 39330 2748
rect 39330 2692 39334 2748
rect 39270 2688 39334 2692
rect 39350 2748 39414 2752
rect 39350 2692 39354 2748
rect 39354 2692 39410 2748
rect 39410 2692 39414 2748
rect 39350 2688 39414 2692
rect 39430 2748 39494 2752
rect 39430 2692 39434 2748
rect 39434 2692 39490 2748
rect 39490 2692 39494 2748
rect 39430 2688 39494 2692
rect 39510 2748 39574 2752
rect 39510 2692 39514 2748
rect 39514 2692 39570 2748
rect 39570 2692 39574 2748
rect 39510 2688 39574 2692
rect 11900 2204 11964 2208
rect 11900 2148 11904 2204
rect 11904 2148 11960 2204
rect 11960 2148 11964 2204
rect 11900 2144 11964 2148
rect 11980 2204 12044 2208
rect 11980 2148 11984 2204
rect 11984 2148 12040 2204
rect 12040 2148 12044 2204
rect 11980 2144 12044 2148
rect 12060 2204 12124 2208
rect 12060 2148 12064 2204
rect 12064 2148 12120 2204
rect 12120 2148 12124 2204
rect 12060 2144 12124 2148
rect 12140 2204 12204 2208
rect 12140 2148 12144 2204
rect 12144 2148 12200 2204
rect 12200 2148 12204 2204
rect 12140 2144 12204 2148
rect 22848 2204 22912 2208
rect 22848 2148 22852 2204
rect 22852 2148 22908 2204
rect 22908 2148 22912 2204
rect 22848 2144 22912 2148
rect 22928 2204 22992 2208
rect 22928 2148 22932 2204
rect 22932 2148 22988 2204
rect 22988 2148 22992 2204
rect 22928 2144 22992 2148
rect 23008 2204 23072 2208
rect 23008 2148 23012 2204
rect 23012 2148 23068 2204
rect 23068 2148 23072 2204
rect 23008 2144 23072 2148
rect 23088 2204 23152 2208
rect 23088 2148 23092 2204
rect 23092 2148 23148 2204
rect 23148 2148 23152 2204
rect 23088 2144 23152 2148
rect 33796 2204 33860 2208
rect 33796 2148 33800 2204
rect 33800 2148 33856 2204
rect 33856 2148 33860 2204
rect 33796 2144 33860 2148
rect 33876 2204 33940 2208
rect 33876 2148 33880 2204
rect 33880 2148 33936 2204
rect 33936 2148 33940 2204
rect 33876 2144 33940 2148
rect 33956 2204 34020 2208
rect 33956 2148 33960 2204
rect 33960 2148 34016 2204
rect 34016 2148 34020 2204
rect 33956 2144 34020 2148
rect 34036 2204 34100 2208
rect 34036 2148 34040 2204
rect 34040 2148 34096 2204
rect 34096 2148 34100 2204
rect 34036 2144 34100 2148
rect 44744 2204 44808 2208
rect 44744 2148 44748 2204
rect 44748 2148 44804 2204
rect 44804 2148 44808 2204
rect 44744 2144 44808 2148
rect 44824 2204 44888 2208
rect 44824 2148 44828 2204
rect 44828 2148 44884 2204
rect 44884 2148 44888 2204
rect 44824 2144 44888 2148
rect 44904 2204 44968 2208
rect 44904 2148 44908 2204
rect 44908 2148 44964 2204
rect 44964 2148 44968 2204
rect 44904 2144 44968 2148
rect 44984 2204 45048 2208
rect 44984 2148 44988 2204
rect 44988 2148 45044 2204
rect 45044 2148 45048 2204
rect 44984 2144 45048 2148
<< metal4 >>
rect 6418 16896 6738 17456
rect 6418 16832 6426 16896
rect 6490 16832 6506 16896
rect 6570 16832 6586 16896
rect 6650 16832 6666 16896
rect 6730 16832 6738 16896
rect 6418 15808 6738 16832
rect 6418 15744 6426 15808
rect 6490 15744 6506 15808
rect 6570 15744 6586 15808
rect 6650 15744 6666 15808
rect 6730 15744 6738 15808
rect 6418 14720 6738 15744
rect 6418 14656 6426 14720
rect 6490 14656 6506 14720
rect 6570 14656 6586 14720
rect 6650 14656 6666 14720
rect 6730 14656 6738 14720
rect 6418 13632 6738 14656
rect 6418 13568 6426 13632
rect 6490 13568 6506 13632
rect 6570 13568 6586 13632
rect 6650 13568 6666 13632
rect 6730 13568 6738 13632
rect 6418 12544 6738 13568
rect 6418 12480 6426 12544
rect 6490 12480 6506 12544
rect 6570 12480 6586 12544
rect 6650 12480 6666 12544
rect 6730 12480 6738 12544
rect 6418 11456 6738 12480
rect 6418 11392 6426 11456
rect 6490 11392 6506 11456
rect 6570 11392 6586 11456
rect 6650 11392 6666 11456
rect 6730 11392 6738 11456
rect 6418 10368 6738 11392
rect 6418 10304 6426 10368
rect 6490 10304 6506 10368
rect 6570 10304 6586 10368
rect 6650 10304 6666 10368
rect 6730 10304 6738 10368
rect 6418 9280 6738 10304
rect 6418 9216 6426 9280
rect 6490 9216 6506 9280
rect 6570 9216 6586 9280
rect 6650 9216 6666 9280
rect 6730 9216 6738 9280
rect 6418 8192 6738 9216
rect 6418 8128 6426 8192
rect 6490 8128 6506 8192
rect 6570 8128 6586 8192
rect 6650 8128 6666 8192
rect 6730 8128 6738 8192
rect 6418 7104 6738 8128
rect 6418 7040 6426 7104
rect 6490 7040 6506 7104
rect 6570 7040 6586 7104
rect 6650 7040 6666 7104
rect 6730 7040 6738 7104
rect 6418 6016 6738 7040
rect 6418 5952 6426 6016
rect 6490 5952 6506 6016
rect 6570 5952 6586 6016
rect 6650 5952 6666 6016
rect 6730 5952 6738 6016
rect 6418 4928 6738 5952
rect 6418 4864 6426 4928
rect 6490 4864 6506 4928
rect 6570 4864 6586 4928
rect 6650 4864 6666 4928
rect 6730 4864 6738 4928
rect 6418 3840 6738 4864
rect 6418 3776 6426 3840
rect 6490 3776 6506 3840
rect 6570 3776 6586 3840
rect 6650 3776 6666 3840
rect 6730 3776 6738 3840
rect 6418 2752 6738 3776
rect 6418 2688 6426 2752
rect 6490 2688 6506 2752
rect 6570 2688 6586 2752
rect 6650 2688 6666 2752
rect 6730 2688 6738 2752
rect 6418 2128 6738 2688
rect 11892 17440 12212 17456
rect 11892 17376 11900 17440
rect 11964 17376 11980 17440
rect 12044 17376 12060 17440
rect 12124 17376 12140 17440
rect 12204 17376 12212 17440
rect 11892 16352 12212 17376
rect 11892 16288 11900 16352
rect 11964 16288 11980 16352
rect 12044 16288 12060 16352
rect 12124 16288 12140 16352
rect 12204 16288 12212 16352
rect 11892 15264 12212 16288
rect 11892 15200 11900 15264
rect 11964 15200 11980 15264
rect 12044 15200 12060 15264
rect 12124 15200 12140 15264
rect 12204 15200 12212 15264
rect 11892 14176 12212 15200
rect 11892 14112 11900 14176
rect 11964 14112 11980 14176
rect 12044 14112 12060 14176
rect 12124 14112 12140 14176
rect 12204 14112 12212 14176
rect 11892 13088 12212 14112
rect 11892 13024 11900 13088
rect 11964 13024 11980 13088
rect 12044 13024 12060 13088
rect 12124 13024 12140 13088
rect 12204 13024 12212 13088
rect 11892 12000 12212 13024
rect 11892 11936 11900 12000
rect 11964 11936 11980 12000
rect 12044 11936 12060 12000
rect 12124 11936 12140 12000
rect 12204 11936 12212 12000
rect 11892 10912 12212 11936
rect 11892 10848 11900 10912
rect 11964 10848 11980 10912
rect 12044 10848 12060 10912
rect 12124 10848 12140 10912
rect 12204 10848 12212 10912
rect 11892 9824 12212 10848
rect 11892 9760 11900 9824
rect 11964 9760 11980 9824
rect 12044 9760 12060 9824
rect 12124 9760 12140 9824
rect 12204 9760 12212 9824
rect 11892 8736 12212 9760
rect 11892 8672 11900 8736
rect 11964 8672 11980 8736
rect 12044 8672 12060 8736
rect 12124 8672 12140 8736
rect 12204 8672 12212 8736
rect 11892 7648 12212 8672
rect 11892 7584 11900 7648
rect 11964 7584 11980 7648
rect 12044 7584 12060 7648
rect 12124 7584 12140 7648
rect 12204 7584 12212 7648
rect 11892 6560 12212 7584
rect 11892 6496 11900 6560
rect 11964 6496 11980 6560
rect 12044 6496 12060 6560
rect 12124 6496 12140 6560
rect 12204 6496 12212 6560
rect 11892 5472 12212 6496
rect 11892 5408 11900 5472
rect 11964 5408 11980 5472
rect 12044 5408 12060 5472
rect 12124 5408 12140 5472
rect 12204 5408 12212 5472
rect 11892 4384 12212 5408
rect 11892 4320 11900 4384
rect 11964 4320 11980 4384
rect 12044 4320 12060 4384
rect 12124 4320 12140 4384
rect 12204 4320 12212 4384
rect 11892 3296 12212 4320
rect 11892 3232 11900 3296
rect 11964 3232 11980 3296
rect 12044 3232 12060 3296
rect 12124 3232 12140 3296
rect 12204 3232 12212 3296
rect 11892 2208 12212 3232
rect 11892 2144 11900 2208
rect 11964 2144 11980 2208
rect 12044 2144 12060 2208
rect 12124 2144 12140 2208
rect 12204 2144 12212 2208
rect 11892 2128 12212 2144
rect 17366 16896 17686 17456
rect 17366 16832 17374 16896
rect 17438 16832 17454 16896
rect 17518 16832 17534 16896
rect 17598 16832 17614 16896
rect 17678 16832 17686 16896
rect 17366 15808 17686 16832
rect 17366 15744 17374 15808
rect 17438 15744 17454 15808
rect 17518 15744 17534 15808
rect 17598 15744 17614 15808
rect 17678 15744 17686 15808
rect 17366 14720 17686 15744
rect 17366 14656 17374 14720
rect 17438 14656 17454 14720
rect 17518 14656 17534 14720
rect 17598 14656 17614 14720
rect 17678 14656 17686 14720
rect 17366 13632 17686 14656
rect 17366 13568 17374 13632
rect 17438 13568 17454 13632
rect 17518 13568 17534 13632
rect 17598 13568 17614 13632
rect 17678 13568 17686 13632
rect 17366 12544 17686 13568
rect 17366 12480 17374 12544
rect 17438 12480 17454 12544
rect 17518 12480 17534 12544
rect 17598 12480 17614 12544
rect 17678 12480 17686 12544
rect 17366 11456 17686 12480
rect 17366 11392 17374 11456
rect 17438 11392 17454 11456
rect 17518 11392 17534 11456
rect 17598 11392 17614 11456
rect 17678 11392 17686 11456
rect 17366 10368 17686 11392
rect 17366 10304 17374 10368
rect 17438 10304 17454 10368
rect 17518 10304 17534 10368
rect 17598 10304 17614 10368
rect 17678 10304 17686 10368
rect 17366 9280 17686 10304
rect 17366 9216 17374 9280
rect 17438 9216 17454 9280
rect 17518 9216 17534 9280
rect 17598 9216 17614 9280
rect 17678 9216 17686 9280
rect 17366 8192 17686 9216
rect 17366 8128 17374 8192
rect 17438 8128 17454 8192
rect 17518 8128 17534 8192
rect 17598 8128 17614 8192
rect 17678 8128 17686 8192
rect 17366 7104 17686 8128
rect 17366 7040 17374 7104
rect 17438 7040 17454 7104
rect 17518 7040 17534 7104
rect 17598 7040 17614 7104
rect 17678 7040 17686 7104
rect 17366 6016 17686 7040
rect 17366 5952 17374 6016
rect 17438 5952 17454 6016
rect 17518 5952 17534 6016
rect 17598 5952 17614 6016
rect 17678 5952 17686 6016
rect 17366 4928 17686 5952
rect 17366 4864 17374 4928
rect 17438 4864 17454 4928
rect 17518 4864 17534 4928
rect 17598 4864 17614 4928
rect 17678 4864 17686 4928
rect 17366 3840 17686 4864
rect 17366 3776 17374 3840
rect 17438 3776 17454 3840
rect 17518 3776 17534 3840
rect 17598 3776 17614 3840
rect 17678 3776 17686 3840
rect 17366 2752 17686 3776
rect 17366 2688 17374 2752
rect 17438 2688 17454 2752
rect 17518 2688 17534 2752
rect 17598 2688 17614 2752
rect 17678 2688 17686 2752
rect 17366 2128 17686 2688
rect 22840 17440 23160 17456
rect 22840 17376 22848 17440
rect 22912 17376 22928 17440
rect 22992 17376 23008 17440
rect 23072 17376 23088 17440
rect 23152 17376 23160 17440
rect 22840 16352 23160 17376
rect 22840 16288 22848 16352
rect 22912 16288 22928 16352
rect 22992 16288 23008 16352
rect 23072 16288 23088 16352
rect 23152 16288 23160 16352
rect 22840 15264 23160 16288
rect 22840 15200 22848 15264
rect 22912 15200 22928 15264
rect 22992 15200 23008 15264
rect 23072 15200 23088 15264
rect 23152 15200 23160 15264
rect 22840 14176 23160 15200
rect 22840 14112 22848 14176
rect 22912 14112 22928 14176
rect 22992 14112 23008 14176
rect 23072 14112 23088 14176
rect 23152 14112 23160 14176
rect 22840 13088 23160 14112
rect 22840 13024 22848 13088
rect 22912 13024 22928 13088
rect 22992 13024 23008 13088
rect 23072 13024 23088 13088
rect 23152 13024 23160 13088
rect 22840 12000 23160 13024
rect 22840 11936 22848 12000
rect 22912 11936 22928 12000
rect 22992 11936 23008 12000
rect 23072 11936 23088 12000
rect 23152 11936 23160 12000
rect 22840 10912 23160 11936
rect 22840 10848 22848 10912
rect 22912 10848 22928 10912
rect 22992 10848 23008 10912
rect 23072 10848 23088 10912
rect 23152 10848 23160 10912
rect 22840 9824 23160 10848
rect 22840 9760 22848 9824
rect 22912 9760 22928 9824
rect 22992 9760 23008 9824
rect 23072 9760 23088 9824
rect 23152 9760 23160 9824
rect 22840 8736 23160 9760
rect 22840 8672 22848 8736
rect 22912 8672 22928 8736
rect 22992 8672 23008 8736
rect 23072 8672 23088 8736
rect 23152 8672 23160 8736
rect 22840 7648 23160 8672
rect 22840 7584 22848 7648
rect 22912 7584 22928 7648
rect 22992 7584 23008 7648
rect 23072 7584 23088 7648
rect 23152 7584 23160 7648
rect 22840 6560 23160 7584
rect 22840 6496 22848 6560
rect 22912 6496 22928 6560
rect 22992 6496 23008 6560
rect 23072 6496 23088 6560
rect 23152 6496 23160 6560
rect 22840 5472 23160 6496
rect 22840 5408 22848 5472
rect 22912 5408 22928 5472
rect 22992 5408 23008 5472
rect 23072 5408 23088 5472
rect 23152 5408 23160 5472
rect 22840 4384 23160 5408
rect 22840 4320 22848 4384
rect 22912 4320 22928 4384
rect 22992 4320 23008 4384
rect 23072 4320 23088 4384
rect 23152 4320 23160 4384
rect 22840 3296 23160 4320
rect 22840 3232 22848 3296
rect 22912 3232 22928 3296
rect 22992 3232 23008 3296
rect 23072 3232 23088 3296
rect 23152 3232 23160 3296
rect 22840 2208 23160 3232
rect 22840 2144 22848 2208
rect 22912 2144 22928 2208
rect 22992 2144 23008 2208
rect 23072 2144 23088 2208
rect 23152 2144 23160 2208
rect 22840 2128 23160 2144
rect 28314 16896 28634 17456
rect 28314 16832 28322 16896
rect 28386 16832 28402 16896
rect 28466 16832 28482 16896
rect 28546 16832 28562 16896
rect 28626 16832 28634 16896
rect 28314 15808 28634 16832
rect 28314 15744 28322 15808
rect 28386 15744 28402 15808
rect 28466 15744 28482 15808
rect 28546 15744 28562 15808
rect 28626 15744 28634 15808
rect 28314 14720 28634 15744
rect 28314 14656 28322 14720
rect 28386 14656 28402 14720
rect 28466 14656 28482 14720
rect 28546 14656 28562 14720
rect 28626 14656 28634 14720
rect 28314 13632 28634 14656
rect 28314 13568 28322 13632
rect 28386 13568 28402 13632
rect 28466 13568 28482 13632
rect 28546 13568 28562 13632
rect 28626 13568 28634 13632
rect 28314 12544 28634 13568
rect 28314 12480 28322 12544
rect 28386 12480 28402 12544
rect 28466 12480 28482 12544
rect 28546 12480 28562 12544
rect 28626 12480 28634 12544
rect 28314 11456 28634 12480
rect 28314 11392 28322 11456
rect 28386 11392 28402 11456
rect 28466 11392 28482 11456
rect 28546 11392 28562 11456
rect 28626 11392 28634 11456
rect 28314 10368 28634 11392
rect 28314 10304 28322 10368
rect 28386 10304 28402 10368
rect 28466 10304 28482 10368
rect 28546 10304 28562 10368
rect 28626 10304 28634 10368
rect 28314 9280 28634 10304
rect 28314 9216 28322 9280
rect 28386 9216 28402 9280
rect 28466 9216 28482 9280
rect 28546 9216 28562 9280
rect 28626 9216 28634 9280
rect 28314 8192 28634 9216
rect 28314 8128 28322 8192
rect 28386 8128 28402 8192
rect 28466 8128 28482 8192
rect 28546 8128 28562 8192
rect 28626 8128 28634 8192
rect 28314 7104 28634 8128
rect 28314 7040 28322 7104
rect 28386 7040 28402 7104
rect 28466 7040 28482 7104
rect 28546 7040 28562 7104
rect 28626 7040 28634 7104
rect 28314 6016 28634 7040
rect 28314 5952 28322 6016
rect 28386 5952 28402 6016
rect 28466 5952 28482 6016
rect 28546 5952 28562 6016
rect 28626 5952 28634 6016
rect 28314 4928 28634 5952
rect 28314 4864 28322 4928
rect 28386 4864 28402 4928
rect 28466 4864 28482 4928
rect 28546 4864 28562 4928
rect 28626 4864 28634 4928
rect 28314 3840 28634 4864
rect 28314 3776 28322 3840
rect 28386 3776 28402 3840
rect 28466 3776 28482 3840
rect 28546 3776 28562 3840
rect 28626 3776 28634 3840
rect 28314 2752 28634 3776
rect 28314 2688 28322 2752
rect 28386 2688 28402 2752
rect 28466 2688 28482 2752
rect 28546 2688 28562 2752
rect 28626 2688 28634 2752
rect 28314 2128 28634 2688
rect 33788 17440 34108 17456
rect 33788 17376 33796 17440
rect 33860 17376 33876 17440
rect 33940 17376 33956 17440
rect 34020 17376 34036 17440
rect 34100 17376 34108 17440
rect 33788 16352 34108 17376
rect 33788 16288 33796 16352
rect 33860 16288 33876 16352
rect 33940 16288 33956 16352
rect 34020 16288 34036 16352
rect 34100 16288 34108 16352
rect 33788 15264 34108 16288
rect 33788 15200 33796 15264
rect 33860 15200 33876 15264
rect 33940 15200 33956 15264
rect 34020 15200 34036 15264
rect 34100 15200 34108 15264
rect 33788 14176 34108 15200
rect 33788 14112 33796 14176
rect 33860 14112 33876 14176
rect 33940 14112 33956 14176
rect 34020 14112 34036 14176
rect 34100 14112 34108 14176
rect 33788 13088 34108 14112
rect 33788 13024 33796 13088
rect 33860 13024 33876 13088
rect 33940 13024 33956 13088
rect 34020 13024 34036 13088
rect 34100 13024 34108 13088
rect 33788 12000 34108 13024
rect 33788 11936 33796 12000
rect 33860 11936 33876 12000
rect 33940 11936 33956 12000
rect 34020 11936 34036 12000
rect 34100 11936 34108 12000
rect 33788 10912 34108 11936
rect 33788 10848 33796 10912
rect 33860 10848 33876 10912
rect 33940 10848 33956 10912
rect 34020 10848 34036 10912
rect 34100 10848 34108 10912
rect 33788 9824 34108 10848
rect 33788 9760 33796 9824
rect 33860 9760 33876 9824
rect 33940 9760 33956 9824
rect 34020 9760 34036 9824
rect 34100 9760 34108 9824
rect 33788 8736 34108 9760
rect 33788 8672 33796 8736
rect 33860 8672 33876 8736
rect 33940 8672 33956 8736
rect 34020 8672 34036 8736
rect 34100 8672 34108 8736
rect 33788 7648 34108 8672
rect 33788 7584 33796 7648
rect 33860 7584 33876 7648
rect 33940 7584 33956 7648
rect 34020 7584 34036 7648
rect 34100 7584 34108 7648
rect 33788 6560 34108 7584
rect 33788 6496 33796 6560
rect 33860 6496 33876 6560
rect 33940 6496 33956 6560
rect 34020 6496 34036 6560
rect 34100 6496 34108 6560
rect 33788 5472 34108 6496
rect 33788 5408 33796 5472
rect 33860 5408 33876 5472
rect 33940 5408 33956 5472
rect 34020 5408 34036 5472
rect 34100 5408 34108 5472
rect 33788 4384 34108 5408
rect 33788 4320 33796 4384
rect 33860 4320 33876 4384
rect 33940 4320 33956 4384
rect 34020 4320 34036 4384
rect 34100 4320 34108 4384
rect 33788 3296 34108 4320
rect 33788 3232 33796 3296
rect 33860 3232 33876 3296
rect 33940 3232 33956 3296
rect 34020 3232 34036 3296
rect 34100 3232 34108 3296
rect 33788 2208 34108 3232
rect 33788 2144 33796 2208
rect 33860 2144 33876 2208
rect 33940 2144 33956 2208
rect 34020 2144 34036 2208
rect 34100 2144 34108 2208
rect 33788 2128 34108 2144
rect 39262 16896 39582 17456
rect 39262 16832 39270 16896
rect 39334 16832 39350 16896
rect 39414 16832 39430 16896
rect 39494 16832 39510 16896
rect 39574 16832 39582 16896
rect 39262 15808 39582 16832
rect 39262 15744 39270 15808
rect 39334 15744 39350 15808
rect 39414 15744 39430 15808
rect 39494 15744 39510 15808
rect 39574 15744 39582 15808
rect 39262 14720 39582 15744
rect 39262 14656 39270 14720
rect 39334 14656 39350 14720
rect 39414 14656 39430 14720
rect 39494 14656 39510 14720
rect 39574 14656 39582 14720
rect 39262 13632 39582 14656
rect 39262 13568 39270 13632
rect 39334 13568 39350 13632
rect 39414 13568 39430 13632
rect 39494 13568 39510 13632
rect 39574 13568 39582 13632
rect 39262 12544 39582 13568
rect 39262 12480 39270 12544
rect 39334 12480 39350 12544
rect 39414 12480 39430 12544
rect 39494 12480 39510 12544
rect 39574 12480 39582 12544
rect 39262 11456 39582 12480
rect 39262 11392 39270 11456
rect 39334 11392 39350 11456
rect 39414 11392 39430 11456
rect 39494 11392 39510 11456
rect 39574 11392 39582 11456
rect 39262 10368 39582 11392
rect 39262 10304 39270 10368
rect 39334 10304 39350 10368
rect 39414 10304 39430 10368
rect 39494 10304 39510 10368
rect 39574 10304 39582 10368
rect 39262 9280 39582 10304
rect 39262 9216 39270 9280
rect 39334 9216 39350 9280
rect 39414 9216 39430 9280
rect 39494 9216 39510 9280
rect 39574 9216 39582 9280
rect 39262 8192 39582 9216
rect 39262 8128 39270 8192
rect 39334 8128 39350 8192
rect 39414 8128 39430 8192
rect 39494 8128 39510 8192
rect 39574 8128 39582 8192
rect 39262 7104 39582 8128
rect 39262 7040 39270 7104
rect 39334 7040 39350 7104
rect 39414 7040 39430 7104
rect 39494 7040 39510 7104
rect 39574 7040 39582 7104
rect 39262 6016 39582 7040
rect 39262 5952 39270 6016
rect 39334 5952 39350 6016
rect 39414 5952 39430 6016
rect 39494 5952 39510 6016
rect 39574 5952 39582 6016
rect 39262 4928 39582 5952
rect 39262 4864 39270 4928
rect 39334 4864 39350 4928
rect 39414 4864 39430 4928
rect 39494 4864 39510 4928
rect 39574 4864 39582 4928
rect 39262 3840 39582 4864
rect 39262 3776 39270 3840
rect 39334 3776 39350 3840
rect 39414 3776 39430 3840
rect 39494 3776 39510 3840
rect 39574 3776 39582 3840
rect 39262 2752 39582 3776
rect 39262 2688 39270 2752
rect 39334 2688 39350 2752
rect 39414 2688 39430 2752
rect 39494 2688 39510 2752
rect 39574 2688 39582 2752
rect 39262 2128 39582 2688
rect 44736 17440 45056 17456
rect 44736 17376 44744 17440
rect 44808 17376 44824 17440
rect 44888 17376 44904 17440
rect 44968 17376 44984 17440
rect 45048 17376 45056 17440
rect 44736 16352 45056 17376
rect 44736 16288 44744 16352
rect 44808 16288 44824 16352
rect 44888 16288 44904 16352
rect 44968 16288 44984 16352
rect 45048 16288 45056 16352
rect 44736 15264 45056 16288
rect 44736 15200 44744 15264
rect 44808 15200 44824 15264
rect 44888 15200 44904 15264
rect 44968 15200 44984 15264
rect 45048 15200 45056 15264
rect 44736 14176 45056 15200
rect 44736 14112 44744 14176
rect 44808 14112 44824 14176
rect 44888 14112 44904 14176
rect 44968 14112 44984 14176
rect 45048 14112 45056 14176
rect 44736 13088 45056 14112
rect 44736 13024 44744 13088
rect 44808 13024 44824 13088
rect 44888 13024 44904 13088
rect 44968 13024 44984 13088
rect 45048 13024 45056 13088
rect 44736 12000 45056 13024
rect 44736 11936 44744 12000
rect 44808 11936 44824 12000
rect 44888 11936 44904 12000
rect 44968 11936 44984 12000
rect 45048 11936 45056 12000
rect 44736 10912 45056 11936
rect 44736 10848 44744 10912
rect 44808 10848 44824 10912
rect 44888 10848 44904 10912
rect 44968 10848 44984 10912
rect 45048 10848 45056 10912
rect 44736 9824 45056 10848
rect 44736 9760 44744 9824
rect 44808 9760 44824 9824
rect 44888 9760 44904 9824
rect 44968 9760 44984 9824
rect 45048 9760 45056 9824
rect 44736 8736 45056 9760
rect 44736 8672 44744 8736
rect 44808 8672 44824 8736
rect 44888 8672 44904 8736
rect 44968 8672 44984 8736
rect 45048 8672 45056 8736
rect 44736 7648 45056 8672
rect 44736 7584 44744 7648
rect 44808 7584 44824 7648
rect 44888 7584 44904 7648
rect 44968 7584 44984 7648
rect 45048 7584 45056 7648
rect 44736 6560 45056 7584
rect 44736 6496 44744 6560
rect 44808 6496 44824 6560
rect 44888 6496 44904 6560
rect 44968 6496 44984 6560
rect 45048 6496 45056 6560
rect 44736 5472 45056 6496
rect 44736 5408 44744 5472
rect 44808 5408 44824 5472
rect 44888 5408 44904 5472
rect 44968 5408 44984 5472
rect 45048 5408 45056 5472
rect 44736 4384 45056 5408
rect 44736 4320 44744 4384
rect 44808 4320 44824 4384
rect 44888 4320 44904 4384
rect 44968 4320 44984 4384
rect 45048 4320 45056 4384
rect 44736 3296 45056 4320
rect 44736 3232 44744 3296
rect 44808 3232 44824 3296
rect 44888 3232 44904 3296
rect 44968 3232 44984 3296
rect 45048 3232 45056 3296
rect 44736 2208 45056 3232
rect 44736 2144 44744 2208
rect 44808 2144 44824 2208
rect 44888 2144 44904 2208
rect 44968 2144 44984 2208
rect 45048 2144 45056 2208
rect 44736 2128 45056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_0 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20148 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1649977179
transform 1 0 33948 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1649977179
transform 1 0 43240 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4048 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71
timestamp 1649977179
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76
timestamp 1649977179
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_116
timestamp 1649977179
transform 1 0 11776 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128
timestamp 1649977179
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1649977179
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146
timestamp 1649977179
transform 1 0 14536 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1649977179
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_202
timestamp 1649977179
transform 1 0 19688 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_210
timestamp 1649977179
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1649977179
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1649977179
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_238
timestamp 1649977179
transform 1 0 23000 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1649977179
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_256
timestamp 1649977179
transform 1 0 24656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_268
timestamp 1649977179
transform 1 0 25760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1649977179
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_287
timestamp 1649977179
transform 1 0 27508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_299
timestamp 1649977179
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1649977179
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_312
timestamp 1649977179
transform 1 0 29808 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1649977179
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1649977179
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_345
timestamp 1649977179
transform 1 0 32844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1649977179
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1649977179
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_373
timestamp 1649977179
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_378
timestamp 1649977179
transform 1 0 35880 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1649977179
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_408
timestamp 1649977179
transform 1 0 38640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_412
timestamp 1649977179
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_426
timestamp 1649977179
transform 1 0 40296 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1649977179
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1649977179
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_457
timestamp 1649977179
transform 1 0 43148 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_469
timestamp 1649977179
transform 1 0 44252 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6
timestamp 1649977179
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_18
timestamp 1649977179
transform 1 0 2760 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_30
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_42
timestamp 1649977179
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_60
timestamp 1649977179
transform 1 0 6624 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_72
timestamp 1649977179
transform 1 0 7728 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_84
timestamp 1649977179
transform 1 0 8832 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_96
timestamp 1649977179
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_131
timestamp 1649977179
transform 1 0 13156 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_143
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_155
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_177
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1649977179
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_209
timestamp 1649977179
transform 1 0 20332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_229
timestamp 1649977179
transform 1 0 22172 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1649977179
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_247
timestamp 1649977179
transform 1 0 23828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_259
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_271
timestamp 1649977179
transform 1 0 26036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1649977179
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_325
timestamp 1649977179
transform 1 0 31004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1649977179
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1649977179
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_349
timestamp 1649977179
transform 1 0 33212 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_359
timestamp 1649977179
transform 1 0 34132 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_364
timestamp 1649977179
transform 1 0 34592 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_376
timestamp 1649977179
transform 1 0 35696 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1649977179
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1649977179
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1649977179
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1649977179
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1649977179
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_449
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_457
timestamp 1649977179
transform 1 0 43148 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1649977179
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_468
timestamp 1649977179
transform 1 0 44160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_472
timestamp 1649977179
transform 1 0 44528 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6
timestamp 1649977179
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1649977179
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_116
timestamp 1649977179
transform 1 0 11776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_129
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1649977179
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_162
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1649977179
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_218
timestamp 1649977179
transform 1 0 21160 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_226
timestamp 1649977179
transform 1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_241
timestamp 1649977179
transform 1 0 23276 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1649977179
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_256
timestamp 1649977179
transform 1 0 24656 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_268
timestamp 1649977179
transform 1 0 25760 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_280
timestamp 1649977179
transform 1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_287
timestamp 1649977179
transform 1 0 27508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_291
timestamp 1649977179
transform 1 0 27876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1649977179
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1649977179
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_313
timestamp 1649977179
transform 1 0 29900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_320
timestamp 1649977179
transform 1 0 30544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_327
timestamp 1649977179
transform 1 0 31188 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_336
timestamp 1649977179
transform 1 0 32016 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_348
timestamp 1649977179
transform 1 0 33120 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1649977179
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1649977179
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_457
timestamp 1649977179
transform 1 0 43148 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_465
timestamp 1649977179
transform 1 0 43884 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_469
timestamp 1649977179
transform 1 0 44252 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_133
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_145
timestamp 1649977179
transform 1 0 14444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_157
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1649977179
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_173
timestamp 1649977179
transform 1 0 17020 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_180
timestamp 1649977179
transform 1 0 17664 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_191
timestamp 1649977179
transform 1 0 18676 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_198
timestamp 1649977179
transform 1 0 19320 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_210
timestamp 1649977179
transform 1 0 20424 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1649977179
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_248
timestamp 1649977179
transform 1 0 23920 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_255
timestamp 1649977179
transform 1 0 24564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_262
timestamp 1649977179
transform 1 0 25208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_270
timestamp 1649977179
transform 1 0 25944 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp 1649977179
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_304
timestamp 1649977179
transform 1 0 29072 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_308
timestamp 1649977179
transform 1 0 29440 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_315
timestamp 1649977179
transform 1 0 30084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_323
timestamp 1649977179
transform 1 0 30820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1649977179
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_357
timestamp 1649977179
transform 1 0 33948 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_369
timestamp 1649977179
transform 1 0 35052 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_381
timestamp 1649977179
transform 1 0 36156 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_389
timestamp 1649977179
transform 1 0 36892 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_103
timestamp 1649977179
transform 1 0 10580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_116
timestamp 1649977179
transform 1 0 11776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1649977179
transform 1 0 14352 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_164
timestamp 1649977179
transform 1 0 16192 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_176
timestamp 1649977179
transform 1 0 17296 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 1649977179
transform 1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_204
timestamp 1649977179
transform 1 0 19872 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_216
timestamp 1649977179
transform 1 0 20976 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_224
timestamp 1649977179
transform 1 0 21712 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_261
timestamp 1649977179
transform 1 0 25116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_268
timestamp 1649977179
transform 1 0 25760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1649977179
transform 1 0 26496 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_282
timestamp 1649977179
transform 1 0 27048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_291
timestamp 1649977179
transform 1 0 27876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_302
timestamp 1649977179
transform 1 0 28888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_329
timestamp 1649977179
transform 1 0 31372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_338
timestamp 1649977179
transform 1 0 32200 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_347
timestamp 1649977179
transform 1 0 33028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_356
timestamp 1649977179
transform 1 0 33856 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_13
timestamp 1649977179
transform 1 0 2300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_25
timestamp 1649977179
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_37
timestamp 1649977179
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1649977179
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_88
timestamp 1649977179
transform 1 0 9200 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1649977179
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_156
timestamp 1649977179
transform 1 0 15456 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_206
timestamp 1649977179
transform 1 0 20056 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1649977179
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_233
timestamp 1649977179
transform 1 0 22540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1649977179
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_253
timestamp 1649977179
transform 1 0 24380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_259
timestamp 1649977179
transform 1 0 24932 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_267
timestamp 1649977179
transform 1 0 25668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_285
timestamp 1649977179
transform 1 0 27324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_302
timestamp 1649977179
transform 1 0 28888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_316
timestamp 1649977179
transform 1 0 30176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_327
timestamp 1649977179
transform 1 0 31188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_342
timestamp 1649977179
transform 1 0 32568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_350
timestamp 1649977179
transform 1 0 33304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_372
timestamp 1649977179
transform 1 0 35328 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_379
timestamp 1649977179
transform 1 0 35972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_456
timestamp 1649977179
transform 1 0 43056 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_460
timestamp 1649977179
transform 1 0 43424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_472
timestamp 1649977179
transform 1 0 44528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_61
timestamp 1649977179
transform 1 0 6716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1649977179
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_88
timestamp 1649977179
transform 1 0 9200 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_149
timestamp 1649977179
transform 1 0 14812 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_160
timestamp 1649977179
transform 1 0 15824 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1649977179
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_204
timestamp 1649977179
transform 1 0 19872 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_216
timestamp 1649977179
transform 1 0 20976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_224
timestamp 1649977179
transform 1 0 21712 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_229
timestamp 1649977179
transform 1 0 22172 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_235
timestamp 1649977179
transform 1 0 22724 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_243
timestamp 1649977179
transform 1 0 23460 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_259
timestamp 1649977179
transform 1 0 24932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_271
timestamp 1649977179
transform 1 0 26036 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_276
timestamp 1649977179
transform 1 0 26496 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_283
timestamp 1649977179
transform 1 0 27140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_291
timestamp 1649977179
transform 1 0 27876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_316
timestamp 1649977179
transform 1 0 30176 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_324
timestamp 1649977179
transform 1 0 30912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_347
timestamp 1649977179
transform 1 0 33028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_354
timestamp 1649977179
transform 1 0 33672 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1649977179
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_368
timestamp 1649977179
transform 1 0 34960 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_375
timestamp 1649977179
transform 1 0 35604 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_382
timestamp 1649977179
transform 1 0 36248 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_394
timestamp 1649977179
transform 1 0 37352 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_406
timestamp 1649977179
transform 1 0 38456 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp 1649977179
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_73
timestamp 1649977179
transform 1 0 7820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_80
timestamp 1649977179
transform 1 0 8464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_84
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_88
timestamp 1649977179
transform 1 0 9200 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_116
timestamp 1649977179
transform 1 0 11776 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_120
timestamp 1649977179
transform 1 0 12144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_145
timestamp 1649977179
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1649977179
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1649977179
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_187
timestamp 1649977179
transform 1 0 18308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_199
timestamp 1649977179
transform 1 0 19412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_211
timestamp 1649977179
transform 1 0 20516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1649977179
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_241
timestamp 1649977179
transform 1 0 23276 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_252
timestamp 1649977179
transform 1 0 24288 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_264
timestamp 1649977179
transform 1 0 25392 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_272
timestamp 1649977179
transform 1 0 26128 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1649977179
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_302
timestamp 1649977179
transform 1 0 28888 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_308
timestamp 1649977179
transform 1 0 29440 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_319
timestamp 1649977179
transform 1 0 30452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1649977179
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_342
timestamp 1649977179
transform 1 0 32568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_366
timestamp 1649977179
transform 1 0 34776 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_380
timestamp 1649977179
transform 1 0 36064 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1649977179
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_91
timestamp 1649977179
transform 1 0 9476 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_100
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_104
timestamp 1649977179
transform 1 0 10672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1649977179
transform 1 0 16100 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_170
timestamp 1649977179
transform 1 0 16744 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_182
timestamp 1649977179
transform 1 0 17848 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_188
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_202
timestamp 1649977179
transform 1 0 19688 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_210
timestamp 1649977179
transform 1 0 20424 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_242
timestamp 1649977179
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1649977179
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_269
timestamp 1649977179
transform 1 0 25852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_297
timestamp 1649977179
transform 1 0 28428 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_305
timestamp 1649977179
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_332
timestamp 1649977179
transform 1 0 31648 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_339
timestamp 1649977179
transform 1 0 32292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 1649977179
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_426
timestamp 1649977179
transform 1 0 40296 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_438
timestamp 1649977179
transform 1 0 41400 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_450
timestamp 1649977179
transform 1 0 42504 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_462
timestamp 1649977179
transform 1 0 43608 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_470
timestamp 1649977179
transform 1 0 44344 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_6
timestamp 1649977179
transform 1 0 1656 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_14
timestamp 1649977179
transform 1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_36
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1649977179
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_124
timestamp 1649977179
transform 1 0 12512 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_132
timestamp 1649977179
transform 1 0 13248 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_180
timestamp 1649977179
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_200
timestamp 1649977179
transform 1 0 19504 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_238
timestamp 1649977179
transform 1 0 23000 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_245
timestamp 1649977179
transform 1 0 23644 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_252
timestamp 1649977179
transform 1 0 24288 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_263
timestamp 1649977179
transform 1 0 25300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1649977179
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_292
timestamp 1649977179
transform 1 0 27968 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_298
timestamp 1649977179
transform 1 0 28520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_319
timestamp 1649977179
transform 1 0 30452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_327
timestamp 1649977179
transform 1 0 31188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_341
timestamp 1649977179
transform 1 0 32476 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_367
timestamp 1649977179
transform 1 0 34868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_379
timestamp 1649977179
transform 1 0 35972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_413
timestamp 1649977179
transform 1 0 39100 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_417
timestamp 1649977179
transform 1 0 39468 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_427
timestamp 1649977179
transform 1 0 40388 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_437
timestamp 1649977179
transform 1 0 41308 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1649977179
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_47
timestamp 1649977179
transform 1 0 5428 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_55
timestamp 1649977179
transform 1 0 6164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 1649977179
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_101
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_108
timestamp 1649977179
transform 1 0 11040 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_116
timestamp 1649977179
transform 1 0 11776 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_171
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_178
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_186
timestamp 1649977179
transform 1 0 18216 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_213
timestamp 1649977179
transform 1 0 20700 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_226
timestamp 1649977179
transform 1 0 21896 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1649977179
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_271
timestamp 1649977179
transform 1 0 26036 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_291
timestamp 1649977179
transform 1 0 27876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1649977179
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_327
timestamp 1649977179
transform 1 0 31188 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_335
timestamp 1649977179
transform 1 0 31924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_353
timestamp 1649977179
transform 1 0 33580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1649977179
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_368
timestamp 1649977179
transform 1 0 34960 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_375
timestamp 1649977179
transform 1 0 35604 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_387
timestamp 1649977179
transform 1 0 36708 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_399
timestamp 1649977179
transform 1 0 37812 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_411
timestamp 1649977179
transform 1 0 38916 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1649977179
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_437
timestamp 1649977179
transform 1 0 41308 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_446
timestamp 1649977179
transform 1 0 42136 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_458
timestamp 1649977179
transform 1 0 43240 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_6
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_22
timestamp 1649977179
transform 1 0 3128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_42
timestamp 1649977179
transform 1 0 4968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_46
timestamp 1649977179
transform 1 0 5336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1649977179
transform 1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_66
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_77
timestamp 1649977179
transform 1 0 8188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_84
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_104
timestamp 1649977179
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_131
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_144
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_200
timestamp 1649977179
transform 1 0 19504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_213
timestamp 1649977179
transform 1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1649977179
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_245
timestamp 1649977179
transform 1 0 23644 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_253
timestamp 1649977179
transform 1 0 24380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_270
timestamp 1649977179
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1649977179
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_290
timestamp 1649977179
transform 1 0 27784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_298
timestamp 1649977179
transform 1 0 28520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_306
timestamp 1649977179
transform 1 0 29256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_310
timestamp 1649977179
transform 1 0 29624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_318
timestamp 1649977179
transform 1 0 30360 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_326
timestamp 1649977179
transform 1 0 31096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1649977179
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_343
timestamp 1649977179
transform 1 0 32660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_351
timestamp 1649977179
transform 1 0 33396 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_369
timestamp 1649977179
transform 1 0 35052 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_381
timestamp 1649977179
transform 1 0 36156 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp 1649977179
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_397
timestamp 1649977179
transform 1 0 37628 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_408
timestamp 1649977179
transform 1 0 38640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_428
timestamp 1649977179
transform 1 0 40480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_442
timestamp 1649977179
transform 1 0 41768 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_454
timestamp 1649977179
transform 1 0 42872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_465
timestamp 1649977179
transform 1 0 43884 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_469
timestamp 1649977179
transform 1 0 44252 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_52
timestamp 1649977179
transform 1 0 5888 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_76
timestamp 1649977179
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_119
timestamp 1649977179
transform 1 0 12052 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_150
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_174
timestamp 1649977179
transform 1 0 17112 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_186
timestamp 1649977179
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1649977179
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_219
timestamp 1649977179
transform 1 0 21252 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_227
timestamp 1649977179
transform 1 0 21988 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1649977179
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1649977179
transform 1 0 24840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_291
timestamp 1649977179
transform 1 0 27876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_299
timestamp 1649977179
transform 1 0 28612 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1649977179
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_314
timestamp 1649977179
transform 1 0 29992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_325
timestamp 1649977179
transform 1 0 31004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_335
timestamp 1649977179
transform 1 0 31924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_343
timestamp 1649977179
transform 1 0 32660 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1649977179
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_371
timestamp 1649977179
transform 1 0 35236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_383
timestamp 1649977179
transform 1 0 36340 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_391
timestamp 1649977179
transform 1 0 37076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_397
timestamp 1649977179
transform 1 0 37628 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_406
timestamp 1649977179
transform 1 0 38456 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_416
timestamp 1649977179
transform 1 0 39376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_427
timestamp 1649977179
transform 1 0 40388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_447
timestamp 1649977179
transform 1 0 42228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_456
timestamp 1649977179
transform 1 0 43056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_463
timestamp 1649977179
transform 1 0 43700 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_471
timestamp 1649977179
transform 1 0 44436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_24
timestamp 1649977179
transform 1 0 3312 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_44
timestamp 1649977179
transform 1 0 5152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_66
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_78
timestamp 1649977179
transform 1 0 8280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_85
timestamp 1649977179
transform 1 0 8924 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1649977179
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_122
timestamp 1649977179
transform 1 0 12328 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_128
timestamp 1649977179
transform 1 0 12880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_172
timestamp 1649977179
transform 1 0 16928 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_198
timestamp 1649977179
transform 1 0 19320 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_208
timestamp 1649977179
transform 1 0 20240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_235
timestamp 1649977179
transform 1 0 22724 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_241
timestamp 1649977179
transform 1 0 23276 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_262
timestamp 1649977179
transform 1 0 25208 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_270
timestamp 1649977179
transform 1 0 25944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1649977179
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_285
timestamp 1649977179
transform 1 0 27324 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_306
timestamp 1649977179
transform 1 0 29256 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_326
timestamp 1649977179
transform 1 0 31096 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1649977179
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_348
timestamp 1649977179
transform 1 0 33120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_371
timestamp 1649977179
transform 1 0 35236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_379
timestamp 1649977179
transform 1 0 35972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_386
timestamp 1649977179
transform 1 0 36616 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_401
timestamp 1649977179
transform 1 0 37996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_411
timestamp 1649977179
transform 1 0 38916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_425
timestamp 1649977179
transform 1 0 40204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_437
timestamp 1649977179
transform 1 0 41308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_444
timestamp 1649977179
transform 1 0 41952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_456
timestamp 1649977179
transform 1 0 43056 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_463
timestamp 1649977179
transform 1 0 43700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_471
timestamp 1649977179
transform 1 0 44436 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_74
timestamp 1649977179
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1649977179
transform 1 0 9200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_92
timestamp 1649977179
transform 1 0 9568 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_125
timestamp 1649977179
transform 1 0 12604 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_131
timestamp 1649977179
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_146
timestamp 1649977179
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_180
timestamp 1649977179
transform 1 0 17664 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_188
timestamp 1649977179
transform 1 0 18400 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_201
timestamp 1649977179
transform 1 0 19596 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_205
timestamp 1649977179
transform 1 0 19964 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_211
timestamp 1649977179
transform 1 0 20516 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1649977179
transform 1 0 22080 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_236
timestamp 1649977179
transform 1 0 22816 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_244
timestamp 1649977179
transform 1 0 23552 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1649977179
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_260
timestamp 1649977179
transform 1 0 25024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_268
timestamp 1649977179
transform 1 0 25760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_282
timestamp 1649977179
transform 1 0 27048 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_300
timestamp 1649977179
transform 1 0 28704 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_329
timestamp 1649977179
transform 1 0 31372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_353
timestamp 1649977179
transform 1 0 33580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 1649977179
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_370
timestamp 1649977179
transform 1 0 35144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_384
timestamp 1649977179
transform 1 0 36432 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_392
timestamp 1649977179
transform 1 0 37168 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_396
timestamp 1649977179
transform 1 0 37536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1649977179
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_429
timestamp 1649977179
transform 1 0 40572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_441
timestamp 1649977179
transform 1 0 41676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_451
timestamp 1649977179
transform 1 0 42596 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_460
timestamp 1649977179
transform 1 0 43424 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_472
timestamp 1649977179
transform 1 0 44528 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_7
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_11
timestamp 1649977179
transform 1 0 2116 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1649977179
transform 1 0 3312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_28
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1649977179
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1649977179
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_101
timestamp 1649977179
transform 1 0 10396 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_121
timestamp 1649977179
transform 1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_129
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_150
timestamp 1649977179
transform 1 0 14904 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_157
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_177
timestamp 1649977179
transform 1 0 17388 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_183
timestamp 1649977179
transform 1 0 17940 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_195
timestamp 1649977179
transform 1 0 19044 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_207
timestamp 1649977179
transform 1 0 20148 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_215
timestamp 1649977179
transform 1 0 20884 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1649977179
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_234
timestamp 1649977179
transform 1 0 22632 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_241
timestamp 1649977179
transform 1 0 23276 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_253
timestamp 1649977179
transform 1 0 24380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1649977179
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_319
timestamp 1649977179
transform 1 0 30452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_326
timestamp 1649977179
transform 1 0 31096 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1649977179
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_341
timestamp 1649977179
transform 1 0 32476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_348
timestamp 1649977179
transform 1 0 33120 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_354
timestamp 1649977179
transform 1 0 33672 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_375
timestamp 1649977179
transform 1 0 35604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_382
timestamp 1649977179
transform 1 0 36248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1649977179
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_398
timestamp 1649977179
transform 1 0 37720 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_407
timestamp 1649977179
transform 1 0 38548 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_421
timestamp 1649977179
transform 1 0 39836 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_436
timestamp 1649977179
transform 1 0 41216 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_443
timestamp 1649977179
transform 1 0 41860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_458
timestamp 1649977179
transform 1 0 43240 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_469
timestamp 1649977179
transform 1 0 44252 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_51
timestamp 1649977179
transform 1 0 5796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_73
timestamp 1649977179
transform 1 0 7820 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1649977179
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_101
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_114
timestamp 1649977179
transform 1 0 11592 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_118
timestamp 1649977179
transform 1 0 11960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_123
timestamp 1649977179
transform 1 0 12420 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_162
timestamp 1649977179
transform 1 0 16008 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_166
timestamp 1649977179
transform 1 0 16376 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_170
timestamp 1649977179
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_185
timestamp 1649977179
transform 1 0 18124 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_214
timestamp 1649977179
transform 1 0 20792 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_226
timestamp 1649977179
transform 1 0 21896 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_237
timestamp 1649977179
transform 1 0 22908 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1649977179
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_263
timestamp 1649977179
transform 1 0 25300 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_271
timestamp 1649977179
transform 1 0 26036 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_280
timestamp 1649977179
transform 1 0 26864 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_288
timestamp 1649977179
transform 1 0 27600 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_300
timestamp 1649977179
transform 1 0 28704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_313
timestamp 1649977179
transform 1 0 29900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_317
timestamp 1649977179
transform 1 0 30268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_326
timestamp 1649977179
transform 1 0 31096 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_334
timestamp 1649977179
transform 1 0 31832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_338
timestamp 1649977179
transform 1 0 32200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1649977179
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_375
timestamp 1649977179
transform 1 0 35604 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_383
timestamp 1649977179
transform 1 0 36340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_388
timestamp 1649977179
transform 1 0 36800 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_396
timestamp 1649977179
transform 1 0 37536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_416
timestamp 1649977179
transform 1 0 39376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_430
timestamp 1649977179
transform 1 0 40664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_440
timestamp 1649977179
transform 1 0 41584 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_447
timestamp 1649977179
transform 1 0 42228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_456
timestamp 1649977179
transform 1 0 43056 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_463
timestamp 1649977179
transform 1 0 43700 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_471
timestamp 1649977179
transform 1 0 44436 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_37
timestamp 1649977179
transform 1 0 4508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_62
timestamp 1649977179
transform 1 0 6808 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_76
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_135
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_141
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1649977179
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_176
timestamp 1649977179
transform 1 0 17296 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_202
timestamp 1649977179
transform 1 0 19688 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_212
timestamp 1649977179
transform 1 0 20608 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_216
timestamp 1649977179
transform 1 0 20976 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1649977179
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_229
timestamp 1649977179
transform 1 0 22172 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_236
timestamp 1649977179
transform 1 0 22816 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_243
timestamp 1649977179
transform 1 0 23460 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_252
timestamp 1649977179
transform 1 0 24288 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1649977179
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_284
timestamp 1649977179
transform 1 0 27232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_291
timestamp 1649977179
transform 1 0 27876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_298
timestamp 1649977179
transform 1 0 28520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_306
timestamp 1649977179
transform 1 0 29256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_314
timestamp 1649977179
transform 1 0 29992 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_320
timestamp 1649977179
transform 1 0 30544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_345
timestamp 1649977179
transform 1 0 32844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_352
timestamp 1649977179
transform 1 0 33488 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_359
timestamp 1649977179
transform 1 0 34132 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_367
timestamp 1649977179
transform 1 0 34868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_379
timestamp 1649977179
transform 1 0 35972 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_388
timestamp 1649977179
transform 1 0 36800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_399
timestamp 1649977179
transform 1 0 37812 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_407
timestamp 1649977179
transform 1 0 38548 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_419
timestamp 1649977179
transform 1 0 39652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_430
timestamp 1649977179
transform 1 0 40664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_440
timestamp 1649977179
transform 1 0 41584 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_459
timestamp 1649977179
transform 1 0 43332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_471
timestamp 1649977179
transform 1 0 44436 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_34
timestamp 1649977179
transform 1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_38
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_55
timestamp 1649977179
transform 1 0 6164 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_67
timestamp 1649977179
transform 1 0 7268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_75
timestamp 1649977179
transform 1 0 8004 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1649977179
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_99
timestamp 1649977179
transform 1 0 10212 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_144
timestamp 1649977179
transform 1 0 14352 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_148
timestamp 1649977179
transform 1 0 14720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_152
timestamp 1649977179
transform 1 0 15088 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_158
timestamp 1649977179
transform 1 0 15640 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_167
timestamp 1649977179
transform 1 0 16468 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_187
timestamp 1649977179
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_206
timestamp 1649977179
transform 1 0 20056 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_210
timestamp 1649977179
transform 1 0 20424 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_232
timestamp 1649977179
transform 1 0 22448 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1649977179
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1649977179
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1649977179
transform 1 0 24840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_268
timestamp 1649977179
transform 1 0 25760 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1649977179
transform 1 0 26312 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_284
timestamp 1649977179
transform 1 0 27232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_288
timestamp 1649977179
transform 1 0 27600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_292
timestamp 1649977179
transform 1 0 27968 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_298
timestamp 1649977179
transform 1 0 28520 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1649977179
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_315
timestamp 1649977179
transform 1 0 30084 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_323
timestamp 1649977179
transform 1 0 30820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_358
timestamp 1649977179
transform 1 0 34040 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_386
timestamp 1649977179
transform 1 0 36616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_406
timestamp 1649977179
transform 1 0 38456 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_416
timestamp 1649977179
transform 1 0 39376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_430
timestamp 1649977179
transform 1 0 40664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_450
timestamp 1649977179
transform 1 0 42504 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_19
timestamp 1649977179
transform 1 0 2852 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_23
timestamp 1649977179
transform 1 0 3220 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_35
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1649977179
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_87
timestamp 1649977179
transform 1 0 9108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_100
timestamp 1649977179
transform 1 0 10304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_121
timestamp 1649977179
transform 1 0 12236 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1649977179
transform 1 0 13064 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_139
timestamp 1649977179
transform 1 0 13892 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_190
timestamp 1649977179
transform 1 0 18584 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_209
timestamp 1649977179
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1649977179
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_235
timestamp 1649977179
transform 1 0 22724 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_243
timestamp 1649977179
transform 1 0 23460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_255
timestamp 1649977179
transform 1 0 24564 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_267
timestamp 1649977179
transform 1 0 25668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1649977179
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_301
timestamp 1649977179
transform 1 0 28796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_325
timestamp 1649977179
transform 1 0 31004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1649977179
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_353
timestamp 1649977179
transform 1 0 33580 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_366
timestamp 1649977179
transform 1 0 34776 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_379
timestamp 1649977179
transform 1 0 35972 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_409
timestamp 1649977179
transform 1 0 38732 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_413
timestamp 1649977179
transform 1 0 39100 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_419
timestamp 1649977179
transform 1 0 39652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_427
timestamp 1649977179
transform 1 0 40388 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_444
timestamp 1649977179
transform 1 0 41952 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_465
timestamp 1649977179
transform 1 0 43884 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_469
timestamp 1649977179
transform 1 0 44252 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_61
timestamp 1649977179
transform 1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1649977179
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_92
timestamp 1649977179
transform 1 0 9568 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_100
timestamp 1649977179
transform 1 0 10304 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_105
timestamp 1649977179
transform 1 0 10764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1649977179
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1649977179
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_144
timestamp 1649977179
transform 1 0 14352 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_148
timestamp 1649977179
transform 1 0 14720 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_157
timestamp 1649977179
transform 1 0 15548 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_168
timestamp 1649977179
transform 1 0 16560 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_176
timestamp 1649977179
transform 1 0 17296 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_184
timestamp 1649977179
transform 1 0 18032 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_188
timestamp 1649977179
transform 1 0 18400 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1649977179
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_200
timestamp 1649977179
transform 1 0 19504 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1649977179
transform 1 0 20608 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_217
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_241
timestamp 1649977179
transform 1 0 23276 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1649977179
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_271
timestamp 1649977179
transform 1 0 26036 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_275
timestamp 1649977179
transform 1 0 26404 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_299
timestamp 1649977179
transform 1 0 28612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_320
timestamp 1649977179
transform 1 0 30544 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_332
timestamp 1649977179
transform 1 0 31648 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1649977179
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_399
timestamp 1649977179
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_408
timestamp 1649977179
transform 1 0 38640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_412
timestamp 1649977179
transform 1 0 39008 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_416
timestamp 1649977179
transform 1 0 39376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_425
timestamp 1649977179
transform 1 0 40204 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_430
timestamp 1649977179
transform 1 0 40664 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_438
timestamp 1649977179
transform 1 0 41400 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_450
timestamp 1649977179
transform 1 0 42504 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_462
timestamp 1649977179
transform 1 0 43608 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_470
timestamp 1649977179
transform 1 0 44344 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_6
timestamp 1649977179
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1649977179
transform 1 0 2760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_25
timestamp 1649977179
transform 1 0 3404 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1649977179
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_65
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_84
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_95
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_122
timestamp 1649977179
transform 1 0 12328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_142
timestamp 1649977179
transform 1 0 14168 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1649977179
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_172
timestamp 1649977179
transform 1 0 16928 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_178
timestamp 1649977179
transform 1 0 17480 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_182
timestamp 1649977179
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_191
timestamp 1649977179
transform 1 0 18676 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_199
timestamp 1649977179
transform 1 0 19412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_208
timestamp 1649977179
transform 1 0 20240 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_216
timestamp 1649977179
transform 1 0 20976 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1649977179
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_243
timestamp 1649977179
transform 1 0 23460 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1649977179
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_263
timestamp 1649977179
transform 1 0 25300 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1649977179
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_359
timestamp 1649977179
transform 1 0 34132 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_371
timestamp 1649977179
transform 1 0 35236 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_383
timestamp 1649977179
transform 1 0 36340 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_71
timestamp 1649977179
transform 1 0 7636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1649977179
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_90
timestamp 1649977179
transform 1 0 9384 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_102
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_114
timestamp 1649977179
transform 1 0 11592 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_123
timestamp 1649977179
transform 1 0 12420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_172
timestamp 1649977179
transform 1 0 16928 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_205
timestamp 1649977179
transform 1 0 19964 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_214
timestamp 1649977179
transform 1 0 20792 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_222
timestamp 1649977179
transform 1 0 21528 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_227
timestamp 1649977179
transform 1 0 21988 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_231
timestamp 1649977179
transform 1 0 22356 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1649977179
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_456
timestamp 1649977179
transform 1 0 43056 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_464
timestamp 1649977179
transform 1 0 43792 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_86
timestamp 1649977179
transform 1 0 9016 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_98
timestamp 1649977179
transform 1 0 10120 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_124
timestamp 1649977179
transform 1 0 12512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1649977179
transform 1 0 13156 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_138
timestamp 1649977179
transform 1 0 13800 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_150
timestamp 1649977179
transform 1 0 14904 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1649977179
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_172
timestamp 1649977179
transform 1 0 16928 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_180
timestamp 1649977179
transform 1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_187
timestamp 1649977179
transform 1 0 18308 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_198
timestamp 1649977179
transform 1 0 19320 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_208
timestamp 1649977179
transform 1 0 20240 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1649977179
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_233
timestamp 1649977179
transform 1 0 22540 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_246
timestamp 1649977179
transform 1 0 23736 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_258
timestamp 1649977179
transform 1 0 24840 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_270
timestamp 1649977179
transform 1 0 25944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1649977179
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1649977179
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_185
timestamp 1649977179
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_201
timestamp 1649977179
transform 1 0 19596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_213
timestamp 1649977179
transform 1 0 20700 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_225
timestamp 1649977179
transform 1 0 21804 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_237
timestamp 1649977179
transform 1 0 22908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 1649977179
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_368
timestamp 1649977179
transform 1 0 34960 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_380
timestamp 1649977179
transform 1 0 36064 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_392
timestamp 1649977179
transform 1 0 37168 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_404
timestamp 1649977179
transform 1 0 38272 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_416
timestamp 1649977179
transform 1 0 39376 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_465
timestamp 1649977179
transform 1 0 43884 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_469
timestamp 1649977179
transform 1 0 44252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_11
timestamp 1649977179
transform 1 0 2116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1649977179
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_32
timestamp 1649977179
transform 1 0 4048 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_44
timestamp 1649977179
transform 1 0 5152 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_56
timestamp 1649977179
transform 1 0 6256 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_68
timestamp 1649977179
transform 1 0 7360 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_168
timestamp 1649977179
transform 1 0 16560 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_175
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 1649977179
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_424
timestamp 1649977179
transform 1 0 40112 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_436
timestamp 1649977179
transform 1 0 41216 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_448
timestamp 1649977179
transform 1 0 42320 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_456
timestamp 1649977179
transform 1 0 43056 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_461
timestamp 1649977179
transform 1 0 43516 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_468
timestamp 1649977179
transform 1 0 44160 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_472
timestamp 1649977179
transform 1 0 44528 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_23
timestamp 1649977179
transform 1 0 3220 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_29
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_34
timestamp 1649977179
transform 1 0 4232 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1649977179
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_62
timestamp 1649977179
transform 1 0 6808 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_70
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_76
timestamp 1649977179
transform 1 0 8096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_85
timestamp 1649977179
transform 1 0 8924 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1649977179
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_123
timestamp 1649977179
transform 1 0 12420 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_132
timestamp 1649977179
transform 1 0 13248 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_146
timestamp 1649977179
transform 1 0 14536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_158
timestamp 1649977179
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_173
timestamp 1649977179
transform 1 0 17020 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_177
timestamp 1649977179
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_182
timestamp 1649977179
transform 1 0 17848 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_194
timestamp 1649977179
transform 1 0 18952 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_197
timestamp 1649977179
transform 1 0 19228 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_202
timestamp 1649977179
transform 1 0 19688 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_210
timestamp 1649977179
transform 1 0 20424 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_233
timestamp 1649977179
transform 1 0 22540 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_256
timestamp 1649977179
transform 1 0 24656 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_268
timestamp 1649977179
transform 1 0 25760 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_272
timestamp 1649977179
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_289
timestamp 1649977179
transform 1 0 27692 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_312
timestamp 1649977179
transform 1 0 29808 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_324
timestamp 1649977179
transform 1 0 30912 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_328
timestamp 1649977179
transform 1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_368
timestamp 1649977179
transform 1 0 34960 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_377
timestamp 1649977179
transform 1 0 35788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1649977179
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_398
timestamp 1649977179
transform 1 0 37720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_406
timestamp 1649977179
transform 1 0 38456 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_413
timestamp 1649977179
transform 1 0 39100 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_419
timestamp 1649977179
transform 1 0 39652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_421
timestamp 1649977179
transform 1 0 39836 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_429
timestamp 1649977179
transform 1 0 40572 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_434
timestamp 1649977179
transform 1 0 41032 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1649977179
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_452
timestamp 1649977179
transform 1 0 42688 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_469
timestamp 1649977179
transform 1 0 44252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 44896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 44896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 44896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 44896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 44896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 44896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 44896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 44896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 44896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 44896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 44896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 44896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 44896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 44896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 44896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 44896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 44896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 44896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 44896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 44896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 44896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 44896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 44896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 44896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 44896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 44896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 44896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 44896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 19136 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 24288 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 29440 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 34592 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 39744 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _370_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _371_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _372_
timestamp 1649977179
transform 1 0 18032 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _373_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _374_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _375_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _376_
timestamp 1649977179
transform 1 0 21896 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _377_
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _378_
timestamp 1649977179
transform 1 0 22816 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _379_
timestamp 1649977179
transform 1 0 23644 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _380_
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _381_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24288 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _382_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _383_
timestamp 1649977179
transform 1 0 29256 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _384_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31004 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _385_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30544 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _386_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 28428 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _387_
timestamp 1649977179
transform 1 0 24656 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _388_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23920 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _389_
timestamp 1649977179
transform 1 0 24932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _390_
timestamp 1649977179
transform 1 0 23368 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _391_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _392_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _393_
timestamp 1649977179
transform 1 0 26036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _395_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25024 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _396_
timestamp 1649977179
transform 1 0 27416 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _397_
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _398_
timestamp 1649977179
transform 1 0 27232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _399_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _400_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _401_
timestamp 1649977179
transform 1 0 28612 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _402_
timestamp 1649977179
transform 1 0 30268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _403_
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _404_
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _405_
timestamp 1649977179
transform 1 0 33396 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _406_
timestamp 1649977179
transform 1 0 35972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _407_
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _408_
timestamp 1649977179
transform 1 0 30820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1649977179
transform 1 0 26220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _410_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _411_
timestamp 1649977179
transform 1 0 32568 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _412_
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _413_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27508 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _414_
timestamp 1649977179
transform 1 0 28244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _415_
timestamp 1649977179
transform 1 0 28428 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _416_
timestamp 1649977179
transform 1 0 26864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _417_
timestamp 1649977179
transform 1 0 33396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _418_
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _419_
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _420_
timestamp 1649977179
transform 1 0 35328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _421_
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1649977179
transform 1 0 17112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _423_
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _424_
timestamp 1649977179
transform 1 0 20240 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _425_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _426_
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _427_
timestamp 1649977179
transform 1 0 12788 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _428_
timestamp 1649977179
transform 1 0 12788 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _429_
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _430_
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _431_
timestamp 1649977179
transform 1 0 11592 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _432_
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _433_
timestamp 1649977179
transform 1 0 20516 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _434_
timestamp 1649977179
transform 1 0 19688 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _435_
timestamp 1649977179
transform 1 0 21896 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _436_
timestamp 1649977179
transform 1 0 20792 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _437_
timestamp 1649977179
transform 1 0 17480 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _438_
timestamp 1649977179
transform 1 0 17020 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _439_
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _440_
timestamp 1649977179
transform 1 0 17848 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 1649977179
transform 1 0 14536 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _443_
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _444_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15180 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _445_
timestamp 1649977179
transform 1 0 23000 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 1649977179
transform 1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _447_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _448_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14812 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _449_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _450_
timestamp 1649977179
transform 1 0 13432 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _451_
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _452_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _453_
timestamp 1649977179
transform 1 0 22816 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _454_
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _455_
timestamp 1649977179
transform 1 0 24840 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _456_
timestamp 1649977179
transform 1 0 23828 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _457_
timestamp 1649977179
transform 1 0 23092 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _458_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _459_
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _460_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26036 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _461_
timestamp 1649977179
transform 1 0 26404 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _462_
timestamp 1649977179
transform 1 0 26128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _463_
timestamp 1649977179
transform 1 0 23184 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _464_
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _465_
timestamp 1649977179
transform 1 0 38180 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 1649977179
transform 1 0 41952 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _467_
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _468_
timestamp 1649977179
transform 1 0 40020 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _469_
timestamp 1649977179
transform 1 0 36524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _470_
timestamp 1649977179
transform 1 0 43424 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _471_
timestamp 1649977179
transform 1 0 40848 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_1  _472_
timestamp 1649977179
transform 1 0 35604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _473_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _474_
timestamp 1649977179
transform 1 0 38088 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _475_
timestamp 1649977179
transform 1 0 32476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _476_
timestamp 1649977179
transform 1 0 29348 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _477_
timestamp 1649977179
transform 1 0 24748 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _478_
timestamp 1649977179
transform 1 0 29624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _479_
timestamp 1649977179
transform 1 0 28888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _480_
timestamp 1649977179
transform 1 0 28152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _481_
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _482_
timestamp 1649977179
transform 1 0 43240 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _483_
timestamp 1649977179
transform 1 0 37352 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _484_
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _485_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _486_
timestamp 1649977179
transform 1 0 41584 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _487_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _488_
timestamp 1649977179
transform 1 0 42596 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _489_
timestamp 1649977179
transform 1 0 43424 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _490_
timestamp 1649977179
transform 1 0 42964 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _491_
timestamp 1649977179
transform 1 0 43424 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _492_
timestamp 1649977179
transform 1 0 42596 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _493_
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _494_
timestamp 1649977179
transform 1 0 35972 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _495_
timestamp 1649977179
transform 1 0 37168 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _496_
timestamp 1649977179
transform 1 0 38916 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _497_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 41032 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _498_
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor4b_1  _499_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _500_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _501_
timestamp 1649977179
transform 1 0 26496 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _502_
timestamp 1649977179
transform 1 0 27232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _503_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26128 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _504_
timestamp 1649977179
transform 1 0 31464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _505_
timestamp 1649977179
transform 1 0 30636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _506_
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _507_
timestamp 1649977179
transform 1 0 36156 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _508_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _509_
timestamp 1649977179
transform 1 0 32568 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _510_
timestamp 1649977179
transform 1 0 9108 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _511_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _512_
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _513_
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _514_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10028 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _515_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _516_
timestamp 1649977179
transform 1 0 33304 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _517_
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _518_
timestamp 1649977179
transform 1 0 11776 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _520_
timestamp 1649977179
transform 1 0 10580 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _522_
timestamp 1649977179
transform 1 0 12696 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _523_
timestamp 1649977179
transform 1 0 42780 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _524_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _525_
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _526_
timestamp 1649977179
transform 1 0 12052 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _527_
timestamp 1649977179
transform 1 0 5428 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _528_
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _529_
timestamp 1649977179
transform 1 0 2852 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _530_
timestamp 1649977179
transform 1 0 3128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _531_
timestamp 1649977179
transform 1 0 33488 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _532_
timestamp 1649977179
transform 1 0 35144 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _533_
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _534_
timestamp 1649977179
transform 1 0 13524 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _535_
timestamp 1649977179
transform 1 0 15364 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _536_
timestamp 1649977179
transform 1 0 16928 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _537_
timestamp 1649977179
transform 1 0 33212 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _538_
timestamp 1649977179
transform 1 0 33948 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _539_
timestamp 1649977179
transform 1 0 2944 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _540_
timestamp 1649977179
transform 1 0 22080 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _541_
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _542_
timestamp 1649977179
transform 1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _543_
timestamp 1649977179
transform 1 0 23828 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _544_
timestamp 1649977179
transform 1 0 16468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _545_
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _546_
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _547_
timestamp 1649977179
transform 1 0 34500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _548_
timestamp 1649977179
transform 1 0 32200 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _549_
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _550_
timestamp 1649977179
transform 1 0 25208 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _551_
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _552_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _553_
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _554_
timestamp 1649977179
transform 1 0 28612 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _555_
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _556_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19688 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _557_
timestamp 1649977179
transform 1 0 19688 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _558_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _559_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _560_
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _561_
timestamp 1649977179
transform 1 0 25392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _562_
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _563_
timestamp 1649977179
transform 1 0 35512 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _564_
timestamp 1649977179
transform 1 0 30268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _565_
timestamp 1649977179
transform 1 0 27600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _566_
timestamp 1649977179
transform 1 0 33856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _567_
timestamp 1649977179
transform 1 0 25576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _568_
timestamp 1649977179
transform 1 0 27416 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _569_
timestamp 1649977179
transform 1 0 29992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _570_
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _571_
timestamp 1649977179
transform 1 0 32016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _572_
timestamp 1649977179
transform 1 0 24748 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _573_
timestamp 1649977179
transform 1 0 20976 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _574_
timestamp 1649977179
transform 1 0 17664 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _575_
timestamp 1649977179
transform 1 0 28428 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _576_
timestamp 1649977179
transform 1 0 30820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _577_
timestamp 1649977179
transform 1 0 28244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _578_
timestamp 1649977179
transform 1 0 27140 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _579_
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _580_
timestamp 1649977179
transform 1 0 25024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _581_
timestamp 1649977179
transform 1 0 28244 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _582_
timestamp 1649977179
transform 1 0 26220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _583_
timestamp 1649977179
transform 1 0 25668 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _584_
timestamp 1649977179
transform 1 0 25576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _585_
timestamp 1649977179
transform 1 0 21068 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _586_
timestamp 1649977179
transform 1 0 19872 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _587_
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _588_
timestamp 1649977179
transform 1 0 16836 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _589_
timestamp 1649977179
transform 1 0 12788 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _590_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _591_
timestamp 1649977179
transform 1 0 16008 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _592_
timestamp 1649977179
transform 1 0 11776 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _593_
timestamp 1649977179
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _594_
timestamp 1649977179
transform 1 0 12788 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _595_
timestamp 1649977179
transform 1 0 11684 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _596_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _597_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _598_
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _599_
timestamp 1649977179
transform 1 0 17204 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _600_
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _601_
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _602_
timestamp 1649977179
transform 1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _603_
timestamp 1649977179
transform 1 0 22540 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _604_
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _605_
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _606_
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _607_
timestamp 1649977179
transform 1 0 22448 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _608_
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _609_
timestamp 1649977179
transform 1 0 15272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _610__1
timestamp 1649977179
transform 1 0 15732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _611__2
timestamp 1649977179
transform 1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _612__3
timestamp 1649977179
transform 1 0 19044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _613_
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _614_
timestamp 1649977179
transform 1 0 19228 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _615_
timestamp 1649977179
transform 1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _616_
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _617_
timestamp 1649977179
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _618_
timestamp 1649977179
transform 1 0 22172 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _619_
timestamp 1649977179
transform 1 0 23368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _620_
timestamp 1649977179
transform 1 0 20700 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _621_
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _622_
timestamp 1649977179
transform 1 0 12788 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _623_
timestamp 1649977179
transform 1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _624_
timestamp 1649977179
transform 1 0 12144 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _625_
timestamp 1649977179
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _626_
timestamp 1649977179
transform 1 0 10948 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _627_
timestamp 1649977179
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _628_
timestamp 1649977179
transform 1 0 14720 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _629_
timestamp 1649977179
transform 1 0 15180 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _630_
timestamp 1649977179
transform 1 0 23000 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _631_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31372 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _632_
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _633_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30360 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _634_
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _635_
timestamp 1649977179
transform 1 0 36340 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _636_
timestamp 1649977179
transform 1 0 34684 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _637_
timestamp 1649977179
transform 1 0 39284 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__o2111a_1  _638_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32292 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _639_
timestamp 1649977179
transform 1 0 37352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _640_
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _641_
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _642_
timestamp 1649977179
transform 1 0 41676 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _643_
timestamp 1649977179
transform 1 0 39192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _644_
timestamp 1649977179
transform 1 0 39836 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _645_
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _646_
timestamp 1649977179
transform 1 0 42596 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _647_
timestamp 1649977179
transform 1 0 40020 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _648_
timestamp 1649977179
transform 1 0 40756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _649_
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _650_
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _651_
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _652_
timestamp 1649977179
transform 1 0 38272 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _653_
timestamp 1649977179
transform 1 0 38916 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _654_
timestamp 1649977179
transform 1 0 37260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _655_
timestamp 1649977179
transform 1 0 38824 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _656_
timestamp 1649977179
transform 1 0 36156 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _657_
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _658_
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _659_
timestamp 1649977179
transform 1 0 38180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _660_
timestamp 1649977179
transform 1 0 38824 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _661_
timestamp 1649977179
transform 1 0 37168 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _662_
timestamp 1649977179
transform 1 0 39192 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _663_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _664_
timestamp 1649977179
transform 1 0 40296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _665_
timestamp 1649977179
transform 1 0 41032 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _666_
timestamp 1649977179
transform 1 0 41032 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _667_
timestamp 1649977179
transform 1 0 40020 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _668_
timestamp 1649977179
transform 1 0 42872 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _669_
timestamp 1649977179
transform 1 0 31188 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _670_
timestamp 1649977179
transform 1 0 35328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _671_
timestamp 1649977179
transform 1 0 20608 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _672_
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _673_
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _674_
timestamp 1649977179
transform 1 0 25208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _675_
timestamp 1649977179
transform 1 0 7268 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _676_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _677_
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _678_
timestamp 1649977179
transform 1 0 9844 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _679_
timestamp 1649977179
transform 1 0 8188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _680_
timestamp 1649977179
transform 1 0 10580 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _681_
timestamp 1649977179
transform 1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _682_
timestamp 1649977179
transform 1 0 7636 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _683_
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _684_
timestamp 1649977179
transform 1 0 15364 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _685_
timestamp 1649977179
transform 1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _686_
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _687_
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _688_
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _689_
timestamp 1649977179
transform 1 0 6532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _690_
timestamp 1649977179
transform 1 0 6624 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _691_
timestamp 1649977179
transform 1 0 8648 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _692_
timestamp 1649977179
transform 1 0 9384 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _693_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _694_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _695_
timestamp 1649977179
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _696_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _697_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _698_
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _699_
timestamp 1649977179
transform 1 0 5520 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _700_
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _701_
timestamp 1649977179
transform 1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _702_
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _703_
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _704_
timestamp 1649977179
transform 1 0 21804 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _705_
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _706_
timestamp 1649977179
transform 1 0 25208 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _707_
timestamp 1649977179
transform 1 0 23828 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _708_
timestamp 1649977179
transform 1 0 13524 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _709_
timestamp 1649977179
transform 1 0 15732 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _710_
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _711_
timestamp 1649977179
transform 1 0 18308 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _712_
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _713_
timestamp 1649977179
transform 1 0 17848 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _714_
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _715_
timestamp 1649977179
transform 1 0 18216 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _716_
timestamp 1649977179
transform 1 0 17572 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _717_
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _718_
timestamp 1649977179
transform 1 0 19688 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _719_
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _720_
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _721_
timestamp 1649977179
transform 1 0 18676 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _722_
timestamp 1649977179
transform 1 0 19320 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _723_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19596 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _724_
timestamp 1649977179
transform 1 0 21712 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _725_
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _726_
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _727_
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _728_
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _729_
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _730_
timestamp 1649977179
transform 1 0 10212 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _731_
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _732_
timestamp 1649977179
transform 1 0 8004 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _733_
timestamp 1649977179
transform 1 0 11960 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _734_
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _735_
timestamp 1649977179
transform 1 0 11868 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _736_
timestamp 1649977179
transform 1 0 12236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _737_
timestamp 1649977179
transform 1 0 12880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _738_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12788 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _739_
timestamp 1649977179
transform 1 0 35788 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _740_
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _741_
timestamp 1649977179
transform 1 0 35144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _742_
timestamp 1649977179
transform 1 0 35696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _743_
timestamp 1649977179
transform 1 0 22172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _744_
timestamp 1649977179
transform 1 0 30912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _745_
timestamp 1649977179
transform 1 0 27968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _746_
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _747_
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _748_
timestamp 1649977179
transform 1 0 31280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _749_
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _750_
timestamp 1649977179
transform 1 0 30820 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _751_
timestamp 1649977179
transform 1 0 29716 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _752_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26772 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _753_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32292 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _754_
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _755_
timestamp 1649977179
transform 1 0 24656 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _756_
timestamp 1649977179
transform 1 0 31004 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _757_
timestamp 1649977179
transform 1 0 26036 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _758_
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _759_
timestamp 1649977179
transform 1 0 24472 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _760_
timestamp 1649977179
transform 1 0 29808 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _761_
timestamp 1649977179
transform 1 0 23368 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _762_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _763_
timestamp 1649977179
transform 1 0 27416 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _764_
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _765_
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _766_ shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26956 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _767_
timestamp 1649977179
transform 1 0 26404 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _768_
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _769_
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _770_
timestamp 1649977179
transform 1 0 11868 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _771_
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _772_
timestamp 1649977179
transform 1 0 14168 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _773_
timestamp 1649977179
transform 1 0 17848 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _774_
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _775_
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _776_
timestamp 1649977179
transform 1 0 20516 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _777_
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _778_
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _779_
timestamp 1649977179
transform 1 0 13064 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _780_
timestamp 1649977179
transform 1 0 14168 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _781__43 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16744 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _781_
timestamp 1649977179
transform 1 0 16376 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _782_
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _783_
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _784_
timestamp 1649977179
transform 1 0 32108 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _785_
timestamp 1649977179
transform 1 0 18032 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _786_
timestamp 1649977179
transform 1 0 22448 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _787_
timestamp 1649977179
transform 1 0 19872 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _788_
timestamp 1649977179
transform 1 0 6900 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _789_
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _790_
timestamp 1649977179
transform 1 0 6440 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _791_
timestamp 1649977179
transform 1 0 14536 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _792_
timestamp 1649977179
transform 1 0 17388 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _793_
timestamp 1649977179
transform 1 0 16928 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _794_
timestamp 1649977179
transform 1 0 21896 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _795_
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _796_
timestamp 1649977179
transform 1 0 12236 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _797_
timestamp 1649977179
transform 1 0 11868 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _798_
timestamp 1649977179
transform 1 0 12144 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _799_
timestamp 1649977179
transform 1 0 14720 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _800_
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _801_
timestamp 1649977179
transform 1 0 29624 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _802_
timestamp 1649977179
transform 1 0 32752 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _803_
timestamp 1649977179
transform 1 0 33580 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _804_
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _805_
timestamp 1649977179
transform 1 0 40756 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _806_
timestamp 1649977179
transform 1 0 39008 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _807_
timestamp 1649977179
transform 1 0 37904 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _808_
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _809_
timestamp 1649977179
transform 1 0 36984 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _810_
timestamp 1649977179
transform 1 0 37904 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _811_
timestamp 1649977179
transform 1 0 41032 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _812_
timestamp 1649977179
transform 1 0 40480 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _813_
timestamp 1649977179
transform 1 0 32752 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _814_
timestamp 1649977179
transform 1 0 14720 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _815_
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _816_
timestamp 1649977179
transform 1 0 20608 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _817_
timestamp 1649977179
transform 1 0 32660 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _818_
timestamp 1649977179
transform 1 0 24472 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _819_
timestamp 1649977179
transform 1 0 24564 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _820_
timestamp 1649977179
transform 1 0 18032 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _821_
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _822_
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _823_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _824_
timestamp 1649977179
transform 1 0 14628 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _825_
timestamp 1649977179
transform 1 0 3036 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _826_
timestamp 1649977179
transform 1 0 4324 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _827_
timestamp 1649977179
transform 1 0 6348 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _828_
timestamp 1649977179
transform 1 0 9660 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _829_
timestamp 1649977179
transform 1 0 9476 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _830_
timestamp 1649977179
transform 1 0 1840 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _831_
timestamp 1649977179
transform 1 0 3496 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _832_
timestamp 1649977179
transform 1 0 3680 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _833_
timestamp 1649977179
transform 1 0 3772 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _834_
timestamp 1649977179
transform 1 0 4692 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _835_
timestamp 1649977179
transform 1 0 9200 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _836_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _837_
timestamp 1649977179
transform 1 0 10580 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _838_
timestamp 1649977179
transform 1 0 4416 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _839_
timestamp 1649977179
transform 1 0 3956 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _840_
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _841_
timestamp 1649977179
transform 1 0 15272 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _842_
timestamp 1649977179
transform 1 0 17480 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _843_
timestamp 1649977179
transform 1 0 19412 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _844_
timestamp 1649977179
transform 1 0 19320 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _845_
timestamp 1649977179
transform 1 0 15456 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _846_
timestamp 1649977179
transform 1 0 17296 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _847_
timestamp 1649977179
transform 1 0 21988 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _848_
timestamp 1649977179
transform 1 0 22448 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _849_
timestamp 1649977179
transform 1 0 7360 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _850_
timestamp 1649977179
transform 1 0 6992 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _851_
timestamp 1649977179
transform 1 0 11776 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _852_
timestamp 1649977179
transform 1 0 12696 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _853_
timestamp 1649977179
transform 1 0 7728 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _854_
timestamp 1649977179
transform 1 0 3956 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _855_
timestamp 1649977179
transform 1 0 4416 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _856_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _857_
timestamp 1649977179
transform 1 0 33028 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _858_
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _859_
timestamp 1649977179
transform 1 0 32936 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _860_
timestamp 1649977179
transform 1 0 33396 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _861_
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _862_
timestamp 1649977179
transform 1 0 27232 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _863_
timestamp 1649977179
transform 1 0 21804 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _864_
timestamp 1649977179
transform 1 0 22080 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _865_
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _866_
timestamp 1649977179
transform 1 0 29716 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _906_
timestamp 1649977179
transform 1 0 42780 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22080 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_scan_clk_in
timestamp 1649977179
transform 1 0 6072 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_scan_clk_in
timestamp 1649977179
transform 1 0 2576 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_scan_clk_in
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1649977179
transform 1 0 28612 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1649977179
transform 1 0 31188 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1649977179
transform 1 0 28612 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1649977179
transform 1 0 33764 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7544 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1649977179
transform 1 0 6532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1649977179
transform 1 0 2392 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1649977179
transform 1 0 2576 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1649977179
transform 1 0 2576 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1649977179
transform 1 0 11500 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1649977179
transform 1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform 1 0 43884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 43240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 31004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 43976 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1649977179
transform 1 0 2116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1649977179
transform 1 0 3864 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1649977179
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform 1 0 32476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1649977179
transform 1 0 32292 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1649977179
transform 1 0 38732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform 1 0 43976 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform 1 0 24380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform 1 0 34684 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 9752 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1649977179
transform 1 0 43884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output28
timestamp 1649977179
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1649977179
transform 1 0 43884 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1649977179
transform 1 0 35512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1649977179
transform 1 0 17480 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1649977179
transform 1 0 43884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1649977179
transform 1 0 43884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1649977179
transform 1 0 40664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1649977179
transform 1 0 20700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform 1 0 43884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater42
timestamp 1649977179
transform 1 0 11868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  scan_controller_44
timestamp 1649977179
transform 1 0 12972 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_45
timestamp 1649977179
transform 1 0 15272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_46
timestamp 1649977179
transform 1 0 43976 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_47
timestamp 1649977179
transform 1 0 35512 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_48
timestamp 1649977179
transform 1 0 43240 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_49
timestamp 1649977179
transform 1 0 19412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_50
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_51
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_52
timestamp 1649977179
transform 1 0 43240 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_53
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_54
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_55
timestamp 1649977179
transform 1 0 43976 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_56
timestamp 1649977179
transform 1 0 43976 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_57
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_58
timestamp 1649977179
transform 1 0 37444 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_59
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_60
timestamp 1649977179
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_61
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_62
timestamp 1649977179
transform 1 0 43884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_63
timestamp 1649977179
transform 1 0 43976 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_64
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_65
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_66
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_67
timestamp 1649977179
transform 1 0 40020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_68
timestamp 1649977179
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_69
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_70
timestamp 1649977179
transform 1 0 14260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_71
timestamp 1649977179
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_72
timestamp 1649977179
transform 1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_73
timestamp 1649977179
transform 1 0 38732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_74
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_75
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_76
timestamp 1649977179
transform 1 0 22632 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_77
timestamp 1649977179
transform 1 0 29532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_78
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_79
timestamp 1649977179
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_80
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  scan_controller_81
timestamp 1649977179
transform 1 0 27784 0 -1 17408
box -38 -48 314 592
<< labels >>
flabel metal2 s 1278 19200 1390 20000 0 FreeSans 448 90 0 0 active_select[0]
port 0 nsew signal input
flabel metal2 s 43782 0 43894 800 0 FreeSans 448 90 0 0 active_select[1]
port 1 nsew signal input
flabel metal2 s 45070 0 45182 800 0 FreeSans 448 90 0 0 active_select[2]
port 2 nsew signal input
flabel metal2 s 36698 0 36810 800 0 FreeSans 448 90 0 0 active_select[3]
port 3 nsew signal input
flabel metal2 s 30902 19200 31014 20000 0 FreeSans 448 90 0 0 active_select[4]
port 4 nsew signal input
flabel metal2 s 25750 0 25862 800 0 FreeSans 448 90 0 0 active_select[5]
port 5 nsew signal input
flabel metal3 s 45200 7428 46000 7668 0 FreeSans 960 0 0 0 active_select[6]
port 6 nsew signal input
flabel metal3 s 0 16948 800 17188 0 FreeSans 960 0 0 0 active_select[7]
port 7 nsew signal input
flabel metal2 s 3210 19200 3322 20000 0 FreeSans 448 90 0 0 active_select[8]
port 8 nsew signal input
flabel metal2 s 33478 0 33590 800 0 FreeSans 448 90 0 0 clk
port 9 nsew signal input
flabel metal2 s 27038 0 27150 800 0 FreeSans 448 90 0 0 driver_sel[0]
port 10 nsew signal input
flabel metal2 s -10 19200 102 20000 0 FreeSans 448 90 0 0 driver_sel[1]
port 11 nsew signal input
flabel metal2 s 32190 0 32302 800 0 FreeSans 448 90 0 0 inputs[0]
port 12 nsew signal input
flabel metal2 s 10938 19200 11050 20000 0 FreeSans 448 90 0 0 inputs[1]
port 13 nsew signal input
flabel metal2 s 32190 19200 32302 20000 0 FreeSans 448 90 0 0 inputs[2]
port 14 nsew signal input
flabel metal2 s 38630 19200 38742 20000 0 FreeSans 448 90 0 0 inputs[3]
port 15 nsew signal input
flabel metal2 s 4498 19200 4610 20000 0 FreeSans 448 90 0 0 inputs[4]
port 16 nsew signal input
flabel metal2 s 12870 0 12982 800 0 FreeSans 448 90 0 0 inputs[5]
port 17 nsew signal input
flabel metal3 s 0 4708 800 4948 0 FreeSans 960 0 0 0 inputs[6]
port 18 nsew signal input
flabel metal2 s 41850 0 41962 800 0 FreeSans 448 90 0 0 inputs[7]
port 19 nsew signal input
flabel metal3 s 45200 8788 46000 9028 0 FreeSans 960 0 0 0 la_scan_clk_in
port 20 nsew signal input
flabel metal3 s 0 8108 800 8348 0 FreeSans 960 0 0 0 la_scan_data_in
port 21 nsew signal input
flabel metal3 s 45200 14228 46000 14468 0 FreeSans 960 0 0 0 la_scan_data_out
port 22 nsew signal tristate
flabel metal2 s 23818 19200 23930 20000 0 FreeSans 448 90 0 0 la_scan_latch_en
port 23 nsew signal input
flabel metal2 s 34122 19200 34234 20000 0 FreeSans 448 90 0 0 la_scan_select
port 24 nsew signal input
flabel metal2 s 12870 19200 12982 20000 0 FreeSans 448 90 0 0 oeb[0]
port 25 nsew signal tristate
flabel metal2 s 20598 0 20710 800 0 FreeSans 448 90 0 0 oeb[10]
port 26 nsew signal tristate
flabel metal3 s 45200 12188 46000 12428 0 FreeSans 960 0 0 0 oeb[11]
port 27 nsew signal tristate
flabel metal3 s 45200 15588 46000 15828 0 FreeSans 960 0 0 0 oeb[12]
port 28 nsew signal tristate
flabel metal2 s 28970 0 29082 800 0 FreeSans 448 90 0 0 oeb[13]
port 29 nsew signal tristate
flabel metal2 s 37342 19200 37454 20000 0 FreeSans 448 90 0 0 oeb[14]
port 30 nsew signal tristate
flabel metal2 s 3210 0 3322 800 0 FreeSans 448 90 0 0 oeb[15]
port 31 nsew signal tristate
flabel metal2 s 7718 19200 7830 20000 0 FreeSans 448 90 0 0 oeb[16]
port 32 nsew signal tristate
flabel metal2 s 10938 0 11050 800 0 FreeSans 448 90 0 0 oeb[17]
port 33 nsew signal tristate
flabel metal2 s 43782 19200 43894 20000 0 FreeSans 448 90 0 0 oeb[18]
port 34 nsew signal tristate
flabel metal3 s 45200 10828 46000 11068 0 FreeSans 960 0 0 0 oeb[19]
port 35 nsew signal tristate
flabel metal2 s 16090 0 16202 800 0 FreeSans 448 90 0 0 oeb[1]
port 36 nsew signal tristate
flabel metal2 s 41850 19200 41962 20000 0 FreeSans 448 90 0 0 oeb[20]
port 37 nsew signal tristate
flabel metal2 s 7718 0 7830 800 0 FreeSans 448 90 0 0 oeb[21]
port 38 nsew signal tristate
flabel metal2 s 23818 0 23930 800 0 FreeSans 448 90 0 0 oeb[22]
port 39 nsew signal tristate
flabel metal2 s 39918 0 40030 800 0 FreeSans 448 90 0 0 oeb[23]
port 40 nsew signal tristate
flabel metal2 s 6430 19200 6542 20000 0 FreeSans 448 90 0 0 oeb[24]
port 41 nsew signal tristate
flabel metal2 s 19310 0 19422 800 0 FreeSans 448 90 0 0 oeb[25]
port 42 nsew signal tristate
flabel metal2 s 14158 19200 14270 20000 0 FreeSans 448 90 0 0 oeb[26]
port 43 nsew signal tristate
flabel metal2 s 30258 0 30370 800 0 FreeSans 448 90 0 0 oeb[27]
port 44 nsew signal tristate
flabel metal2 s 25750 19200 25862 20000 0 FreeSans 448 90 0 0 oeb[28]
port 45 nsew signal tristate
flabel metal2 s 38630 0 38742 800 0 FreeSans 448 90 0 0 oeb[29]
port 46 nsew signal tristate
flabel metal3 s 45200 628 46000 868 0 FreeSans 960 0 0 0 oeb[2]
port 47 nsew signal tristate
flabel metal3 s 0 6748 800 6988 0 FreeSans 960 0 0 0 oeb[30]
port 48 nsew signal tristate
flabel metal3 s 0 1308 800 1548 0 FreeSans 960 0 0 0 oeb[31]
port 49 nsew signal tristate
flabel metal2 s 22530 19200 22642 20000 0 FreeSans 448 90 0 0 oeb[32]
port 50 nsew signal tristate
flabel metal2 s 28970 19200 29082 20000 0 FreeSans 448 90 0 0 oeb[33]
port 51 nsew signal tristate
flabel metal3 s 0 3348 800 3588 0 FreeSans 960 0 0 0 oeb[34]
port 52 nsew signal tristate
flabel metal2 s -10 0 102 800 0 FreeSans 448 90 0 0 oeb[35]
port 53 nsew signal tristate
flabel metal3 s 0 18308 800 18548 0 FreeSans 960 0 0 0 oeb[36]
port 54 nsew signal tristate
flabel metal2 s 27682 19200 27794 20000 0 FreeSans 448 90 0 0 oeb[37]
port 55 nsew signal tristate
flabel metal2 s 35410 19200 35522 20000 0 FreeSans 448 90 0 0 oeb[3]
port 56 nsew signal tristate
flabel metal2 s 45070 19200 45182 20000 0 FreeSans 448 90 0 0 oeb[4]
port 57 nsew signal tristate
flabel metal2 s 19310 19200 19422 20000 0 FreeSans 448 90 0 0 oeb[5]
port 58 nsew signal tristate
flabel metal2 s 4498 0 4610 800 0 FreeSans 448 90 0 0 oeb[6]
port 59 nsew signal tristate
flabel metal2 s 1278 0 1390 800 0 FreeSans 448 90 0 0 oeb[7]
port 60 nsew signal tristate
flabel metal3 s 45200 18988 46000 19228 0 FreeSans 960 0 0 0 oeb[8]
port 61 nsew signal tristate
flabel metal3 s 0 13548 800 13788 0 FreeSans 960 0 0 0 oeb[9]
port 62 nsew signal tristate
flabel metal2 s 14158 0 14270 800 0 FreeSans 448 90 0 0 outputs[0]
port 63 nsew signal tristate
flabel metal3 s 45200 17628 46000 17868 0 FreeSans 960 0 0 0 outputs[1]
port 64 nsew signal tristate
flabel metal2 s 35410 0 35522 800 0 FreeSans 448 90 0 0 outputs[2]
port 65 nsew signal tristate
flabel metal2 s 17378 19200 17490 20000 0 FreeSans 448 90 0 0 outputs[3]
port 66 nsew signal tristate
flabel metal3 s 45200 4028 46000 4268 0 FreeSans 960 0 0 0 outputs[4]
port 67 nsew signal tristate
flabel metal2 s 6430 0 6542 800 0 FreeSans 448 90 0 0 outputs[5]
port 68 nsew signal tristate
flabel metal2 s 9650 0 9762 800 0 FreeSans 448 90 0 0 outputs[6]
port 69 nsew signal tristate
flabel metal3 s 0 14908 800 15148 0 FreeSans 960 0 0 0 outputs[7]
port 70 nsew signal tristate
flabel metal3 s 45200 5388 46000 5628 0 FreeSans 960 0 0 0 ready
port 71 nsew signal tristate
flabel metal2 s 17378 0 17490 800 0 FreeSans 448 90 0 0 reset
port 72 nsew signal input
flabel metal3 s 0 11508 800 11748 0 FreeSans 960 0 0 0 scan_clk_in
port 73 nsew signal input
flabel metal2 s 40562 19200 40674 20000 0 FreeSans 448 90 0 0 scan_clk_out
port 74 nsew signal tristate
flabel metal2 s 16090 19200 16202 20000 0 FreeSans 448 90 0 0 scan_data_in
port 75 nsew signal input
flabel metal2 s 20598 19200 20710 20000 0 FreeSans 448 90 0 0 scan_data_out
port 76 nsew signal tristate
flabel metal2 s 22530 0 22642 800 0 FreeSans 448 90 0 0 scan_latch_en
port 77 nsew signal tristate
flabel metal3 s 0 10148 800 10388 0 FreeSans 960 0 0 0 scan_select
port 78 nsew signal tristate
flabel metal2 s 9650 19200 9762 20000 0 FreeSans 448 90 0 0 set_clk_div
port 79 nsew signal input
flabel metal3 s 45200 1988 46000 2228 0 FreeSans 960 0 0 0 slow_clk
port 80 nsew signal tristate
flabel metal4 s 6418 2128 6738 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 17366 2128 17686 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 28314 2128 28634 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 39262 2128 39582 17456 0 FreeSans 1920 90 0 0 vccd1
port 81 nsew power bidirectional
flabel metal4 s 11892 2128 12212 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
flabel metal4 s 22840 2128 23160 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
flabel metal4 s 33788 2128 34108 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
flabel metal4 s 44736 2128 45056 17456 0 FreeSans 1920 90 0 0 vssd1
port 82 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 46000 20000
<< end >>
