module user_project_wrapper (user_clock2,
    vccd1,
    vccd2,
    vdda1,
    vdda2,
    vssa1,
    vssa2,
    vssd1,
    vssd2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input vccd1;
 input vccd2;
 input vdda1;
 input vdda2;
 input vssa1;
 input vssa2;
 input vssd1;
 input vssd2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire sc_clk_in;
 wire sc_clk_out;
 wire sc_data_in;
 wire sc_data_out;
 wire sc_latch_out;
 wire sc_scan_out;
 wire sw_000_clk_out;
 wire sw_000_data_out;
 wire sw_000_latch_out;
 wire \sw_000_module_data_in[0] ;
 wire \sw_000_module_data_in[1] ;
 wire \sw_000_module_data_in[2] ;
 wire \sw_000_module_data_in[3] ;
 wire \sw_000_module_data_in[4] ;
 wire \sw_000_module_data_in[5] ;
 wire \sw_000_module_data_in[6] ;
 wire \sw_000_module_data_in[7] ;
 wire \sw_000_module_data_out[0] ;
 wire \sw_000_module_data_out[1] ;
 wire \sw_000_module_data_out[2] ;
 wire \sw_000_module_data_out[3] ;
 wire \sw_000_module_data_out[4] ;
 wire \sw_000_module_data_out[5] ;
 wire \sw_000_module_data_out[6] ;
 wire \sw_000_module_data_out[7] ;
 wire sw_000_scan_out;
 wire sw_001_clk_out;
 wire sw_001_data_out;
 wire sw_001_latch_out;
 wire \sw_001_module_data_in[0] ;
 wire \sw_001_module_data_in[1] ;
 wire \sw_001_module_data_in[2] ;
 wire \sw_001_module_data_in[3] ;
 wire \sw_001_module_data_in[4] ;
 wire \sw_001_module_data_in[5] ;
 wire \sw_001_module_data_in[6] ;
 wire \sw_001_module_data_in[7] ;
 wire \sw_001_module_data_out[0] ;
 wire \sw_001_module_data_out[1] ;
 wire \sw_001_module_data_out[2] ;
 wire \sw_001_module_data_out[3] ;
 wire \sw_001_module_data_out[4] ;
 wire \sw_001_module_data_out[5] ;
 wire \sw_001_module_data_out[6] ;
 wire \sw_001_module_data_out[7] ;
 wire sw_001_scan_out;
 wire sw_002_clk_out;
 wire sw_002_data_out;
 wire sw_002_latch_out;
 wire \sw_002_module_data_in[0] ;
 wire \sw_002_module_data_in[1] ;
 wire \sw_002_module_data_in[2] ;
 wire \sw_002_module_data_in[3] ;
 wire \sw_002_module_data_in[4] ;
 wire \sw_002_module_data_in[5] ;
 wire \sw_002_module_data_in[6] ;
 wire \sw_002_module_data_in[7] ;
 wire \sw_002_module_data_out[0] ;
 wire \sw_002_module_data_out[1] ;
 wire \sw_002_module_data_out[2] ;
 wire \sw_002_module_data_out[3] ;
 wire \sw_002_module_data_out[4] ;
 wire \sw_002_module_data_out[5] ;
 wire \sw_002_module_data_out[6] ;
 wire \sw_002_module_data_out[7] ;
 wire sw_002_scan_out;
 wire sw_003_clk_out;
 wire sw_003_data_out;
 wire sw_003_latch_out;
 wire \sw_003_module_data_in[0] ;
 wire \sw_003_module_data_in[1] ;
 wire \sw_003_module_data_in[2] ;
 wire \sw_003_module_data_in[3] ;
 wire \sw_003_module_data_in[4] ;
 wire \sw_003_module_data_in[5] ;
 wire \sw_003_module_data_in[6] ;
 wire \sw_003_module_data_in[7] ;
 wire \sw_003_module_data_out[0] ;
 wire \sw_003_module_data_out[1] ;
 wire \sw_003_module_data_out[2] ;
 wire \sw_003_module_data_out[3] ;
 wire \sw_003_module_data_out[4] ;
 wire \sw_003_module_data_out[5] ;
 wire \sw_003_module_data_out[6] ;
 wire \sw_003_module_data_out[7] ;
 wire sw_003_scan_out;
 wire sw_004_clk_out;
 wire sw_004_data_out;
 wire sw_004_latch_out;
 wire \sw_004_module_data_in[0] ;
 wire \sw_004_module_data_in[1] ;
 wire \sw_004_module_data_in[2] ;
 wire \sw_004_module_data_in[3] ;
 wire \sw_004_module_data_in[4] ;
 wire \sw_004_module_data_in[5] ;
 wire \sw_004_module_data_in[6] ;
 wire \sw_004_module_data_in[7] ;
 wire \sw_004_module_data_out[0] ;
 wire \sw_004_module_data_out[1] ;
 wire \sw_004_module_data_out[2] ;
 wire \sw_004_module_data_out[3] ;
 wire \sw_004_module_data_out[4] ;
 wire \sw_004_module_data_out[5] ;
 wire \sw_004_module_data_out[6] ;
 wire \sw_004_module_data_out[7] ;
 wire sw_004_scan_out;
 wire sw_005_clk_out;
 wire sw_005_data_out;
 wire sw_005_latch_out;
 wire \sw_005_module_data_in[0] ;
 wire \sw_005_module_data_in[1] ;
 wire \sw_005_module_data_in[2] ;
 wire \sw_005_module_data_in[3] ;
 wire \sw_005_module_data_in[4] ;
 wire \sw_005_module_data_in[5] ;
 wire \sw_005_module_data_in[6] ;
 wire \sw_005_module_data_in[7] ;
 wire \sw_005_module_data_out[0] ;
 wire \sw_005_module_data_out[1] ;
 wire \sw_005_module_data_out[2] ;
 wire \sw_005_module_data_out[3] ;
 wire \sw_005_module_data_out[4] ;
 wire \sw_005_module_data_out[5] ;
 wire \sw_005_module_data_out[6] ;
 wire \sw_005_module_data_out[7] ;
 wire sw_005_scan_out;
 wire sw_006_clk_out;
 wire sw_006_data_out;
 wire sw_006_latch_out;
 wire \sw_006_module_data_in[0] ;
 wire \sw_006_module_data_in[1] ;
 wire \sw_006_module_data_in[2] ;
 wire \sw_006_module_data_in[3] ;
 wire \sw_006_module_data_in[4] ;
 wire \sw_006_module_data_in[5] ;
 wire \sw_006_module_data_in[6] ;
 wire \sw_006_module_data_in[7] ;
 wire \sw_006_module_data_out[0] ;
 wire \sw_006_module_data_out[1] ;
 wire \sw_006_module_data_out[2] ;
 wire \sw_006_module_data_out[3] ;
 wire \sw_006_module_data_out[4] ;
 wire \sw_006_module_data_out[5] ;
 wire \sw_006_module_data_out[6] ;
 wire \sw_006_module_data_out[7] ;
 wire sw_006_scan_out;
 wire sw_007_clk_out;
 wire sw_007_data_out;
 wire sw_007_latch_out;
 wire \sw_007_module_data_in[0] ;
 wire \sw_007_module_data_in[1] ;
 wire \sw_007_module_data_in[2] ;
 wire \sw_007_module_data_in[3] ;
 wire \sw_007_module_data_in[4] ;
 wire \sw_007_module_data_in[5] ;
 wire \sw_007_module_data_in[6] ;
 wire \sw_007_module_data_in[7] ;
 wire \sw_007_module_data_out[0] ;
 wire \sw_007_module_data_out[1] ;
 wire \sw_007_module_data_out[2] ;
 wire \sw_007_module_data_out[3] ;
 wire \sw_007_module_data_out[4] ;
 wire \sw_007_module_data_out[5] ;
 wire \sw_007_module_data_out[6] ;
 wire \sw_007_module_data_out[7] ;
 wire sw_007_scan_out;
 wire sw_008_clk_out;
 wire sw_008_data_out;
 wire sw_008_latch_out;
 wire \sw_008_module_data_in[0] ;
 wire \sw_008_module_data_in[1] ;
 wire \sw_008_module_data_in[2] ;
 wire \sw_008_module_data_in[3] ;
 wire \sw_008_module_data_in[4] ;
 wire \sw_008_module_data_in[5] ;
 wire \sw_008_module_data_in[6] ;
 wire \sw_008_module_data_in[7] ;
 wire \sw_008_module_data_out[0] ;
 wire \sw_008_module_data_out[1] ;
 wire \sw_008_module_data_out[2] ;
 wire \sw_008_module_data_out[3] ;
 wire \sw_008_module_data_out[4] ;
 wire \sw_008_module_data_out[5] ;
 wire \sw_008_module_data_out[6] ;
 wire \sw_008_module_data_out[7] ;
 wire sw_008_scan_out;
 wire sw_009_clk_out;
 wire sw_009_data_out;
 wire sw_009_latch_out;
 wire \sw_009_module_data_in[0] ;
 wire \sw_009_module_data_in[1] ;
 wire \sw_009_module_data_in[2] ;
 wire \sw_009_module_data_in[3] ;
 wire \sw_009_module_data_in[4] ;
 wire \sw_009_module_data_in[5] ;
 wire \sw_009_module_data_in[6] ;
 wire \sw_009_module_data_in[7] ;
 wire \sw_009_module_data_out[0] ;
 wire \sw_009_module_data_out[1] ;
 wire \sw_009_module_data_out[2] ;
 wire \sw_009_module_data_out[3] ;
 wire \sw_009_module_data_out[4] ;
 wire \sw_009_module_data_out[5] ;
 wire \sw_009_module_data_out[6] ;
 wire \sw_009_module_data_out[7] ;
 wire sw_009_scan_out;
 wire sw_010_clk_out;
 wire sw_010_data_out;
 wire sw_010_latch_out;
 wire \sw_010_module_data_in[0] ;
 wire \sw_010_module_data_in[1] ;
 wire \sw_010_module_data_in[2] ;
 wire \sw_010_module_data_in[3] ;
 wire \sw_010_module_data_in[4] ;
 wire \sw_010_module_data_in[5] ;
 wire \sw_010_module_data_in[6] ;
 wire \sw_010_module_data_in[7] ;
 wire \sw_010_module_data_out[0] ;
 wire \sw_010_module_data_out[1] ;
 wire \sw_010_module_data_out[2] ;
 wire \sw_010_module_data_out[3] ;
 wire \sw_010_module_data_out[4] ;
 wire \sw_010_module_data_out[5] ;
 wire \sw_010_module_data_out[6] ;
 wire \sw_010_module_data_out[7] ;
 wire sw_010_scan_out;
 wire sw_011_clk_out;
 wire sw_011_data_out;
 wire sw_011_latch_out;
 wire \sw_011_module_data_in[0] ;
 wire \sw_011_module_data_in[1] ;
 wire \sw_011_module_data_in[2] ;
 wire \sw_011_module_data_in[3] ;
 wire \sw_011_module_data_in[4] ;
 wire \sw_011_module_data_in[5] ;
 wire \sw_011_module_data_in[6] ;
 wire \sw_011_module_data_in[7] ;
 wire \sw_011_module_data_out[0] ;
 wire \sw_011_module_data_out[1] ;
 wire \sw_011_module_data_out[2] ;
 wire \sw_011_module_data_out[3] ;
 wire \sw_011_module_data_out[4] ;
 wire \sw_011_module_data_out[5] ;
 wire \sw_011_module_data_out[6] ;
 wire \sw_011_module_data_out[7] ;
 wire sw_011_scan_out;
 wire sw_012_clk_out;
 wire sw_012_data_out;
 wire sw_012_latch_out;
 wire \sw_012_module_data_in[0] ;
 wire \sw_012_module_data_in[1] ;
 wire \sw_012_module_data_in[2] ;
 wire \sw_012_module_data_in[3] ;
 wire \sw_012_module_data_in[4] ;
 wire \sw_012_module_data_in[5] ;
 wire \sw_012_module_data_in[6] ;
 wire \sw_012_module_data_in[7] ;
 wire \sw_012_module_data_out[0] ;
 wire \sw_012_module_data_out[1] ;
 wire \sw_012_module_data_out[2] ;
 wire \sw_012_module_data_out[3] ;
 wire \sw_012_module_data_out[4] ;
 wire \sw_012_module_data_out[5] ;
 wire \sw_012_module_data_out[6] ;
 wire \sw_012_module_data_out[7] ;
 wire sw_012_scan_out;
 wire sw_013_clk_out;
 wire sw_013_data_out;
 wire sw_013_latch_out;
 wire \sw_013_module_data_in[0] ;
 wire \sw_013_module_data_in[1] ;
 wire \sw_013_module_data_in[2] ;
 wire \sw_013_module_data_in[3] ;
 wire \sw_013_module_data_in[4] ;
 wire \sw_013_module_data_in[5] ;
 wire \sw_013_module_data_in[6] ;
 wire \sw_013_module_data_in[7] ;
 wire \sw_013_module_data_out[0] ;
 wire \sw_013_module_data_out[1] ;
 wire \sw_013_module_data_out[2] ;
 wire \sw_013_module_data_out[3] ;
 wire \sw_013_module_data_out[4] ;
 wire \sw_013_module_data_out[5] ;
 wire \sw_013_module_data_out[6] ;
 wire \sw_013_module_data_out[7] ;
 wire sw_013_scan_out;
 wire sw_014_clk_out;
 wire sw_014_data_out;
 wire sw_014_latch_out;
 wire \sw_014_module_data_in[0] ;
 wire \sw_014_module_data_in[1] ;
 wire \sw_014_module_data_in[2] ;
 wire \sw_014_module_data_in[3] ;
 wire \sw_014_module_data_in[4] ;
 wire \sw_014_module_data_in[5] ;
 wire \sw_014_module_data_in[6] ;
 wire \sw_014_module_data_in[7] ;
 wire \sw_014_module_data_out[0] ;
 wire \sw_014_module_data_out[1] ;
 wire \sw_014_module_data_out[2] ;
 wire \sw_014_module_data_out[3] ;
 wire \sw_014_module_data_out[4] ;
 wire \sw_014_module_data_out[5] ;
 wire \sw_014_module_data_out[6] ;
 wire \sw_014_module_data_out[7] ;
 wire sw_014_scan_out;
 wire sw_015_clk_out;
 wire sw_015_data_out;
 wire sw_015_latch_out;
 wire \sw_015_module_data_in[0] ;
 wire \sw_015_module_data_in[1] ;
 wire \sw_015_module_data_in[2] ;
 wire \sw_015_module_data_in[3] ;
 wire \sw_015_module_data_in[4] ;
 wire \sw_015_module_data_in[5] ;
 wire \sw_015_module_data_in[6] ;
 wire \sw_015_module_data_in[7] ;
 wire \sw_015_module_data_out[0] ;
 wire \sw_015_module_data_out[1] ;
 wire \sw_015_module_data_out[2] ;
 wire \sw_015_module_data_out[3] ;
 wire \sw_015_module_data_out[4] ;
 wire \sw_015_module_data_out[5] ;
 wire \sw_015_module_data_out[6] ;
 wire \sw_015_module_data_out[7] ;
 wire sw_015_scan_out;
 wire sw_016_clk_out;
 wire sw_016_data_out;
 wire sw_016_latch_out;
 wire \sw_016_module_data_in[0] ;
 wire \sw_016_module_data_in[1] ;
 wire \sw_016_module_data_in[2] ;
 wire \sw_016_module_data_in[3] ;
 wire \sw_016_module_data_in[4] ;
 wire \sw_016_module_data_in[5] ;
 wire \sw_016_module_data_in[6] ;
 wire \sw_016_module_data_in[7] ;
 wire \sw_016_module_data_out[0] ;
 wire \sw_016_module_data_out[1] ;
 wire \sw_016_module_data_out[2] ;
 wire \sw_016_module_data_out[3] ;
 wire \sw_016_module_data_out[4] ;
 wire \sw_016_module_data_out[5] ;
 wire \sw_016_module_data_out[6] ;
 wire \sw_016_module_data_out[7] ;
 wire sw_016_scan_out;
 wire sw_017_clk_out;
 wire sw_017_data_out;
 wire sw_017_latch_out;
 wire \sw_017_module_data_in[0] ;
 wire \sw_017_module_data_in[1] ;
 wire \sw_017_module_data_in[2] ;
 wire \sw_017_module_data_in[3] ;
 wire \sw_017_module_data_in[4] ;
 wire \sw_017_module_data_in[5] ;
 wire \sw_017_module_data_in[6] ;
 wire \sw_017_module_data_in[7] ;
 wire \sw_017_module_data_out[0] ;
 wire \sw_017_module_data_out[1] ;
 wire \sw_017_module_data_out[2] ;
 wire \sw_017_module_data_out[3] ;
 wire \sw_017_module_data_out[4] ;
 wire \sw_017_module_data_out[5] ;
 wire \sw_017_module_data_out[6] ;
 wire \sw_017_module_data_out[7] ;
 wire sw_017_scan_out;
 wire sw_018_clk_out;
 wire sw_018_data_out;
 wire sw_018_latch_out;
 wire \sw_018_module_data_in[0] ;
 wire \sw_018_module_data_in[1] ;
 wire \sw_018_module_data_in[2] ;
 wire \sw_018_module_data_in[3] ;
 wire \sw_018_module_data_in[4] ;
 wire \sw_018_module_data_in[5] ;
 wire \sw_018_module_data_in[6] ;
 wire \sw_018_module_data_in[7] ;
 wire \sw_018_module_data_out[0] ;
 wire \sw_018_module_data_out[1] ;
 wire \sw_018_module_data_out[2] ;
 wire \sw_018_module_data_out[3] ;
 wire \sw_018_module_data_out[4] ;
 wire \sw_018_module_data_out[5] ;
 wire \sw_018_module_data_out[6] ;
 wire \sw_018_module_data_out[7] ;
 wire sw_018_scan_out;
 wire sw_019_clk_out;
 wire sw_019_data_out;
 wire sw_019_latch_out;
 wire \sw_019_module_data_in[0] ;
 wire \sw_019_module_data_in[1] ;
 wire \sw_019_module_data_in[2] ;
 wire \sw_019_module_data_in[3] ;
 wire \sw_019_module_data_in[4] ;
 wire \sw_019_module_data_in[5] ;
 wire \sw_019_module_data_in[6] ;
 wire \sw_019_module_data_in[7] ;
 wire \sw_019_module_data_out[0] ;
 wire \sw_019_module_data_out[1] ;
 wire \sw_019_module_data_out[2] ;
 wire \sw_019_module_data_out[3] ;
 wire \sw_019_module_data_out[4] ;
 wire \sw_019_module_data_out[5] ;
 wire \sw_019_module_data_out[6] ;
 wire \sw_019_module_data_out[7] ;
 wire sw_019_scan_out;
 wire sw_020_clk_out;
 wire sw_020_data_out;
 wire sw_020_latch_out;
 wire \sw_020_module_data_in[0] ;
 wire \sw_020_module_data_in[1] ;
 wire \sw_020_module_data_in[2] ;
 wire \sw_020_module_data_in[3] ;
 wire \sw_020_module_data_in[4] ;
 wire \sw_020_module_data_in[5] ;
 wire \sw_020_module_data_in[6] ;
 wire \sw_020_module_data_in[7] ;
 wire \sw_020_module_data_out[0] ;
 wire \sw_020_module_data_out[1] ;
 wire \sw_020_module_data_out[2] ;
 wire \sw_020_module_data_out[3] ;
 wire \sw_020_module_data_out[4] ;
 wire \sw_020_module_data_out[5] ;
 wire \sw_020_module_data_out[6] ;
 wire \sw_020_module_data_out[7] ;
 wire sw_020_scan_out;
 wire sw_021_clk_out;
 wire sw_021_data_out;
 wire sw_021_latch_out;
 wire \sw_021_module_data_in[0] ;
 wire \sw_021_module_data_in[1] ;
 wire \sw_021_module_data_in[2] ;
 wire \sw_021_module_data_in[3] ;
 wire \sw_021_module_data_in[4] ;
 wire \sw_021_module_data_in[5] ;
 wire \sw_021_module_data_in[6] ;
 wire \sw_021_module_data_in[7] ;
 wire \sw_021_module_data_out[0] ;
 wire \sw_021_module_data_out[1] ;
 wire \sw_021_module_data_out[2] ;
 wire \sw_021_module_data_out[3] ;
 wire \sw_021_module_data_out[4] ;
 wire \sw_021_module_data_out[5] ;
 wire \sw_021_module_data_out[6] ;
 wire \sw_021_module_data_out[7] ;
 wire sw_021_scan_out;
 wire sw_022_clk_out;
 wire sw_022_data_out;
 wire sw_022_latch_out;
 wire \sw_022_module_data_in[0] ;
 wire \sw_022_module_data_in[1] ;
 wire \sw_022_module_data_in[2] ;
 wire \sw_022_module_data_in[3] ;
 wire \sw_022_module_data_in[4] ;
 wire \sw_022_module_data_in[5] ;
 wire \sw_022_module_data_in[6] ;
 wire \sw_022_module_data_in[7] ;
 wire \sw_022_module_data_out[0] ;
 wire \sw_022_module_data_out[1] ;
 wire \sw_022_module_data_out[2] ;
 wire \sw_022_module_data_out[3] ;
 wire \sw_022_module_data_out[4] ;
 wire \sw_022_module_data_out[5] ;
 wire \sw_022_module_data_out[6] ;
 wire \sw_022_module_data_out[7] ;
 wire sw_022_scan_out;
 wire sw_023_clk_out;
 wire sw_023_data_out;
 wire sw_023_latch_out;
 wire \sw_023_module_data_in[0] ;
 wire \sw_023_module_data_in[1] ;
 wire \sw_023_module_data_in[2] ;
 wire \sw_023_module_data_in[3] ;
 wire \sw_023_module_data_in[4] ;
 wire \sw_023_module_data_in[5] ;
 wire \sw_023_module_data_in[6] ;
 wire \sw_023_module_data_in[7] ;
 wire \sw_023_module_data_out[0] ;
 wire \sw_023_module_data_out[1] ;
 wire \sw_023_module_data_out[2] ;
 wire \sw_023_module_data_out[3] ;
 wire \sw_023_module_data_out[4] ;
 wire \sw_023_module_data_out[5] ;
 wire \sw_023_module_data_out[6] ;
 wire \sw_023_module_data_out[7] ;
 wire sw_023_scan_out;
 wire sw_024_clk_out;
 wire sw_024_data_out;
 wire sw_024_latch_out;
 wire \sw_024_module_data_in[0] ;
 wire \sw_024_module_data_in[1] ;
 wire \sw_024_module_data_in[2] ;
 wire \sw_024_module_data_in[3] ;
 wire \sw_024_module_data_in[4] ;
 wire \sw_024_module_data_in[5] ;
 wire \sw_024_module_data_in[6] ;
 wire \sw_024_module_data_in[7] ;
 wire \sw_024_module_data_out[0] ;
 wire \sw_024_module_data_out[1] ;
 wire \sw_024_module_data_out[2] ;
 wire \sw_024_module_data_out[3] ;
 wire \sw_024_module_data_out[4] ;
 wire \sw_024_module_data_out[5] ;
 wire \sw_024_module_data_out[6] ;
 wire \sw_024_module_data_out[7] ;
 wire sw_024_scan_out;
 wire sw_025_clk_out;
 wire sw_025_data_out;
 wire sw_025_latch_out;
 wire \sw_025_module_data_in[0] ;
 wire \sw_025_module_data_in[1] ;
 wire \sw_025_module_data_in[2] ;
 wire \sw_025_module_data_in[3] ;
 wire \sw_025_module_data_in[4] ;
 wire \sw_025_module_data_in[5] ;
 wire \sw_025_module_data_in[6] ;
 wire \sw_025_module_data_in[7] ;
 wire \sw_025_module_data_out[0] ;
 wire \sw_025_module_data_out[1] ;
 wire \sw_025_module_data_out[2] ;
 wire \sw_025_module_data_out[3] ;
 wire \sw_025_module_data_out[4] ;
 wire \sw_025_module_data_out[5] ;
 wire \sw_025_module_data_out[6] ;
 wire \sw_025_module_data_out[7] ;
 wire sw_025_scan_out;
 wire sw_026_clk_out;
 wire sw_026_data_out;
 wire sw_026_latch_out;
 wire \sw_026_module_data_in[0] ;
 wire \sw_026_module_data_in[1] ;
 wire \sw_026_module_data_in[2] ;
 wire \sw_026_module_data_in[3] ;
 wire \sw_026_module_data_in[4] ;
 wire \sw_026_module_data_in[5] ;
 wire \sw_026_module_data_in[6] ;
 wire \sw_026_module_data_in[7] ;
 wire \sw_026_module_data_out[0] ;
 wire \sw_026_module_data_out[1] ;
 wire \sw_026_module_data_out[2] ;
 wire \sw_026_module_data_out[3] ;
 wire \sw_026_module_data_out[4] ;
 wire \sw_026_module_data_out[5] ;
 wire \sw_026_module_data_out[6] ;
 wire \sw_026_module_data_out[7] ;
 wire sw_026_scan_out;
 wire sw_027_clk_out;
 wire sw_027_data_out;
 wire sw_027_latch_out;
 wire \sw_027_module_data_in[0] ;
 wire \sw_027_module_data_in[1] ;
 wire \sw_027_module_data_in[2] ;
 wire \sw_027_module_data_in[3] ;
 wire \sw_027_module_data_in[4] ;
 wire \sw_027_module_data_in[5] ;
 wire \sw_027_module_data_in[6] ;
 wire \sw_027_module_data_in[7] ;
 wire \sw_027_module_data_out[0] ;
 wire \sw_027_module_data_out[1] ;
 wire \sw_027_module_data_out[2] ;
 wire \sw_027_module_data_out[3] ;
 wire \sw_027_module_data_out[4] ;
 wire \sw_027_module_data_out[5] ;
 wire \sw_027_module_data_out[6] ;
 wire \sw_027_module_data_out[7] ;
 wire sw_027_scan_out;
 wire sw_028_clk_out;
 wire sw_028_data_out;
 wire sw_028_latch_out;
 wire \sw_028_module_data_in[0] ;
 wire \sw_028_module_data_in[1] ;
 wire \sw_028_module_data_in[2] ;
 wire \sw_028_module_data_in[3] ;
 wire \sw_028_module_data_in[4] ;
 wire \sw_028_module_data_in[5] ;
 wire \sw_028_module_data_in[6] ;
 wire \sw_028_module_data_in[7] ;
 wire \sw_028_module_data_out[0] ;
 wire \sw_028_module_data_out[1] ;
 wire \sw_028_module_data_out[2] ;
 wire \sw_028_module_data_out[3] ;
 wire \sw_028_module_data_out[4] ;
 wire \sw_028_module_data_out[5] ;
 wire \sw_028_module_data_out[6] ;
 wire \sw_028_module_data_out[7] ;
 wire sw_028_scan_out;
 wire sw_029_clk_out;
 wire sw_029_data_out;
 wire sw_029_latch_out;
 wire \sw_029_module_data_in[0] ;
 wire \sw_029_module_data_in[1] ;
 wire \sw_029_module_data_in[2] ;
 wire \sw_029_module_data_in[3] ;
 wire \sw_029_module_data_in[4] ;
 wire \sw_029_module_data_in[5] ;
 wire \sw_029_module_data_in[6] ;
 wire \sw_029_module_data_in[7] ;
 wire \sw_029_module_data_out[0] ;
 wire \sw_029_module_data_out[1] ;
 wire \sw_029_module_data_out[2] ;
 wire \sw_029_module_data_out[3] ;
 wire \sw_029_module_data_out[4] ;
 wire \sw_029_module_data_out[5] ;
 wire \sw_029_module_data_out[6] ;
 wire \sw_029_module_data_out[7] ;
 wire sw_029_scan_out;
 wire sw_030_clk_out;
 wire sw_030_data_out;
 wire sw_030_latch_out;
 wire \sw_030_module_data_in[0] ;
 wire \sw_030_module_data_in[1] ;
 wire \sw_030_module_data_in[2] ;
 wire \sw_030_module_data_in[3] ;
 wire \sw_030_module_data_in[4] ;
 wire \sw_030_module_data_in[5] ;
 wire \sw_030_module_data_in[6] ;
 wire \sw_030_module_data_in[7] ;
 wire \sw_030_module_data_out[0] ;
 wire \sw_030_module_data_out[1] ;
 wire \sw_030_module_data_out[2] ;
 wire \sw_030_module_data_out[3] ;
 wire \sw_030_module_data_out[4] ;
 wire \sw_030_module_data_out[5] ;
 wire \sw_030_module_data_out[6] ;
 wire \sw_030_module_data_out[7] ;
 wire sw_030_scan_out;
 wire sw_031_clk_out;
 wire sw_031_data_out;
 wire sw_031_latch_out;
 wire \sw_031_module_data_in[0] ;
 wire \sw_031_module_data_in[1] ;
 wire \sw_031_module_data_in[2] ;
 wire \sw_031_module_data_in[3] ;
 wire \sw_031_module_data_in[4] ;
 wire \sw_031_module_data_in[5] ;
 wire \sw_031_module_data_in[6] ;
 wire \sw_031_module_data_in[7] ;
 wire \sw_031_module_data_out[0] ;
 wire \sw_031_module_data_out[1] ;
 wire \sw_031_module_data_out[2] ;
 wire \sw_031_module_data_out[3] ;
 wire \sw_031_module_data_out[4] ;
 wire \sw_031_module_data_out[5] ;
 wire \sw_031_module_data_out[6] ;
 wire \sw_031_module_data_out[7] ;
 wire sw_031_scan_out;
 wire sw_032_clk_out;
 wire sw_032_data_out;
 wire sw_032_latch_out;
 wire \sw_032_module_data_in[0] ;
 wire \sw_032_module_data_in[1] ;
 wire \sw_032_module_data_in[2] ;
 wire \sw_032_module_data_in[3] ;
 wire \sw_032_module_data_in[4] ;
 wire \sw_032_module_data_in[5] ;
 wire \sw_032_module_data_in[6] ;
 wire \sw_032_module_data_in[7] ;
 wire \sw_032_module_data_out[0] ;
 wire \sw_032_module_data_out[1] ;
 wire \sw_032_module_data_out[2] ;
 wire \sw_032_module_data_out[3] ;
 wire \sw_032_module_data_out[4] ;
 wire \sw_032_module_data_out[5] ;
 wire \sw_032_module_data_out[6] ;
 wire \sw_032_module_data_out[7] ;
 wire sw_032_scan_out;
 wire sw_033_clk_out;
 wire sw_033_data_out;
 wire sw_033_latch_out;
 wire \sw_033_module_data_in[0] ;
 wire \sw_033_module_data_in[1] ;
 wire \sw_033_module_data_in[2] ;
 wire \sw_033_module_data_in[3] ;
 wire \sw_033_module_data_in[4] ;
 wire \sw_033_module_data_in[5] ;
 wire \sw_033_module_data_in[6] ;
 wire \sw_033_module_data_in[7] ;
 wire \sw_033_module_data_out[0] ;
 wire \sw_033_module_data_out[1] ;
 wire \sw_033_module_data_out[2] ;
 wire \sw_033_module_data_out[3] ;
 wire \sw_033_module_data_out[4] ;
 wire \sw_033_module_data_out[5] ;
 wire \sw_033_module_data_out[6] ;
 wire \sw_033_module_data_out[7] ;
 wire sw_033_scan_out;
 wire sw_034_clk_out;
 wire sw_034_data_out;
 wire sw_034_latch_out;
 wire \sw_034_module_data_in[0] ;
 wire \sw_034_module_data_in[1] ;
 wire \sw_034_module_data_in[2] ;
 wire \sw_034_module_data_in[3] ;
 wire \sw_034_module_data_in[4] ;
 wire \sw_034_module_data_in[5] ;
 wire \sw_034_module_data_in[6] ;
 wire \sw_034_module_data_in[7] ;
 wire \sw_034_module_data_out[0] ;
 wire \sw_034_module_data_out[1] ;
 wire \sw_034_module_data_out[2] ;
 wire \sw_034_module_data_out[3] ;
 wire \sw_034_module_data_out[4] ;
 wire \sw_034_module_data_out[5] ;
 wire \sw_034_module_data_out[6] ;
 wire \sw_034_module_data_out[7] ;
 wire sw_034_scan_out;
 wire sw_035_clk_out;
 wire sw_035_data_out;
 wire sw_035_latch_out;
 wire \sw_035_module_data_in[0] ;
 wire \sw_035_module_data_in[1] ;
 wire \sw_035_module_data_in[2] ;
 wire \sw_035_module_data_in[3] ;
 wire \sw_035_module_data_in[4] ;
 wire \sw_035_module_data_in[5] ;
 wire \sw_035_module_data_in[6] ;
 wire \sw_035_module_data_in[7] ;
 wire \sw_035_module_data_out[0] ;
 wire \sw_035_module_data_out[1] ;
 wire \sw_035_module_data_out[2] ;
 wire \sw_035_module_data_out[3] ;
 wire \sw_035_module_data_out[4] ;
 wire \sw_035_module_data_out[5] ;
 wire \sw_035_module_data_out[6] ;
 wire \sw_035_module_data_out[7] ;
 wire sw_035_scan_out;
 wire sw_036_clk_out;
 wire sw_036_data_out;
 wire sw_036_latch_out;
 wire \sw_036_module_data_in[0] ;
 wire \sw_036_module_data_in[1] ;
 wire \sw_036_module_data_in[2] ;
 wire \sw_036_module_data_in[3] ;
 wire \sw_036_module_data_in[4] ;
 wire \sw_036_module_data_in[5] ;
 wire \sw_036_module_data_in[6] ;
 wire \sw_036_module_data_in[7] ;
 wire \sw_036_module_data_out[0] ;
 wire \sw_036_module_data_out[1] ;
 wire \sw_036_module_data_out[2] ;
 wire \sw_036_module_data_out[3] ;
 wire \sw_036_module_data_out[4] ;
 wire \sw_036_module_data_out[5] ;
 wire \sw_036_module_data_out[6] ;
 wire \sw_036_module_data_out[7] ;
 wire sw_036_scan_out;
 wire sw_037_clk_out;
 wire sw_037_data_out;
 wire sw_037_latch_out;
 wire \sw_037_module_data_in[0] ;
 wire \sw_037_module_data_in[1] ;
 wire \sw_037_module_data_in[2] ;
 wire \sw_037_module_data_in[3] ;
 wire \sw_037_module_data_in[4] ;
 wire \sw_037_module_data_in[5] ;
 wire \sw_037_module_data_in[6] ;
 wire \sw_037_module_data_in[7] ;
 wire \sw_037_module_data_out[0] ;
 wire \sw_037_module_data_out[1] ;
 wire \sw_037_module_data_out[2] ;
 wire \sw_037_module_data_out[3] ;
 wire \sw_037_module_data_out[4] ;
 wire \sw_037_module_data_out[5] ;
 wire \sw_037_module_data_out[6] ;
 wire \sw_037_module_data_out[7] ;
 wire sw_037_scan_out;
 wire sw_038_clk_out;
 wire sw_038_data_out;
 wire sw_038_latch_out;
 wire \sw_038_module_data_in[0] ;
 wire \sw_038_module_data_in[1] ;
 wire \sw_038_module_data_in[2] ;
 wire \sw_038_module_data_in[3] ;
 wire \sw_038_module_data_in[4] ;
 wire \sw_038_module_data_in[5] ;
 wire \sw_038_module_data_in[6] ;
 wire \sw_038_module_data_in[7] ;
 wire \sw_038_module_data_out[0] ;
 wire \sw_038_module_data_out[1] ;
 wire \sw_038_module_data_out[2] ;
 wire \sw_038_module_data_out[3] ;
 wire \sw_038_module_data_out[4] ;
 wire \sw_038_module_data_out[5] ;
 wire \sw_038_module_data_out[6] ;
 wire \sw_038_module_data_out[7] ;
 wire sw_038_scan_out;
 wire sw_039_clk_out;
 wire sw_039_data_out;
 wire sw_039_latch_out;
 wire \sw_039_module_data_in[0] ;
 wire \sw_039_module_data_in[1] ;
 wire \sw_039_module_data_in[2] ;
 wire \sw_039_module_data_in[3] ;
 wire \sw_039_module_data_in[4] ;
 wire \sw_039_module_data_in[5] ;
 wire \sw_039_module_data_in[6] ;
 wire \sw_039_module_data_in[7] ;
 wire \sw_039_module_data_out[0] ;
 wire \sw_039_module_data_out[1] ;
 wire \sw_039_module_data_out[2] ;
 wire \sw_039_module_data_out[3] ;
 wire \sw_039_module_data_out[4] ;
 wire \sw_039_module_data_out[5] ;
 wire \sw_039_module_data_out[6] ;
 wire \sw_039_module_data_out[7] ;
 wire sw_039_scan_out;
 wire sw_040_clk_out;
 wire sw_040_data_out;
 wire sw_040_latch_out;
 wire \sw_040_module_data_in[0] ;
 wire \sw_040_module_data_in[1] ;
 wire \sw_040_module_data_in[2] ;
 wire \sw_040_module_data_in[3] ;
 wire \sw_040_module_data_in[4] ;
 wire \sw_040_module_data_in[5] ;
 wire \sw_040_module_data_in[6] ;
 wire \sw_040_module_data_in[7] ;
 wire \sw_040_module_data_out[0] ;
 wire \sw_040_module_data_out[1] ;
 wire \sw_040_module_data_out[2] ;
 wire \sw_040_module_data_out[3] ;
 wire \sw_040_module_data_out[4] ;
 wire \sw_040_module_data_out[5] ;
 wire \sw_040_module_data_out[6] ;
 wire \sw_040_module_data_out[7] ;
 wire sw_040_scan_out;
 wire sw_041_clk_out;
 wire sw_041_data_out;
 wire sw_041_latch_out;
 wire \sw_041_module_data_in[0] ;
 wire \sw_041_module_data_in[1] ;
 wire \sw_041_module_data_in[2] ;
 wire \sw_041_module_data_in[3] ;
 wire \sw_041_module_data_in[4] ;
 wire \sw_041_module_data_in[5] ;
 wire \sw_041_module_data_in[6] ;
 wire \sw_041_module_data_in[7] ;
 wire \sw_041_module_data_out[0] ;
 wire \sw_041_module_data_out[1] ;
 wire \sw_041_module_data_out[2] ;
 wire \sw_041_module_data_out[3] ;
 wire \sw_041_module_data_out[4] ;
 wire \sw_041_module_data_out[5] ;
 wire \sw_041_module_data_out[6] ;
 wire \sw_041_module_data_out[7] ;
 wire sw_041_scan_out;
 wire sw_042_clk_out;
 wire sw_042_data_out;
 wire sw_042_latch_out;
 wire \sw_042_module_data_in[0] ;
 wire \sw_042_module_data_in[1] ;
 wire \sw_042_module_data_in[2] ;
 wire \sw_042_module_data_in[3] ;
 wire \sw_042_module_data_in[4] ;
 wire \sw_042_module_data_in[5] ;
 wire \sw_042_module_data_in[6] ;
 wire \sw_042_module_data_in[7] ;
 wire \sw_042_module_data_out[0] ;
 wire \sw_042_module_data_out[1] ;
 wire \sw_042_module_data_out[2] ;
 wire \sw_042_module_data_out[3] ;
 wire \sw_042_module_data_out[4] ;
 wire \sw_042_module_data_out[5] ;
 wire \sw_042_module_data_out[6] ;
 wire \sw_042_module_data_out[7] ;
 wire sw_042_scan_out;
 wire sw_043_clk_out;
 wire sw_043_data_out;
 wire sw_043_latch_out;
 wire \sw_043_module_data_in[0] ;
 wire \sw_043_module_data_in[1] ;
 wire \sw_043_module_data_in[2] ;
 wire \sw_043_module_data_in[3] ;
 wire \sw_043_module_data_in[4] ;
 wire \sw_043_module_data_in[5] ;
 wire \sw_043_module_data_in[6] ;
 wire \sw_043_module_data_in[7] ;
 wire \sw_043_module_data_out[0] ;
 wire \sw_043_module_data_out[1] ;
 wire \sw_043_module_data_out[2] ;
 wire \sw_043_module_data_out[3] ;
 wire \sw_043_module_data_out[4] ;
 wire \sw_043_module_data_out[5] ;
 wire \sw_043_module_data_out[6] ;
 wire \sw_043_module_data_out[7] ;
 wire sw_043_scan_out;
 wire sw_044_clk_out;
 wire sw_044_data_out;
 wire sw_044_latch_out;
 wire \sw_044_module_data_in[0] ;
 wire \sw_044_module_data_in[1] ;
 wire \sw_044_module_data_in[2] ;
 wire \sw_044_module_data_in[3] ;
 wire \sw_044_module_data_in[4] ;
 wire \sw_044_module_data_in[5] ;
 wire \sw_044_module_data_in[6] ;
 wire \sw_044_module_data_in[7] ;
 wire \sw_044_module_data_out[0] ;
 wire \sw_044_module_data_out[1] ;
 wire \sw_044_module_data_out[2] ;
 wire \sw_044_module_data_out[3] ;
 wire \sw_044_module_data_out[4] ;
 wire \sw_044_module_data_out[5] ;
 wire \sw_044_module_data_out[6] ;
 wire \sw_044_module_data_out[7] ;
 wire sw_044_scan_out;
 wire sw_045_clk_out;
 wire sw_045_data_out;
 wire sw_045_latch_out;
 wire \sw_045_module_data_in[0] ;
 wire \sw_045_module_data_in[1] ;
 wire \sw_045_module_data_in[2] ;
 wire \sw_045_module_data_in[3] ;
 wire \sw_045_module_data_in[4] ;
 wire \sw_045_module_data_in[5] ;
 wire \sw_045_module_data_in[6] ;
 wire \sw_045_module_data_in[7] ;
 wire \sw_045_module_data_out[0] ;
 wire \sw_045_module_data_out[1] ;
 wire \sw_045_module_data_out[2] ;
 wire \sw_045_module_data_out[3] ;
 wire \sw_045_module_data_out[4] ;
 wire \sw_045_module_data_out[5] ;
 wire \sw_045_module_data_out[6] ;
 wire \sw_045_module_data_out[7] ;
 wire sw_045_scan_out;
 wire sw_046_clk_out;
 wire sw_046_data_out;
 wire sw_046_latch_out;
 wire \sw_046_module_data_in[0] ;
 wire \sw_046_module_data_in[1] ;
 wire \sw_046_module_data_in[2] ;
 wire \sw_046_module_data_in[3] ;
 wire \sw_046_module_data_in[4] ;
 wire \sw_046_module_data_in[5] ;
 wire \sw_046_module_data_in[6] ;
 wire \sw_046_module_data_in[7] ;
 wire \sw_046_module_data_out[0] ;
 wire \sw_046_module_data_out[1] ;
 wire \sw_046_module_data_out[2] ;
 wire \sw_046_module_data_out[3] ;
 wire \sw_046_module_data_out[4] ;
 wire \sw_046_module_data_out[5] ;
 wire \sw_046_module_data_out[6] ;
 wire \sw_046_module_data_out[7] ;
 wire sw_046_scan_out;
 wire sw_047_clk_out;
 wire sw_047_data_out;
 wire sw_047_latch_out;
 wire \sw_047_module_data_in[0] ;
 wire \sw_047_module_data_in[1] ;
 wire \sw_047_module_data_in[2] ;
 wire \sw_047_module_data_in[3] ;
 wire \sw_047_module_data_in[4] ;
 wire \sw_047_module_data_in[5] ;
 wire \sw_047_module_data_in[6] ;
 wire \sw_047_module_data_in[7] ;
 wire \sw_047_module_data_out[0] ;
 wire \sw_047_module_data_out[1] ;
 wire \sw_047_module_data_out[2] ;
 wire \sw_047_module_data_out[3] ;
 wire \sw_047_module_data_out[4] ;
 wire \sw_047_module_data_out[5] ;
 wire \sw_047_module_data_out[6] ;
 wire \sw_047_module_data_out[7] ;
 wire sw_047_scan_out;
 wire sw_048_clk_out;
 wire sw_048_data_out;
 wire sw_048_latch_out;
 wire \sw_048_module_data_in[0] ;
 wire \sw_048_module_data_in[1] ;
 wire \sw_048_module_data_in[2] ;
 wire \sw_048_module_data_in[3] ;
 wire \sw_048_module_data_in[4] ;
 wire \sw_048_module_data_in[5] ;
 wire \sw_048_module_data_in[6] ;
 wire \sw_048_module_data_in[7] ;
 wire \sw_048_module_data_out[0] ;
 wire \sw_048_module_data_out[1] ;
 wire \sw_048_module_data_out[2] ;
 wire \sw_048_module_data_out[3] ;
 wire \sw_048_module_data_out[4] ;
 wire \sw_048_module_data_out[5] ;
 wire \sw_048_module_data_out[6] ;
 wire \sw_048_module_data_out[7] ;
 wire sw_048_scan_out;
 wire sw_049_clk_out;
 wire sw_049_data_out;
 wire sw_049_latch_out;
 wire \sw_049_module_data_in[0] ;
 wire \sw_049_module_data_in[1] ;
 wire \sw_049_module_data_in[2] ;
 wire \sw_049_module_data_in[3] ;
 wire \sw_049_module_data_in[4] ;
 wire \sw_049_module_data_in[5] ;
 wire \sw_049_module_data_in[6] ;
 wire \sw_049_module_data_in[7] ;
 wire \sw_049_module_data_out[0] ;
 wire \sw_049_module_data_out[1] ;
 wire \sw_049_module_data_out[2] ;
 wire \sw_049_module_data_out[3] ;
 wire \sw_049_module_data_out[4] ;
 wire \sw_049_module_data_out[5] ;
 wire \sw_049_module_data_out[6] ;
 wire \sw_049_module_data_out[7] ;
 wire sw_049_scan_out;
 wire sw_050_clk_out;
 wire sw_050_data_out;
 wire sw_050_latch_out;
 wire \sw_050_module_data_in[0] ;
 wire \sw_050_module_data_in[1] ;
 wire \sw_050_module_data_in[2] ;
 wire \sw_050_module_data_in[3] ;
 wire \sw_050_module_data_in[4] ;
 wire \sw_050_module_data_in[5] ;
 wire \sw_050_module_data_in[6] ;
 wire \sw_050_module_data_in[7] ;
 wire \sw_050_module_data_out[0] ;
 wire \sw_050_module_data_out[1] ;
 wire \sw_050_module_data_out[2] ;
 wire \sw_050_module_data_out[3] ;
 wire \sw_050_module_data_out[4] ;
 wire \sw_050_module_data_out[5] ;
 wire \sw_050_module_data_out[6] ;
 wire \sw_050_module_data_out[7] ;
 wire sw_050_scan_out;
 wire sw_051_clk_out;
 wire sw_051_data_out;
 wire sw_051_latch_out;
 wire \sw_051_module_data_in[0] ;
 wire \sw_051_module_data_in[1] ;
 wire \sw_051_module_data_in[2] ;
 wire \sw_051_module_data_in[3] ;
 wire \sw_051_module_data_in[4] ;
 wire \sw_051_module_data_in[5] ;
 wire \sw_051_module_data_in[6] ;
 wire \sw_051_module_data_in[7] ;
 wire \sw_051_module_data_out[0] ;
 wire \sw_051_module_data_out[1] ;
 wire \sw_051_module_data_out[2] ;
 wire \sw_051_module_data_out[3] ;
 wire \sw_051_module_data_out[4] ;
 wire \sw_051_module_data_out[5] ;
 wire \sw_051_module_data_out[6] ;
 wire \sw_051_module_data_out[7] ;
 wire sw_051_scan_out;
 wire sw_052_clk_out;
 wire sw_052_data_out;
 wire sw_052_latch_out;
 wire \sw_052_module_data_in[0] ;
 wire \sw_052_module_data_in[1] ;
 wire \sw_052_module_data_in[2] ;
 wire \sw_052_module_data_in[3] ;
 wire \sw_052_module_data_in[4] ;
 wire \sw_052_module_data_in[5] ;
 wire \sw_052_module_data_in[6] ;
 wire \sw_052_module_data_in[7] ;
 wire \sw_052_module_data_out[0] ;
 wire \sw_052_module_data_out[1] ;
 wire \sw_052_module_data_out[2] ;
 wire \sw_052_module_data_out[3] ;
 wire \sw_052_module_data_out[4] ;
 wire \sw_052_module_data_out[5] ;
 wire \sw_052_module_data_out[6] ;
 wire \sw_052_module_data_out[7] ;
 wire sw_052_scan_out;
 wire sw_053_clk_out;
 wire sw_053_data_out;
 wire sw_053_latch_out;
 wire \sw_053_module_data_in[0] ;
 wire \sw_053_module_data_in[1] ;
 wire \sw_053_module_data_in[2] ;
 wire \sw_053_module_data_in[3] ;
 wire \sw_053_module_data_in[4] ;
 wire \sw_053_module_data_in[5] ;
 wire \sw_053_module_data_in[6] ;
 wire \sw_053_module_data_in[7] ;
 wire \sw_053_module_data_out[0] ;
 wire \sw_053_module_data_out[1] ;
 wire \sw_053_module_data_out[2] ;
 wire \sw_053_module_data_out[3] ;
 wire \sw_053_module_data_out[4] ;
 wire \sw_053_module_data_out[5] ;
 wire \sw_053_module_data_out[6] ;
 wire \sw_053_module_data_out[7] ;
 wire sw_053_scan_out;
 wire sw_054_clk_out;
 wire sw_054_data_out;
 wire sw_054_latch_out;
 wire \sw_054_module_data_in[0] ;
 wire \sw_054_module_data_in[1] ;
 wire \sw_054_module_data_in[2] ;
 wire \sw_054_module_data_in[3] ;
 wire \sw_054_module_data_in[4] ;
 wire \sw_054_module_data_in[5] ;
 wire \sw_054_module_data_in[6] ;
 wire \sw_054_module_data_in[7] ;
 wire \sw_054_module_data_out[0] ;
 wire \sw_054_module_data_out[1] ;
 wire \sw_054_module_data_out[2] ;
 wire \sw_054_module_data_out[3] ;
 wire \sw_054_module_data_out[4] ;
 wire \sw_054_module_data_out[5] ;
 wire \sw_054_module_data_out[6] ;
 wire \sw_054_module_data_out[7] ;
 wire sw_054_scan_out;
 wire sw_055_clk_out;
 wire sw_055_data_out;
 wire sw_055_latch_out;
 wire \sw_055_module_data_in[0] ;
 wire \sw_055_module_data_in[1] ;
 wire \sw_055_module_data_in[2] ;
 wire \sw_055_module_data_in[3] ;
 wire \sw_055_module_data_in[4] ;
 wire \sw_055_module_data_in[5] ;
 wire \sw_055_module_data_in[6] ;
 wire \sw_055_module_data_in[7] ;
 wire \sw_055_module_data_out[0] ;
 wire \sw_055_module_data_out[1] ;
 wire \sw_055_module_data_out[2] ;
 wire \sw_055_module_data_out[3] ;
 wire \sw_055_module_data_out[4] ;
 wire \sw_055_module_data_out[5] ;
 wire \sw_055_module_data_out[6] ;
 wire \sw_055_module_data_out[7] ;
 wire sw_055_scan_out;
 wire sw_056_clk_out;
 wire sw_056_data_out;
 wire sw_056_latch_out;
 wire \sw_056_module_data_in[0] ;
 wire \sw_056_module_data_in[1] ;
 wire \sw_056_module_data_in[2] ;
 wire \sw_056_module_data_in[3] ;
 wire \sw_056_module_data_in[4] ;
 wire \sw_056_module_data_in[5] ;
 wire \sw_056_module_data_in[6] ;
 wire \sw_056_module_data_in[7] ;
 wire \sw_056_module_data_out[0] ;
 wire \sw_056_module_data_out[1] ;
 wire \sw_056_module_data_out[2] ;
 wire \sw_056_module_data_out[3] ;
 wire \sw_056_module_data_out[4] ;
 wire \sw_056_module_data_out[5] ;
 wire \sw_056_module_data_out[6] ;
 wire \sw_056_module_data_out[7] ;
 wire sw_056_scan_out;
 wire sw_057_clk_out;
 wire sw_057_data_out;
 wire sw_057_latch_out;
 wire \sw_057_module_data_in[0] ;
 wire \sw_057_module_data_in[1] ;
 wire \sw_057_module_data_in[2] ;
 wire \sw_057_module_data_in[3] ;
 wire \sw_057_module_data_in[4] ;
 wire \sw_057_module_data_in[5] ;
 wire \sw_057_module_data_in[6] ;
 wire \sw_057_module_data_in[7] ;
 wire \sw_057_module_data_out[0] ;
 wire \sw_057_module_data_out[1] ;
 wire \sw_057_module_data_out[2] ;
 wire \sw_057_module_data_out[3] ;
 wire \sw_057_module_data_out[4] ;
 wire \sw_057_module_data_out[5] ;
 wire \sw_057_module_data_out[6] ;
 wire \sw_057_module_data_out[7] ;
 wire sw_057_scan_out;
 wire sw_058_clk_out;
 wire sw_058_data_out;
 wire sw_058_latch_out;
 wire \sw_058_module_data_in[0] ;
 wire \sw_058_module_data_in[1] ;
 wire \sw_058_module_data_in[2] ;
 wire \sw_058_module_data_in[3] ;
 wire \sw_058_module_data_in[4] ;
 wire \sw_058_module_data_in[5] ;
 wire \sw_058_module_data_in[6] ;
 wire \sw_058_module_data_in[7] ;
 wire \sw_058_module_data_out[0] ;
 wire \sw_058_module_data_out[1] ;
 wire \sw_058_module_data_out[2] ;
 wire \sw_058_module_data_out[3] ;
 wire \sw_058_module_data_out[4] ;
 wire \sw_058_module_data_out[5] ;
 wire \sw_058_module_data_out[6] ;
 wire \sw_058_module_data_out[7] ;
 wire sw_058_scan_out;
 wire sw_059_clk_out;
 wire sw_059_data_out;
 wire sw_059_latch_out;
 wire \sw_059_module_data_in[0] ;
 wire \sw_059_module_data_in[1] ;
 wire \sw_059_module_data_in[2] ;
 wire \sw_059_module_data_in[3] ;
 wire \sw_059_module_data_in[4] ;
 wire \sw_059_module_data_in[5] ;
 wire \sw_059_module_data_in[6] ;
 wire \sw_059_module_data_in[7] ;
 wire \sw_059_module_data_out[0] ;
 wire \sw_059_module_data_out[1] ;
 wire \sw_059_module_data_out[2] ;
 wire \sw_059_module_data_out[3] ;
 wire \sw_059_module_data_out[4] ;
 wire \sw_059_module_data_out[5] ;
 wire \sw_059_module_data_out[6] ;
 wire \sw_059_module_data_out[7] ;
 wire sw_059_scan_out;
 wire sw_060_clk_out;
 wire sw_060_data_out;
 wire sw_060_latch_out;
 wire \sw_060_module_data_in[0] ;
 wire \sw_060_module_data_in[1] ;
 wire \sw_060_module_data_in[2] ;
 wire \sw_060_module_data_in[3] ;
 wire \sw_060_module_data_in[4] ;
 wire \sw_060_module_data_in[5] ;
 wire \sw_060_module_data_in[6] ;
 wire \sw_060_module_data_in[7] ;
 wire \sw_060_module_data_out[0] ;
 wire \sw_060_module_data_out[1] ;
 wire \sw_060_module_data_out[2] ;
 wire \sw_060_module_data_out[3] ;
 wire \sw_060_module_data_out[4] ;
 wire \sw_060_module_data_out[5] ;
 wire \sw_060_module_data_out[6] ;
 wire \sw_060_module_data_out[7] ;
 wire sw_060_scan_out;
 wire sw_061_clk_out;
 wire sw_061_data_out;
 wire sw_061_latch_out;
 wire \sw_061_module_data_in[0] ;
 wire \sw_061_module_data_in[1] ;
 wire \sw_061_module_data_in[2] ;
 wire \sw_061_module_data_in[3] ;
 wire \sw_061_module_data_in[4] ;
 wire \sw_061_module_data_in[5] ;
 wire \sw_061_module_data_in[6] ;
 wire \sw_061_module_data_in[7] ;
 wire \sw_061_module_data_out[0] ;
 wire \sw_061_module_data_out[1] ;
 wire \sw_061_module_data_out[2] ;
 wire \sw_061_module_data_out[3] ;
 wire \sw_061_module_data_out[4] ;
 wire \sw_061_module_data_out[5] ;
 wire \sw_061_module_data_out[6] ;
 wire \sw_061_module_data_out[7] ;
 wire sw_061_scan_out;
 wire sw_062_clk_out;
 wire sw_062_data_out;
 wire sw_062_latch_out;
 wire \sw_062_module_data_in[0] ;
 wire \sw_062_module_data_in[1] ;
 wire \sw_062_module_data_in[2] ;
 wire \sw_062_module_data_in[3] ;
 wire \sw_062_module_data_in[4] ;
 wire \sw_062_module_data_in[5] ;
 wire \sw_062_module_data_in[6] ;
 wire \sw_062_module_data_in[7] ;
 wire \sw_062_module_data_out[0] ;
 wire \sw_062_module_data_out[1] ;
 wire \sw_062_module_data_out[2] ;
 wire \sw_062_module_data_out[3] ;
 wire \sw_062_module_data_out[4] ;
 wire \sw_062_module_data_out[5] ;
 wire \sw_062_module_data_out[6] ;
 wire \sw_062_module_data_out[7] ;
 wire sw_062_scan_out;
 wire sw_063_clk_out;
 wire sw_063_data_out;
 wire sw_063_latch_out;
 wire \sw_063_module_data_in[0] ;
 wire \sw_063_module_data_in[1] ;
 wire \sw_063_module_data_in[2] ;
 wire \sw_063_module_data_in[3] ;
 wire \sw_063_module_data_in[4] ;
 wire \sw_063_module_data_in[5] ;
 wire \sw_063_module_data_in[6] ;
 wire \sw_063_module_data_in[7] ;
 wire \sw_063_module_data_out[0] ;
 wire \sw_063_module_data_out[1] ;
 wire \sw_063_module_data_out[2] ;
 wire \sw_063_module_data_out[3] ;
 wire \sw_063_module_data_out[4] ;
 wire \sw_063_module_data_out[5] ;
 wire \sw_063_module_data_out[6] ;
 wire \sw_063_module_data_out[7] ;
 wire sw_063_scan_out;
 wire sw_064_clk_out;
 wire sw_064_data_out;
 wire sw_064_latch_out;
 wire \sw_064_module_data_in[0] ;
 wire \sw_064_module_data_in[1] ;
 wire \sw_064_module_data_in[2] ;
 wire \sw_064_module_data_in[3] ;
 wire \sw_064_module_data_in[4] ;
 wire \sw_064_module_data_in[5] ;
 wire \sw_064_module_data_in[6] ;
 wire \sw_064_module_data_in[7] ;
 wire \sw_064_module_data_out[0] ;
 wire \sw_064_module_data_out[1] ;
 wire \sw_064_module_data_out[2] ;
 wire \sw_064_module_data_out[3] ;
 wire \sw_064_module_data_out[4] ;
 wire \sw_064_module_data_out[5] ;
 wire \sw_064_module_data_out[6] ;
 wire \sw_064_module_data_out[7] ;
 wire sw_064_scan_out;
 wire sw_065_clk_out;
 wire sw_065_data_out;
 wire sw_065_latch_out;
 wire \sw_065_module_data_in[0] ;
 wire \sw_065_module_data_in[1] ;
 wire \sw_065_module_data_in[2] ;
 wire \sw_065_module_data_in[3] ;
 wire \sw_065_module_data_in[4] ;
 wire \sw_065_module_data_in[5] ;
 wire \sw_065_module_data_in[6] ;
 wire \sw_065_module_data_in[7] ;
 wire \sw_065_module_data_out[0] ;
 wire \sw_065_module_data_out[1] ;
 wire \sw_065_module_data_out[2] ;
 wire \sw_065_module_data_out[3] ;
 wire \sw_065_module_data_out[4] ;
 wire \sw_065_module_data_out[5] ;
 wire \sw_065_module_data_out[6] ;
 wire \sw_065_module_data_out[7] ;
 wire sw_065_scan_out;
 wire sw_066_clk_out;
 wire sw_066_data_out;
 wire sw_066_latch_out;
 wire \sw_066_module_data_in[0] ;
 wire \sw_066_module_data_in[1] ;
 wire \sw_066_module_data_in[2] ;
 wire \sw_066_module_data_in[3] ;
 wire \sw_066_module_data_in[4] ;
 wire \sw_066_module_data_in[5] ;
 wire \sw_066_module_data_in[6] ;
 wire \sw_066_module_data_in[7] ;
 wire \sw_066_module_data_out[0] ;
 wire \sw_066_module_data_out[1] ;
 wire \sw_066_module_data_out[2] ;
 wire \sw_066_module_data_out[3] ;
 wire \sw_066_module_data_out[4] ;
 wire \sw_066_module_data_out[5] ;
 wire \sw_066_module_data_out[6] ;
 wire \sw_066_module_data_out[7] ;
 wire sw_066_scan_out;
 wire sw_067_clk_out;
 wire sw_067_data_out;
 wire sw_067_latch_out;
 wire \sw_067_module_data_in[0] ;
 wire \sw_067_module_data_in[1] ;
 wire \sw_067_module_data_in[2] ;
 wire \sw_067_module_data_in[3] ;
 wire \sw_067_module_data_in[4] ;
 wire \sw_067_module_data_in[5] ;
 wire \sw_067_module_data_in[6] ;
 wire \sw_067_module_data_in[7] ;
 wire \sw_067_module_data_out[0] ;
 wire \sw_067_module_data_out[1] ;
 wire \sw_067_module_data_out[2] ;
 wire \sw_067_module_data_out[3] ;
 wire \sw_067_module_data_out[4] ;
 wire \sw_067_module_data_out[5] ;
 wire \sw_067_module_data_out[6] ;
 wire \sw_067_module_data_out[7] ;
 wire sw_067_scan_out;
 wire sw_068_clk_out;
 wire sw_068_data_out;
 wire sw_068_latch_out;
 wire \sw_068_module_data_in[0] ;
 wire \sw_068_module_data_in[1] ;
 wire \sw_068_module_data_in[2] ;
 wire \sw_068_module_data_in[3] ;
 wire \sw_068_module_data_in[4] ;
 wire \sw_068_module_data_in[5] ;
 wire \sw_068_module_data_in[6] ;
 wire \sw_068_module_data_in[7] ;
 wire \sw_068_module_data_out[0] ;
 wire \sw_068_module_data_out[1] ;
 wire \sw_068_module_data_out[2] ;
 wire \sw_068_module_data_out[3] ;
 wire \sw_068_module_data_out[4] ;
 wire \sw_068_module_data_out[5] ;
 wire \sw_068_module_data_out[6] ;
 wire \sw_068_module_data_out[7] ;
 wire sw_068_scan_out;
 wire sw_069_clk_out;
 wire sw_069_data_out;
 wire sw_069_latch_out;
 wire \sw_069_module_data_in[0] ;
 wire \sw_069_module_data_in[1] ;
 wire \sw_069_module_data_in[2] ;
 wire \sw_069_module_data_in[3] ;
 wire \sw_069_module_data_in[4] ;
 wire \sw_069_module_data_in[5] ;
 wire \sw_069_module_data_in[6] ;
 wire \sw_069_module_data_in[7] ;
 wire \sw_069_module_data_out[0] ;
 wire \sw_069_module_data_out[1] ;
 wire \sw_069_module_data_out[2] ;
 wire \sw_069_module_data_out[3] ;
 wire \sw_069_module_data_out[4] ;
 wire \sw_069_module_data_out[5] ;
 wire \sw_069_module_data_out[6] ;
 wire \sw_069_module_data_out[7] ;
 wire sw_069_scan_out;
 wire sw_070_clk_out;
 wire sw_070_data_out;
 wire sw_070_latch_out;
 wire \sw_070_module_data_in[0] ;
 wire \sw_070_module_data_in[1] ;
 wire \sw_070_module_data_in[2] ;
 wire \sw_070_module_data_in[3] ;
 wire \sw_070_module_data_in[4] ;
 wire \sw_070_module_data_in[5] ;
 wire \sw_070_module_data_in[6] ;
 wire \sw_070_module_data_in[7] ;
 wire \sw_070_module_data_out[0] ;
 wire \sw_070_module_data_out[1] ;
 wire \sw_070_module_data_out[2] ;
 wire \sw_070_module_data_out[3] ;
 wire \sw_070_module_data_out[4] ;
 wire \sw_070_module_data_out[5] ;
 wire \sw_070_module_data_out[6] ;
 wire \sw_070_module_data_out[7] ;
 wire sw_070_scan_out;
 wire sw_071_clk_out;
 wire sw_071_data_out;
 wire sw_071_latch_out;
 wire \sw_071_module_data_in[0] ;
 wire \sw_071_module_data_in[1] ;
 wire \sw_071_module_data_in[2] ;
 wire \sw_071_module_data_in[3] ;
 wire \sw_071_module_data_in[4] ;
 wire \sw_071_module_data_in[5] ;
 wire \sw_071_module_data_in[6] ;
 wire \sw_071_module_data_in[7] ;
 wire \sw_071_module_data_out[0] ;
 wire \sw_071_module_data_out[1] ;
 wire \sw_071_module_data_out[2] ;
 wire \sw_071_module_data_out[3] ;
 wire \sw_071_module_data_out[4] ;
 wire \sw_071_module_data_out[5] ;
 wire \sw_071_module_data_out[6] ;
 wire \sw_071_module_data_out[7] ;
 wire sw_071_scan_out;
 wire sw_072_clk_out;
 wire sw_072_data_out;
 wire sw_072_latch_out;
 wire \sw_072_module_data_in[0] ;
 wire \sw_072_module_data_in[1] ;
 wire \sw_072_module_data_in[2] ;
 wire \sw_072_module_data_in[3] ;
 wire \sw_072_module_data_in[4] ;
 wire \sw_072_module_data_in[5] ;
 wire \sw_072_module_data_in[6] ;
 wire \sw_072_module_data_in[7] ;
 wire \sw_072_module_data_out[0] ;
 wire \sw_072_module_data_out[1] ;
 wire \sw_072_module_data_out[2] ;
 wire \sw_072_module_data_out[3] ;
 wire \sw_072_module_data_out[4] ;
 wire \sw_072_module_data_out[5] ;
 wire \sw_072_module_data_out[6] ;
 wire \sw_072_module_data_out[7] ;
 wire sw_072_scan_out;
 wire sw_073_clk_out;
 wire sw_073_data_out;
 wire sw_073_latch_out;
 wire \sw_073_module_data_in[0] ;
 wire \sw_073_module_data_in[1] ;
 wire \sw_073_module_data_in[2] ;
 wire \sw_073_module_data_in[3] ;
 wire \sw_073_module_data_in[4] ;
 wire \sw_073_module_data_in[5] ;
 wire \sw_073_module_data_in[6] ;
 wire \sw_073_module_data_in[7] ;
 wire \sw_073_module_data_out[0] ;
 wire \sw_073_module_data_out[1] ;
 wire \sw_073_module_data_out[2] ;
 wire \sw_073_module_data_out[3] ;
 wire \sw_073_module_data_out[4] ;
 wire \sw_073_module_data_out[5] ;
 wire \sw_073_module_data_out[6] ;
 wire \sw_073_module_data_out[7] ;
 wire sw_073_scan_out;
 wire sw_074_clk_out;
 wire sw_074_data_out;
 wire sw_074_latch_out;
 wire \sw_074_module_data_in[0] ;
 wire \sw_074_module_data_in[1] ;
 wire \sw_074_module_data_in[2] ;
 wire \sw_074_module_data_in[3] ;
 wire \sw_074_module_data_in[4] ;
 wire \sw_074_module_data_in[5] ;
 wire \sw_074_module_data_in[6] ;
 wire \sw_074_module_data_in[7] ;
 wire \sw_074_module_data_out[0] ;
 wire \sw_074_module_data_out[1] ;
 wire \sw_074_module_data_out[2] ;
 wire \sw_074_module_data_out[3] ;
 wire \sw_074_module_data_out[4] ;
 wire \sw_074_module_data_out[5] ;
 wire \sw_074_module_data_out[6] ;
 wire \sw_074_module_data_out[7] ;
 wire sw_074_scan_out;
 wire sw_075_clk_out;
 wire sw_075_data_out;
 wire sw_075_latch_out;
 wire \sw_075_module_data_in[0] ;
 wire \sw_075_module_data_in[1] ;
 wire \sw_075_module_data_in[2] ;
 wire \sw_075_module_data_in[3] ;
 wire \sw_075_module_data_in[4] ;
 wire \sw_075_module_data_in[5] ;
 wire \sw_075_module_data_in[6] ;
 wire \sw_075_module_data_in[7] ;
 wire \sw_075_module_data_out[0] ;
 wire \sw_075_module_data_out[1] ;
 wire \sw_075_module_data_out[2] ;
 wire \sw_075_module_data_out[3] ;
 wire \sw_075_module_data_out[4] ;
 wire \sw_075_module_data_out[5] ;
 wire \sw_075_module_data_out[6] ;
 wire \sw_075_module_data_out[7] ;
 wire sw_075_scan_out;
 wire sw_076_clk_out;
 wire sw_076_data_out;
 wire sw_076_latch_out;
 wire \sw_076_module_data_in[0] ;
 wire \sw_076_module_data_in[1] ;
 wire \sw_076_module_data_in[2] ;
 wire \sw_076_module_data_in[3] ;
 wire \sw_076_module_data_in[4] ;
 wire \sw_076_module_data_in[5] ;
 wire \sw_076_module_data_in[6] ;
 wire \sw_076_module_data_in[7] ;
 wire \sw_076_module_data_out[0] ;
 wire \sw_076_module_data_out[1] ;
 wire \sw_076_module_data_out[2] ;
 wire \sw_076_module_data_out[3] ;
 wire \sw_076_module_data_out[4] ;
 wire \sw_076_module_data_out[5] ;
 wire \sw_076_module_data_out[6] ;
 wire \sw_076_module_data_out[7] ;
 wire sw_076_scan_out;
 wire sw_077_clk_out;
 wire sw_077_data_out;
 wire sw_077_latch_out;
 wire \sw_077_module_data_in[0] ;
 wire \sw_077_module_data_in[1] ;
 wire \sw_077_module_data_in[2] ;
 wire \sw_077_module_data_in[3] ;
 wire \sw_077_module_data_in[4] ;
 wire \sw_077_module_data_in[5] ;
 wire \sw_077_module_data_in[6] ;
 wire \sw_077_module_data_in[7] ;
 wire \sw_077_module_data_out[0] ;
 wire \sw_077_module_data_out[1] ;
 wire \sw_077_module_data_out[2] ;
 wire \sw_077_module_data_out[3] ;
 wire \sw_077_module_data_out[4] ;
 wire \sw_077_module_data_out[5] ;
 wire \sw_077_module_data_out[6] ;
 wire \sw_077_module_data_out[7] ;
 wire sw_077_scan_out;
 wire sw_078_clk_out;
 wire sw_078_data_out;
 wire sw_078_latch_out;
 wire \sw_078_module_data_in[0] ;
 wire \sw_078_module_data_in[1] ;
 wire \sw_078_module_data_in[2] ;
 wire \sw_078_module_data_in[3] ;
 wire \sw_078_module_data_in[4] ;
 wire \sw_078_module_data_in[5] ;
 wire \sw_078_module_data_in[6] ;
 wire \sw_078_module_data_in[7] ;
 wire \sw_078_module_data_out[0] ;
 wire \sw_078_module_data_out[1] ;
 wire \sw_078_module_data_out[2] ;
 wire \sw_078_module_data_out[3] ;
 wire \sw_078_module_data_out[4] ;
 wire \sw_078_module_data_out[5] ;
 wire \sw_078_module_data_out[6] ;
 wire \sw_078_module_data_out[7] ;
 wire sw_078_scan_out;
 wire sw_079_clk_out;
 wire sw_079_data_out;
 wire sw_079_latch_out;
 wire \sw_079_module_data_in[0] ;
 wire \sw_079_module_data_in[1] ;
 wire \sw_079_module_data_in[2] ;
 wire \sw_079_module_data_in[3] ;
 wire \sw_079_module_data_in[4] ;
 wire \sw_079_module_data_in[5] ;
 wire \sw_079_module_data_in[6] ;
 wire \sw_079_module_data_in[7] ;
 wire \sw_079_module_data_out[0] ;
 wire \sw_079_module_data_out[1] ;
 wire \sw_079_module_data_out[2] ;
 wire \sw_079_module_data_out[3] ;
 wire \sw_079_module_data_out[4] ;
 wire \sw_079_module_data_out[5] ;
 wire \sw_079_module_data_out[6] ;
 wire \sw_079_module_data_out[7] ;
 wire sw_079_scan_out;
 wire sw_080_clk_out;
 wire sw_080_data_out;
 wire sw_080_latch_out;
 wire \sw_080_module_data_in[0] ;
 wire \sw_080_module_data_in[1] ;
 wire \sw_080_module_data_in[2] ;
 wire \sw_080_module_data_in[3] ;
 wire \sw_080_module_data_in[4] ;
 wire \sw_080_module_data_in[5] ;
 wire \sw_080_module_data_in[6] ;
 wire \sw_080_module_data_in[7] ;
 wire \sw_080_module_data_out[0] ;
 wire \sw_080_module_data_out[1] ;
 wire \sw_080_module_data_out[2] ;
 wire \sw_080_module_data_out[3] ;
 wire \sw_080_module_data_out[4] ;
 wire \sw_080_module_data_out[5] ;
 wire \sw_080_module_data_out[6] ;
 wire \sw_080_module_data_out[7] ;
 wire sw_080_scan_out;
 wire sw_081_clk_out;
 wire sw_081_data_out;
 wire sw_081_latch_out;
 wire \sw_081_module_data_in[0] ;
 wire \sw_081_module_data_in[1] ;
 wire \sw_081_module_data_in[2] ;
 wire \sw_081_module_data_in[3] ;
 wire \sw_081_module_data_in[4] ;
 wire \sw_081_module_data_in[5] ;
 wire \sw_081_module_data_in[6] ;
 wire \sw_081_module_data_in[7] ;
 wire \sw_081_module_data_out[0] ;
 wire \sw_081_module_data_out[1] ;
 wire \sw_081_module_data_out[2] ;
 wire \sw_081_module_data_out[3] ;
 wire \sw_081_module_data_out[4] ;
 wire \sw_081_module_data_out[5] ;
 wire \sw_081_module_data_out[6] ;
 wire \sw_081_module_data_out[7] ;
 wire sw_081_scan_out;
 wire sw_082_clk_out;
 wire sw_082_data_out;
 wire sw_082_latch_out;
 wire \sw_082_module_data_in[0] ;
 wire \sw_082_module_data_in[1] ;
 wire \sw_082_module_data_in[2] ;
 wire \sw_082_module_data_in[3] ;
 wire \sw_082_module_data_in[4] ;
 wire \sw_082_module_data_in[5] ;
 wire \sw_082_module_data_in[6] ;
 wire \sw_082_module_data_in[7] ;
 wire \sw_082_module_data_out[0] ;
 wire \sw_082_module_data_out[1] ;
 wire \sw_082_module_data_out[2] ;
 wire \sw_082_module_data_out[3] ;
 wire \sw_082_module_data_out[4] ;
 wire \sw_082_module_data_out[5] ;
 wire \sw_082_module_data_out[6] ;
 wire \sw_082_module_data_out[7] ;
 wire sw_082_scan_out;
 wire sw_083_clk_out;
 wire sw_083_data_out;
 wire sw_083_latch_out;
 wire \sw_083_module_data_in[0] ;
 wire \sw_083_module_data_in[1] ;
 wire \sw_083_module_data_in[2] ;
 wire \sw_083_module_data_in[3] ;
 wire \sw_083_module_data_in[4] ;
 wire \sw_083_module_data_in[5] ;
 wire \sw_083_module_data_in[6] ;
 wire \sw_083_module_data_in[7] ;
 wire \sw_083_module_data_out[0] ;
 wire \sw_083_module_data_out[1] ;
 wire \sw_083_module_data_out[2] ;
 wire \sw_083_module_data_out[3] ;
 wire \sw_083_module_data_out[4] ;
 wire \sw_083_module_data_out[5] ;
 wire \sw_083_module_data_out[6] ;
 wire \sw_083_module_data_out[7] ;
 wire sw_083_scan_out;
 wire sw_084_clk_out;
 wire sw_084_data_out;
 wire sw_084_latch_out;
 wire \sw_084_module_data_in[0] ;
 wire \sw_084_module_data_in[1] ;
 wire \sw_084_module_data_in[2] ;
 wire \sw_084_module_data_in[3] ;
 wire \sw_084_module_data_in[4] ;
 wire \sw_084_module_data_in[5] ;
 wire \sw_084_module_data_in[6] ;
 wire \sw_084_module_data_in[7] ;
 wire \sw_084_module_data_out[0] ;
 wire \sw_084_module_data_out[1] ;
 wire \sw_084_module_data_out[2] ;
 wire \sw_084_module_data_out[3] ;
 wire \sw_084_module_data_out[4] ;
 wire \sw_084_module_data_out[5] ;
 wire \sw_084_module_data_out[6] ;
 wire \sw_084_module_data_out[7] ;
 wire sw_084_scan_out;
 wire sw_085_clk_out;
 wire sw_085_data_out;
 wire sw_085_latch_out;
 wire \sw_085_module_data_in[0] ;
 wire \sw_085_module_data_in[1] ;
 wire \sw_085_module_data_in[2] ;
 wire \sw_085_module_data_in[3] ;
 wire \sw_085_module_data_in[4] ;
 wire \sw_085_module_data_in[5] ;
 wire \sw_085_module_data_in[6] ;
 wire \sw_085_module_data_in[7] ;
 wire \sw_085_module_data_out[0] ;
 wire \sw_085_module_data_out[1] ;
 wire \sw_085_module_data_out[2] ;
 wire \sw_085_module_data_out[3] ;
 wire \sw_085_module_data_out[4] ;
 wire \sw_085_module_data_out[5] ;
 wire \sw_085_module_data_out[6] ;
 wire \sw_085_module_data_out[7] ;
 wire sw_085_scan_out;
 wire sw_086_clk_out;
 wire sw_086_data_out;
 wire sw_086_latch_out;
 wire \sw_086_module_data_in[0] ;
 wire \sw_086_module_data_in[1] ;
 wire \sw_086_module_data_in[2] ;
 wire \sw_086_module_data_in[3] ;
 wire \sw_086_module_data_in[4] ;
 wire \sw_086_module_data_in[5] ;
 wire \sw_086_module_data_in[6] ;
 wire \sw_086_module_data_in[7] ;
 wire \sw_086_module_data_out[0] ;
 wire \sw_086_module_data_out[1] ;
 wire \sw_086_module_data_out[2] ;
 wire \sw_086_module_data_out[3] ;
 wire \sw_086_module_data_out[4] ;
 wire \sw_086_module_data_out[5] ;
 wire \sw_086_module_data_out[6] ;
 wire \sw_086_module_data_out[7] ;
 wire sw_086_scan_out;
 wire sw_087_clk_out;
 wire sw_087_data_out;
 wire sw_087_latch_out;
 wire \sw_087_module_data_in[0] ;
 wire \sw_087_module_data_in[1] ;
 wire \sw_087_module_data_in[2] ;
 wire \sw_087_module_data_in[3] ;
 wire \sw_087_module_data_in[4] ;
 wire \sw_087_module_data_in[5] ;
 wire \sw_087_module_data_in[6] ;
 wire \sw_087_module_data_in[7] ;
 wire \sw_087_module_data_out[0] ;
 wire \sw_087_module_data_out[1] ;
 wire \sw_087_module_data_out[2] ;
 wire \sw_087_module_data_out[3] ;
 wire \sw_087_module_data_out[4] ;
 wire \sw_087_module_data_out[5] ;
 wire \sw_087_module_data_out[6] ;
 wire \sw_087_module_data_out[7] ;
 wire sw_087_scan_out;
 wire sw_088_clk_out;
 wire sw_088_data_out;
 wire sw_088_latch_out;
 wire \sw_088_module_data_in[0] ;
 wire \sw_088_module_data_in[1] ;
 wire \sw_088_module_data_in[2] ;
 wire \sw_088_module_data_in[3] ;
 wire \sw_088_module_data_in[4] ;
 wire \sw_088_module_data_in[5] ;
 wire \sw_088_module_data_in[6] ;
 wire \sw_088_module_data_in[7] ;
 wire \sw_088_module_data_out[0] ;
 wire \sw_088_module_data_out[1] ;
 wire \sw_088_module_data_out[2] ;
 wire \sw_088_module_data_out[3] ;
 wire \sw_088_module_data_out[4] ;
 wire \sw_088_module_data_out[5] ;
 wire \sw_088_module_data_out[6] ;
 wire \sw_088_module_data_out[7] ;
 wire sw_088_scan_out;
 wire sw_089_clk_out;
 wire sw_089_data_out;
 wire sw_089_latch_out;
 wire \sw_089_module_data_in[0] ;
 wire \sw_089_module_data_in[1] ;
 wire \sw_089_module_data_in[2] ;
 wire \sw_089_module_data_in[3] ;
 wire \sw_089_module_data_in[4] ;
 wire \sw_089_module_data_in[5] ;
 wire \sw_089_module_data_in[6] ;
 wire \sw_089_module_data_in[7] ;
 wire \sw_089_module_data_out[0] ;
 wire \sw_089_module_data_out[1] ;
 wire \sw_089_module_data_out[2] ;
 wire \sw_089_module_data_out[3] ;
 wire \sw_089_module_data_out[4] ;
 wire \sw_089_module_data_out[5] ;
 wire \sw_089_module_data_out[6] ;
 wire \sw_089_module_data_out[7] ;
 wire sw_089_scan_out;
 wire sw_090_clk_out;
 wire sw_090_data_out;
 wire sw_090_latch_out;
 wire \sw_090_module_data_in[0] ;
 wire \sw_090_module_data_in[1] ;
 wire \sw_090_module_data_in[2] ;
 wire \sw_090_module_data_in[3] ;
 wire \sw_090_module_data_in[4] ;
 wire \sw_090_module_data_in[5] ;
 wire \sw_090_module_data_in[6] ;
 wire \sw_090_module_data_in[7] ;
 wire \sw_090_module_data_out[0] ;
 wire \sw_090_module_data_out[1] ;
 wire \sw_090_module_data_out[2] ;
 wire \sw_090_module_data_out[3] ;
 wire \sw_090_module_data_out[4] ;
 wire \sw_090_module_data_out[5] ;
 wire \sw_090_module_data_out[6] ;
 wire \sw_090_module_data_out[7] ;
 wire sw_090_scan_out;
 wire sw_091_clk_out;
 wire sw_091_data_out;
 wire sw_091_latch_out;
 wire \sw_091_module_data_in[0] ;
 wire \sw_091_module_data_in[1] ;
 wire \sw_091_module_data_in[2] ;
 wire \sw_091_module_data_in[3] ;
 wire \sw_091_module_data_in[4] ;
 wire \sw_091_module_data_in[5] ;
 wire \sw_091_module_data_in[6] ;
 wire \sw_091_module_data_in[7] ;
 wire \sw_091_module_data_out[0] ;
 wire \sw_091_module_data_out[1] ;
 wire \sw_091_module_data_out[2] ;
 wire \sw_091_module_data_out[3] ;
 wire \sw_091_module_data_out[4] ;
 wire \sw_091_module_data_out[5] ;
 wire \sw_091_module_data_out[6] ;
 wire \sw_091_module_data_out[7] ;
 wire sw_091_scan_out;
 wire sw_092_clk_out;
 wire sw_092_data_out;
 wire sw_092_latch_out;
 wire \sw_092_module_data_in[0] ;
 wire \sw_092_module_data_in[1] ;
 wire \sw_092_module_data_in[2] ;
 wire \sw_092_module_data_in[3] ;
 wire \sw_092_module_data_in[4] ;
 wire \sw_092_module_data_in[5] ;
 wire \sw_092_module_data_in[6] ;
 wire \sw_092_module_data_in[7] ;
 wire \sw_092_module_data_out[0] ;
 wire \sw_092_module_data_out[1] ;
 wire \sw_092_module_data_out[2] ;
 wire \sw_092_module_data_out[3] ;
 wire \sw_092_module_data_out[4] ;
 wire \sw_092_module_data_out[5] ;
 wire \sw_092_module_data_out[6] ;
 wire \sw_092_module_data_out[7] ;
 wire sw_092_scan_out;
 wire sw_093_clk_out;
 wire sw_093_data_out;
 wire sw_093_latch_out;
 wire \sw_093_module_data_in[0] ;
 wire \sw_093_module_data_in[1] ;
 wire \sw_093_module_data_in[2] ;
 wire \sw_093_module_data_in[3] ;
 wire \sw_093_module_data_in[4] ;
 wire \sw_093_module_data_in[5] ;
 wire \sw_093_module_data_in[6] ;
 wire \sw_093_module_data_in[7] ;
 wire \sw_093_module_data_out[0] ;
 wire \sw_093_module_data_out[1] ;
 wire \sw_093_module_data_out[2] ;
 wire \sw_093_module_data_out[3] ;
 wire \sw_093_module_data_out[4] ;
 wire \sw_093_module_data_out[5] ;
 wire \sw_093_module_data_out[6] ;
 wire \sw_093_module_data_out[7] ;
 wire sw_093_scan_out;
 wire sw_094_clk_out;
 wire sw_094_data_out;
 wire sw_094_latch_out;
 wire \sw_094_module_data_in[0] ;
 wire \sw_094_module_data_in[1] ;
 wire \sw_094_module_data_in[2] ;
 wire \sw_094_module_data_in[3] ;
 wire \sw_094_module_data_in[4] ;
 wire \sw_094_module_data_in[5] ;
 wire \sw_094_module_data_in[6] ;
 wire \sw_094_module_data_in[7] ;
 wire \sw_094_module_data_out[0] ;
 wire \sw_094_module_data_out[1] ;
 wire \sw_094_module_data_out[2] ;
 wire \sw_094_module_data_out[3] ;
 wire \sw_094_module_data_out[4] ;
 wire \sw_094_module_data_out[5] ;
 wire \sw_094_module_data_out[6] ;
 wire \sw_094_module_data_out[7] ;
 wire sw_094_scan_out;
 wire sw_095_clk_out;
 wire sw_095_data_out;
 wire sw_095_latch_out;
 wire \sw_095_module_data_in[0] ;
 wire \sw_095_module_data_in[1] ;
 wire \sw_095_module_data_in[2] ;
 wire \sw_095_module_data_in[3] ;
 wire \sw_095_module_data_in[4] ;
 wire \sw_095_module_data_in[5] ;
 wire \sw_095_module_data_in[6] ;
 wire \sw_095_module_data_in[7] ;
 wire \sw_095_module_data_out[0] ;
 wire \sw_095_module_data_out[1] ;
 wire \sw_095_module_data_out[2] ;
 wire \sw_095_module_data_out[3] ;
 wire \sw_095_module_data_out[4] ;
 wire \sw_095_module_data_out[5] ;
 wire \sw_095_module_data_out[6] ;
 wire \sw_095_module_data_out[7] ;
 wire sw_095_scan_out;
 wire sw_096_clk_out;
 wire sw_096_data_out;
 wire sw_096_latch_out;
 wire \sw_096_module_data_in[0] ;
 wire \sw_096_module_data_in[1] ;
 wire \sw_096_module_data_in[2] ;
 wire \sw_096_module_data_in[3] ;
 wire \sw_096_module_data_in[4] ;
 wire \sw_096_module_data_in[5] ;
 wire \sw_096_module_data_in[6] ;
 wire \sw_096_module_data_in[7] ;
 wire \sw_096_module_data_out[0] ;
 wire \sw_096_module_data_out[1] ;
 wire \sw_096_module_data_out[2] ;
 wire \sw_096_module_data_out[3] ;
 wire \sw_096_module_data_out[4] ;
 wire \sw_096_module_data_out[5] ;
 wire \sw_096_module_data_out[6] ;
 wire \sw_096_module_data_out[7] ;
 wire sw_096_scan_out;
 wire sw_097_clk_out;
 wire sw_097_data_out;
 wire sw_097_latch_out;
 wire \sw_097_module_data_in[0] ;
 wire \sw_097_module_data_in[1] ;
 wire \sw_097_module_data_in[2] ;
 wire \sw_097_module_data_in[3] ;
 wire \sw_097_module_data_in[4] ;
 wire \sw_097_module_data_in[5] ;
 wire \sw_097_module_data_in[6] ;
 wire \sw_097_module_data_in[7] ;
 wire \sw_097_module_data_out[0] ;
 wire \sw_097_module_data_out[1] ;
 wire \sw_097_module_data_out[2] ;
 wire \sw_097_module_data_out[3] ;
 wire \sw_097_module_data_out[4] ;
 wire \sw_097_module_data_out[5] ;
 wire \sw_097_module_data_out[6] ;
 wire \sw_097_module_data_out[7] ;
 wire sw_097_scan_out;
 wire sw_098_clk_out;
 wire sw_098_data_out;
 wire sw_098_latch_out;
 wire \sw_098_module_data_in[0] ;
 wire \sw_098_module_data_in[1] ;
 wire \sw_098_module_data_in[2] ;
 wire \sw_098_module_data_in[3] ;
 wire \sw_098_module_data_in[4] ;
 wire \sw_098_module_data_in[5] ;
 wire \sw_098_module_data_in[6] ;
 wire \sw_098_module_data_in[7] ;
 wire \sw_098_module_data_out[0] ;
 wire \sw_098_module_data_out[1] ;
 wire \sw_098_module_data_out[2] ;
 wire \sw_098_module_data_out[3] ;
 wire \sw_098_module_data_out[4] ;
 wire \sw_098_module_data_out[5] ;
 wire \sw_098_module_data_out[6] ;
 wire \sw_098_module_data_out[7] ;
 wire sw_098_scan_out;
 wire sw_099_clk_out;
 wire sw_099_data_out;
 wire sw_099_latch_out;
 wire \sw_099_module_data_in[0] ;
 wire \sw_099_module_data_in[1] ;
 wire \sw_099_module_data_in[2] ;
 wire \sw_099_module_data_in[3] ;
 wire \sw_099_module_data_in[4] ;
 wire \sw_099_module_data_in[5] ;
 wire \sw_099_module_data_in[6] ;
 wire \sw_099_module_data_in[7] ;
 wire \sw_099_module_data_out[0] ;
 wire \sw_099_module_data_out[1] ;
 wire \sw_099_module_data_out[2] ;
 wire \sw_099_module_data_out[3] ;
 wire \sw_099_module_data_out[4] ;
 wire \sw_099_module_data_out[5] ;
 wire \sw_099_module_data_out[6] ;
 wire \sw_099_module_data_out[7] ;
 wire sw_099_scan_out;
 wire sw_100_clk_out;
 wire sw_100_data_out;
 wire sw_100_latch_out;
 wire \sw_100_module_data_in[0] ;
 wire \sw_100_module_data_in[1] ;
 wire \sw_100_module_data_in[2] ;
 wire \sw_100_module_data_in[3] ;
 wire \sw_100_module_data_in[4] ;
 wire \sw_100_module_data_in[5] ;
 wire \sw_100_module_data_in[6] ;
 wire \sw_100_module_data_in[7] ;
 wire \sw_100_module_data_out[0] ;
 wire \sw_100_module_data_out[1] ;
 wire \sw_100_module_data_out[2] ;
 wire \sw_100_module_data_out[3] ;
 wire \sw_100_module_data_out[4] ;
 wire \sw_100_module_data_out[5] ;
 wire \sw_100_module_data_out[6] ;
 wire \sw_100_module_data_out[7] ;
 wire sw_100_scan_out;
 wire sw_101_clk_out;
 wire sw_101_data_out;
 wire sw_101_latch_out;
 wire \sw_101_module_data_in[0] ;
 wire \sw_101_module_data_in[1] ;
 wire \sw_101_module_data_in[2] ;
 wire \sw_101_module_data_in[3] ;
 wire \sw_101_module_data_in[4] ;
 wire \sw_101_module_data_in[5] ;
 wire \sw_101_module_data_in[6] ;
 wire \sw_101_module_data_in[7] ;
 wire \sw_101_module_data_out[0] ;
 wire \sw_101_module_data_out[1] ;
 wire \sw_101_module_data_out[2] ;
 wire \sw_101_module_data_out[3] ;
 wire \sw_101_module_data_out[4] ;
 wire \sw_101_module_data_out[5] ;
 wire \sw_101_module_data_out[6] ;
 wire \sw_101_module_data_out[7] ;
 wire sw_101_scan_out;
 wire sw_102_clk_out;
 wire sw_102_data_out;
 wire sw_102_latch_out;
 wire \sw_102_module_data_in[0] ;
 wire \sw_102_module_data_in[1] ;
 wire \sw_102_module_data_in[2] ;
 wire \sw_102_module_data_in[3] ;
 wire \sw_102_module_data_in[4] ;
 wire \sw_102_module_data_in[5] ;
 wire \sw_102_module_data_in[6] ;
 wire \sw_102_module_data_in[7] ;
 wire \sw_102_module_data_out[0] ;
 wire \sw_102_module_data_out[1] ;
 wire \sw_102_module_data_out[2] ;
 wire \sw_102_module_data_out[3] ;
 wire \sw_102_module_data_out[4] ;
 wire \sw_102_module_data_out[5] ;
 wire \sw_102_module_data_out[6] ;
 wire \sw_102_module_data_out[7] ;
 wire sw_102_scan_out;
 wire sw_103_clk_out;
 wire sw_103_data_out;
 wire sw_103_latch_out;
 wire \sw_103_module_data_in[0] ;
 wire \sw_103_module_data_in[1] ;
 wire \sw_103_module_data_in[2] ;
 wire \sw_103_module_data_in[3] ;
 wire \sw_103_module_data_in[4] ;
 wire \sw_103_module_data_in[5] ;
 wire \sw_103_module_data_in[6] ;
 wire \sw_103_module_data_in[7] ;
 wire \sw_103_module_data_out[0] ;
 wire \sw_103_module_data_out[1] ;
 wire \sw_103_module_data_out[2] ;
 wire \sw_103_module_data_out[3] ;
 wire \sw_103_module_data_out[4] ;
 wire \sw_103_module_data_out[5] ;
 wire \sw_103_module_data_out[6] ;
 wire \sw_103_module_data_out[7] ;
 wire sw_103_scan_out;
 wire sw_104_clk_out;
 wire sw_104_data_out;
 wire sw_104_latch_out;
 wire \sw_104_module_data_in[0] ;
 wire \sw_104_module_data_in[1] ;
 wire \sw_104_module_data_in[2] ;
 wire \sw_104_module_data_in[3] ;
 wire \sw_104_module_data_in[4] ;
 wire \sw_104_module_data_in[5] ;
 wire \sw_104_module_data_in[6] ;
 wire \sw_104_module_data_in[7] ;
 wire \sw_104_module_data_out[0] ;
 wire \sw_104_module_data_out[1] ;
 wire \sw_104_module_data_out[2] ;
 wire \sw_104_module_data_out[3] ;
 wire \sw_104_module_data_out[4] ;
 wire \sw_104_module_data_out[5] ;
 wire \sw_104_module_data_out[6] ;
 wire \sw_104_module_data_out[7] ;
 wire sw_104_scan_out;
 wire sw_105_clk_out;
 wire sw_105_data_out;
 wire sw_105_latch_out;
 wire \sw_105_module_data_in[0] ;
 wire \sw_105_module_data_in[1] ;
 wire \sw_105_module_data_in[2] ;
 wire \sw_105_module_data_in[3] ;
 wire \sw_105_module_data_in[4] ;
 wire \sw_105_module_data_in[5] ;
 wire \sw_105_module_data_in[6] ;
 wire \sw_105_module_data_in[7] ;
 wire \sw_105_module_data_out[0] ;
 wire \sw_105_module_data_out[1] ;
 wire \sw_105_module_data_out[2] ;
 wire \sw_105_module_data_out[3] ;
 wire \sw_105_module_data_out[4] ;
 wire \sw_105_module_data_out[5] ;
 wire \sw_105_module_data_out[6] ;
 wire \sw_105_module_data_out[7] ;
 wire sw_105_scan_out;
 wire sw_106_clk_out;
 wire sw_106_data_out;
 wire sw_106_latch_out;
 wire \sw_106_module_data_in[0] ;
 wire \sw_106_module_data_in[1] ;
 wire \sw_106_module_data_in[2] ;
 wire \sw_106_module_data_in[3] ;
 wire \sw_106_module_data_in[4] ;
 wire \sw_106_module_data_in[5] ;
 wire \sw_106_module_data_in[6] ;
 wire \sw_106_module_data_in[7] ;
 wire \sw_106_module_data_out[0] ;
 wire \sw_106_module_data_out[1] ;
 wire \sw_106_module_data_out[2] ;
 wire \sw_106_module_data_out[3] ;
 wire \sw_106_module_data_out[4] ;
 wire \sw_106_module_data_out[5] ;
 wire \sw_106_module_data_out[6] ;
 wire \sw_106_module_data_out[7] ;
 wire sw_106_scan_out;
 wire sw_107_clk_out;
 wire sw_107_data_out;
 wire sw_107_latch_out;
 wire \sw_107_module_data_in[0] ;
 wire \sw_107_module_data_in[1] ;
 wire \sw_107_module_data_in[2] ;
 wire \sw_107_module_data_in[3] ;
 wire \sw_107_module_data_in[4] ;
 wire \sw_107_module_data_in[5] ;
 wire \sw_107_module_data_in[6] ;
 wire \sw_107_module_data_in[7] ;
 wire \sw_107_module_data_out[0] ;
 wire \sw_107_module_data_out[1] ;
 wire \sw_107_module_data_out[2] ;
 wire \sw_107_module_data_out[3] ;
 wire \sw_107_module_data_out[4] ;
 wire \sw_107_module_data_out[5] ;
 wire \sw_107_module_data_out[6] ;
 wire \sw_107_module_data_out[7] ;
 wire sw_107_scan_out;
 wire sw_108_clk_out;
 wire sw_108_data_out;
 wire sw_108_latch_out;
 wire \sw_108_module_data_in[0] ;
 wire \sw_108_module_data_in[1] ;
 wire \sw_108_module_data_in[2] ;
 wire \sw_108_module_data_in[3] ;
 wire \sw_108_module_data_in[4] ;
 wire \sw_108_module_data_in[5] ;
 wire \sw_108_module_data_in[6] ;
 wire \sw_108_module_data_in[7] ;
 wire \sw_108_module_data_out[0] ;
 wire \sw_108_module_data_out[1] ;
 wire \sw_108_module_data_out[2] ;
 wire \sw_108_module_data_out[3] ;
 wire \sw_108_module_data_out[4] ;
 wire \sw_108_module_data_out[5] ;
 wire \sw_108_module_data_out[6] ;
 wire \sw_108_module_data_out[7] ;
 wire sw_108_scan_out;
 wire sw_109_clk_out;
 wire sw_109_data_out;
 wire sw_109_latch_out;
 wire \sw_109_module_data_in[0] ;
 wire \sw_109_module_data_in[1] ;
 wire \sw_109_module_data_in[2] ;
 wire \sw_109_module_data_in[3] ;
 wire \sw_109_module_data_in[4] ;
 wire \sw_109_module_data_in[5] ;
 wire \sw_109_module_data_in[6] ;
 wire \sw_109_module_data_in[7] ;
 wire \sw_109_module_data_out[0] ;
 wire \sw_109_module_data_out[1] ;
 wire \sw_109_module_data_out[2] ;
 wire \sw_109_module_data_out[3] ;
 wire \sw_109_module_data_out[4] ;
 wire \sw_109_module_data_out[5] ;
 wire \sw_109_module_data_out[6] ;
 wire \sw_109_module_data_out[7] ;
 wire sw_109_scan_out;
 wire sw_110_clk_out;
 wire sw_110_data_out;
 wire sw_110_latch_out;
 wire \sw_110_module_data_in[0] ;
 wire \sw_110_module_data_in[1] ;
 wire \sw_110_module_data_in[2] ;
 wire \sw_110_module_data_in[3] ;
 wire \sw_110_module_data_in[4] ;
 wire \sw_110_module_data_in[5] ;
 wire \sw_110_module_data_in[6] ;
 wire \sw_110_module_data_in[7] ;
 wire \sw_110_module_data_out[0] ;
 wire \sw_110_module_data_out[1] ;
 wire \sw_110_module_data_out[2] ;
 wire \sw_110_module_data_out[3] ;
 wire \sw_110_module_data_out[4] ;
 wire \sw_110_module_data_out[5] ;
 wire \sw_110_module_data_out[6] ;
 wire \sw_110_module_data_out[7] ;
 wire sw_110_scan_out;
 wire sw_111_clk_out;
 wire sw_111_data_out;
 wire sw_111_latch_out;
 wire \sw_111_module_data_in[0] ;
 wire \sw_111_module_data_in[1] ;
 wire \sw_111_module_data_in[2] ;
 wire \sw_111_module_data_in[3] ;
 wire \sw_111_module_data_in[4] ;
 wire \sw_111_module_data_in[5] ;
 wire \sw_111_module_data_in[6] ;
 wire \sw_111_module_data_in[7] ;
 wire \sw_111_module_data_out[0] ;
 wire \sw_111_module_data_out[1] ;
 wire \sw_111_module_data_out[2] ;
 wire \sw_111_module_data_out[3] ;
 wire \sw_111_module_data_out[4] ;
 wire \sw_111_module_data_out[5] ;
 wire \sw_111_module_data_out[6] ;
 wire \sw_111_module_data_out[7] ;
 wire sw_111_scan_out;
 wire sw_112_clk_out;
 wire sw_112_data_out;
 wire sw_112_latch_out;
 wire \sw_112_module_data_in[0] ;
 wire \sw_112_module_data_in[1] ;
 wire \sw_112_module_data_in[2] ;
 wire \sw_112_module_data_in[3] ;
 wire \sw_112_module_data_in[4] ;
 wire \sw_112_module_data_in[5] ;
 wire \sw_112_module_data_in[6] ;
 wire \sw_112_module_data_in[7] ;
 wire \sw_112_module_data_out[0] ;
 wire \sw_112_module_data_out[1] ;
 wire \sw_112_module_data_out[2] ;
 wire \sw_112_module_data_out[3] ;
 wire \sw_112_module_data_out[4] ;
 wire \sw_112_module_data_out[5] ;
 wire \sw_112_module_data_out[6] ;
 wire \sw_112_module_data_out[7] ;
 wire sw_112_scan_out;
 wire sw_113_clk_out;
 wire sw_113_data_out;
 wire sw_113_latch_out;
 wire \sw_113_module_data_in[0] ;
 wire \sw_113_module_data_in[1] ;
 wire \sw_113_module_data_in[2] ;
 wire \sw_113_module_data_in[3] ;
 wire \sw_113_module_data_in[4] ;
 wire \sw_113_module_data_in[5] ;
 wire \sw_113_module_data_in[6] ;
 wire \sw_113_module_data_in[7] ;
 wire \sw_113_module_data_out[0] ;
 wire \sw_113_module_data_out[1] ;
 wire \sw_113_module_data_out[2] ;
 wire \sw_113_module_data_out[3] ;
 wire \sw_113_module_data_out[4] ;
 wire \sw_113_module_data_out[5] ;
 wire \sw_113_module_data_out[6] ;
 wire \sw_113_module_data_out[7] ;
 wire sw_113_scan_out;
 wire sw_114_clk_out;
 wire sw_114_data_out;
 wire sw_114_latch_out;
 wire \sw_114_module_data_in[0] ;
 wire \sw_114_module_data_in[1] ;
 wire \sw_114_module_data_in[2] ;
 wire \sw_114_module_data_in[3] ;
 wire \sw_114_module_data_in[4] ;
 wire \sw_114_module_data_in[5] ;
 wire \sw_114_module_data_in[6] ;
 wire \sw_114_module_data_in[7] ;
 wire \sw_114_module_data_out[0] ;
 wire \sw_114_module_data_out[1] ;
 wire \sw_114_module_data_out[2] ;
 wire \sw_114_module_data_out[3] ;
 wire \sw_114_module_data_out[4] ;
 wire \sw_114_module_data_out[5] ;
 wire \sw_114_module_data_out[6] ;
 wire \sw_114_module_data_out[7] ;
 wire sw_114_scan_out;
 wire sw_115_clk_out;
 wire sw_115_data_out;
 wire sw_115_latch_out;
 wire \sw_115_module_data_in[0] ;
 wire \sw_115_module_data_in[1] ;
 wire \sw_115_module_data_in[2] ;
 wire \sw_115_module_data_in[3] ;
 wire \sw_115_module_data_in[4] ;
 wire \sw_115_module_data_in[5] ;
 wire \sw_115_module_data_in[6] ;
 wire \sw_115_module_data_in[7] ;
 wire \sw_115_module_data_out[0] ;
 wire \sw_115_module_data_out[1] ;
 wire \sw_115_module_data_out[2] ;
 wire \sw_115_module_data_out[3] ;
 wire \sw_115_module_data_out[4] ;
 wire \sw_115_module_data_out[5] ;
 wire \sw_115_module_data_out[6] ;
 wire \sw_115_module_data_out[7] ;
 wire sw_115_scan_out;
 wire sw_116_clk_out;
 wire sw_116_data_out;
 wire sw_116_latch_out;
 wire \sw_116_module_data_in[0] ;
 wire \sw_116_module_data_in[1] ;
 wire \sw_116_module_data_in[2] ;
 wire \sw_116_module_data_in[3] ;
 wire \sw_116_module_data_in[4] ;
 wire \sw_116_module_data_in[5] ;
 wire \sw_116_module_data_in[6] ;
 wire \sw_116_module_data_in[7] ;
 wire \sw_116_module_data_out[0] ;
 wire \sw_116_module_data_out[1] ;
 wire \sw_116_module_data_out[2] ;
 wire \sw_116_module_data_out[3] ;
 wire \sw_116_module_data_out[4] ;
 wire \sw_116_module_data_out[5] ;
 wire \sw_116_module_data_out[6] ;
 wire \sw_116_module_data_out[7] ;
 wire sw_116_scan_out;
 wire sw_117_clk_out;
 wire sw_117_data_out;
 wire sw_117_latch_out;
 wire \sw_117_module_data_in[0] ;
 wire \sw_117_module_data_in[1] ;
 wire \sw_117_module_data_in[2] ;
 wire \sw_117_module_data_in[3] ;
 wire \sw_117_module_data_in[4] ;
 wire \sw_117_module_data_in[5] ;
 wire \sw_117_module_data_in[6] ;
 wire \sw_117_module_data_in[7] ;
 wire \sw_117_module_data_out[0] ;
 wire \sw_117_module_data_out[1] ;
 wire \sw_117_module_data_out[2] ;
 wire \sw_117_module_data_out[3] ;
 wire \sw_117_module_data_out[4] ;
 wire \sw_117_module_data_out[5] ;
 wire \sw_117_module_data_out[6] ;
 wire \sw_117_module_data_out[7] ;
 wire sw_117_scan_out;
 wire sw_118_clk_out;
 wire sw_118_data_out;
 wire sw_118_latch_out;
 wire \sw_118_module_data_in[0] ;
 wire \sw_118_module_data_in[1] ;
 wire \sw_118_module_data_in[2] ;
 wire \sw_118_module_data_in[3] ;
 wire \sw_118_module_data_in[4] ;
 wire \sw_118_module_data_in[5] ;
 wire \sw_118_module_data_in[6] ;
 wire \sw_118_module_data_in[7] ;
 wire \sw_118_module_data_out[0] ;
 wire \sw_118_module_data_out[1] ;
 wire \sw_118_module_data_out[2] ;
 wire \sw_118_module_data_out[3] ;
 wire \sw_118_module_data_out[4] ;
 wire \sw_118_module_data_out[5] ;
 wire \sw_118_module_data_out[6] ;
 wire \sw_118_module_data_out[7] ;
 wire sw_118_scan_out;
 wire sw_119_clk_out;
 wire sw_119_data_out;
 wire sw_119_latch_out;
 wire \sw_119_module_data_in[0] ;
 wire \sw_119_module_data_in[1] ;
 wire \sw_119_module_data_in[2] ;
 wire \sw_119_module_data_in[3] ;
 wire \sw_119_module_data_in[4] ;
 wire \sw_119_module_data_in[5] ;
 wire \sw_119_module_data_in[6] ;
 wire \sw_119_module_data_in[7] ;
 wire \sw_119_module_data_out[0] ;
 wire \sw_119_module_data_out[1] ;
 wire \sw_119_module_data_out[2] ;
 wire \sw_119_module_data_out[3] ;
 wire \sw_119_module_data_out[4] ;
 wire \sw_119_module_data_out[5] ;
 wire \sw_119_module_data_out[6] ;
 wire \sw_119_module_data_out[7] ;
 wire sw_119_scan_out;
 wire sw_120_clk_out;
 wire sw_120_data_out;
 wire sw_120_latch_out;
 wire \sw_120_module_data_in[0] ;
 wire \sw_120_module_data_in[1] ;
 wire \sw_120_module_data_in[2] ;
 wire \sw_120_module_data_in[3] ;
 wire \sw_120_module_data_in[4] ;
 wire \sw_120_module_data_in[5] ;
 wire \sw_120_module_data_in[6] ;
 wire \sw_120_module_data_in[7] ;
 wire \sw_120_module_data_out[0] ;
 wire \sw_120_module_data_out[1] ;
 wire \sw_120_module_data_out[2] ;
 wire \sw_120_module_data_out[3] ;
 wire \sw_120_module_data_out[4] ;
 wire \sw_120_module_data_out[5] ;
 wire \sw_120_module_data_out[6] ;
 wire \sw_120_module_data_out[7] ;
 wire sw_120_scan_out;
 wire sw_121_clk_out;
 wire sw_121_data_out;
 wire sw_121_latch_out;
 wire \sw_121_module_data_in[0] ;
 wire \sw_121_module_data_in[1] ;
 wire \sw_121_module_data_in[2] ;
 wire \sw_121_module_data_in[3] ;
 wire \sw_121_module_data_in[4] ;
 wire \sw_121_module_data_in[5] ;
 wire \sw_121_module_data_in[6] ;
 wire \sw_121_module_data_in[7] ;
 wire \sw_121_module_data_out[0] ;
 wire \sw_121_module_data_out[1] ;
 wire \sw_121_module_data_out[2] ;
 wire \sw_121_module_data_out[3] ;
 wire \sw_121_module_data_out[4] ;
 wire \sw_121_module_data_out[5] ;
 wire \sw_121_module_data_out[6] ;
 wire \sw_121_module_data_out[7] ;
 wire sw_121_scan_out;
 wire sw_122_clk_out;
 wire sw_122_data_out;
 wire sw_122_latch_out;
 wire \sw_122_module_data_in[0] ;
 wire \sw_122_module_data_in[1] ;
 wire \sw_122_module_data_in[2] ;
 wire \sw_122_module_data_in[3] ;
 wire \sw_122_module_data_in[4] ;
 wire \sw_122_module_data_in[5] ;
 wire \sw_122_module_data_in[6] ;
 wire \sw_122_module_data_in[7] ;
 wire \sw_122_module_data_out[0] ;
 wire \sw_122_module_data_out[1] ;
 wire \sw_122_module_data_out[2] ;
 wire \sw_122_module_data_out[3] ;
 wire \sw_122_module_data_out[4] ;
 wire \sw_122_module_data_out[5] ;
 wire \sw_122_module_data_out[6] ;
 wire \sw_122_module_data_out[7] ;
 wire sw_122_scan_out;
 wire sw_123_clk_out;
 wire sw_123_data_out;
 wire sw_123_latch_out;
 wire \sw_123_module_data_in[0] ;
 wire \sw_123_module_data_in[1] ;
 wire \sw_123_module_data_in[2] ;
 wire \sw_123_module_data_in[3] ;
 wire \sw_123_module_data_in[4] ;
 wire \sw_123_module_data_in[5] ;
 wire \sw_123_module_data_in[6] ;
 wire \sw_123_module_data_in[7] ;
 wire \sw_123_module_data_out[0] ;
 wire \sw_123_module_data_out[1] ;
 wire \sw_123_module_data_out[2] ;
 wire \sw_123_module_data_out[3] ;
 wire \sw_123_module_data_out[4] ;
 wire \sw_123_module_data_out[5] ;
 wire \sw_123_module_data_out[6] ;
 wire \sw_123_module_data_out[7] ;
 wire sw_123_scan_out;
 wire sw_124_clk_out;
 wire sw_124_data_out;
 wire sw_124_latch_out;
 wire \sw_124_module_data_in[0] ;
 wire \sw_124_module_data_in[1] ;
 wire \sw_124_module_data_in[2] ;
 wire \sw_124_module_data_in[3] ;
 wire \sw_124_module_data_in[4] ;
 wire \sw_124_module_data_in[5] ;
 wire \sw_124_module_data_in[6] ;
 wire \sw_124_module_data_in[7] ;
 wire \sw_124_module_data_out[0] ;
 wire \sw_124_module_data_out[1] ;
 wire \sw_124_module_data_out[2] ;
 wire \sw_124_module_data_out[3] ;
 wire \sw_124_module_data_out[4] ;
 wire \sw_124_module_data_out[5] ;
 wire \sw_124_module_data_out[6] ;
 wire \sw_124_module_data_out[7] ;
 wire sw_124_scan_out;
 wire sw_125_clk_out;
 wire sw_125_data_out;
 wire sw_125_latch_out;
 wire \sw_125_module_data_in[0] ;
 wire \sw_125_module_data_in[1] ;
 wire \sw_125_module_data_in[2] ;
 wire \sw_125_module_data_in[3] ;
 wire \sw_125_module_data_in[4] ;
 wire \sw_125_module_data_in[5] ;
 wire \sw_125_module_data_in[6] ;
 wire \sw_125_module_data_in[7] ;
 wire \sw_125_module_data_out[0] ;
 wire \sw_125_module_data_out[1] ;
 wire \sw_125_module_data_out[2] ;
 wire \sw_125_module_data_out[3] ;
 wire \sw_125_module_data_out[4] ;
 wire \sw_125_module_data_out[5] ;
 wire \sw_125_module_data_out[6] ;
 wire \sw_125_module_data_out[7] ;
 wire sw_125_scan_out;
 wire sw_126_clk_out;
 wire sw_126_data_out;
 wire sw_126_latch_out;
 wire \sw_126_module_data_in[0] ;
 wire \sw_126_module_data_in[1] ;
 wire \sw_126_module_data_in[2] ;
 wire \sw_126_module_data_in[3] ;
 wire \sw_126_module_data_in[4] ;
 wire \sw_126_module_data_in[5] ;
 wire \sw_126_module_data_in[6] ;
 wire \sw_126_module_data_in[7] ;
 wire \sw_126_module_data_out[0] ;
 wire \sw_126_module_data_out[1] ;
 wire \sw_126_module_data_out[2] ;
 wire \sw_126_module_data_out[3] ;
 wire \sw_126_module_data_out[4] ;
 wire \sw_126_module_data_out[5] ;
 wire \sw_126_module_data_out[6] ;
 wire \sw_126_module_data_out[7] ;
 wire sw_126_scan_out;
 wire sw_127_clk_out;
 wire sw_127_data_out;
 wire sw_127_latch_out;
 wire \sw_127_module_data_in[0] ;
 wire \sw_127_module_data_in[1] ;
 wire \sw_127_module_data_in[2] ;
 wire \sw_127_module_data_in[3] ;
 wire \sw_127_module_data_in[4] ;
 wire \sw_127_module_data_in[5] ;
 wire \sw_127_module_data_in[6] ;
 wire \sw_127_module_data_in[7] ;
 wire \sw_127_module_data_out[0] ;
 wire \sw_127_module_data_out[1] ;
 wire \sw_127_module_data_out[2] ;
 wire \sw_127_module_data_out[3] ;
 wire \sw_127_module_data_out[4] ;
 wire \sw_127_module_data_out[5] ;
 wire \sw_127_module_data_out[6] ;
 wire \sw_127_module_data_out[7] ;
 wire sw_127_scan_out;
 wire sw_128_clk_out;
 wire sw_128_data_out;
 wire sw_128_latch_out;
 wire \sw_128_module_data_in[0] ;
 wire \sw_128_module_data_in[1] ;
 wire \sw_128_module_data_in[2] ;
 wire \sw_128_module_data_in[3] ;
 wire \sw_128_module_data_in[4] ;
 wire \sw_128_module_data_in[5] ;
 wire \sw_128_module_data_in[6] ;
 wire \sw_128_module_data_in[7] ;
 wire \sw_128_module_data_out[0] ;
 wire \sw_128_module_data_out[1] ;
 wire \sw_128_module_data_out[2] ;
 wire \sw_128_module_data_out[3] ;
 wire \sw_128_module_data_out[4] ;
 wire \sw_128_module_data_out[5] ;
 wire \sw_128_module_data_out[6] ;
 wire \sw_128_module_data_out[7] ;
 wire sw_128_scan_out;
 wire sw_129_clk_out;
 wire sw_129_data_out;
 wire sw_129_latch_out;
 wire \sw_129_module_data_in[0] ;
 wire \sw_129_module_data_in[1] ;
 wire \sw_129_module_data_in[2] ;
 wire \sw_129_module_data_in[3] ;
 wire \sw_129_module_data_in[4] ;
 wire \sw_129_module_data_in[5] ;
 wire \sw_129_module_data_in[6] ;
 wire \sw_129_module_data_in[7] ;
 wire \sw_129_module_data_out[0] ;
 wire \sw_129_module_data_out[1] ;
 wire \sw_129_module_data_out[2] ;
 wire \sw_129_module_data_out[3] ;
 wire \sw_129_module_data_out[4] ;
 wire \sw_129_module_data_out[5] ;
 wire \sw_129_module_data_out[6] ;
 wire \sw_129_module_data_out[7] ;
 wire sw_129_scan_out;
 wire sw_130_clk_out;
 wire sw_130_data_out;
 wire sw_130_latch_out;
 wire \sw_130_module_data_in[0] ;
 wire \sw_130_module_data_in[1] ;
 wire \sw_130_module_data_in[2] ;
 wire \sw_130_module_data_in[3] ;
 wire \sw_130_module_data_in[4] ;
 wire \sw_130_module_data_in[5] ;
 wire \sw_130_module_data_in[6] ;
 wire \sw_130_module_data_in[7] ;
 wire \sw_130_module_data_out[0] ;
 wire \sw_130_module_data_out[1] ;
 wire \sw_130_module_data_out[2] ;
 wire \sw_130_module_data_out[3] ;
 wire \sw_130_module_data_out[4] ;
 wire \sw_130_module_data_out[5] ;
 wire \sw_130_module_data_out[6] ;
 wire \sw_130_module_data_out[7] ;
 wire sw_130_scan_out;
 wire sw_131_clk_out;
 wire sw_131_data_out;
 wire sw_131_latch_out;
 wire \sw_131_module_data_in[0] ;
 wire \sw_131_module_data_in[1] ;
 wire \sw_131_module_data_in[2] ;
 wire \sw_131_module_data_in[3] ;
 wire \sw_131_module_data_in[4] ;
 wire \sw_131_module_data_in[5] ;
 wire \sw_131_module_data_in[6] ;
 wire \sw_131_module_data_in[7] ;
 wire \sw_131_module_data_out[0] ;
 wire \sw_131_module_data_out[1] ;
 wire \sw_131_module_data_out[2] ;
 wire \sw_131_module_data_out[3] ;
 wire \sw_131_module_data_out[4] ;
 wire \sw_131_module_data_out[5] ;
 wire \sw_131_module_data_out[6] ;
 wire \sw_131_module_data_out[7] ;
 wire sw_131_scan_out;
 wire sw_132_clk_out;
 wire sw_132_data_out;
 wire sw_132_latch_out;
 wire \sw_132_module_data_in[0] ;
 wire \sw_132_module_data_in[1] ;
 wire \sw_132_module_data_in[2] ;
 wire \sw_132_module_data_in[3] ;
 wire \sw_132_module_data_in[4] ;
 wire \sw_132_module_data_in[5] ;
 wire \sw_132_module_data_in[6] ;
 wire \sw_132_module_data_in[7] ;
 wire \sw_132_module_data_out[0] ;
 wire \sw_132_module_data_out[1] ;
 wire \sw_132_module_data_out[2] ;
 wire \sw_132_module_data_out[3] ;
 wire \sw_132_module_data_out[4] ;
 wire \sw_132_module_data_out[5] ;
 wire \sw_132_module_data_out[6] ;
 wire \sw_132_module_data_out[7] ;
 wire sw_132_scan_out;
 wire sw_133_clk_out;
 wire sw_133_data_out;
 wire sw_133_latch_out;
 wire \sw_133_module_data_in[0] ;
 wire \sw_133_module_data_in[1] ;
 wire \sw_133_module_data_in[2] ;
 wire \sw_133_module_data_in[3] ;
 wire \sw_133_module_data_in[4] ;
 wire \sw_133_module_data_in[5] ;
 wire \sw_133_module_data_in[6] ;
 wire \sw_133_module_data_in[7] ;
 wire \sw_133_module_data_out[0] ;
 wire \sw_133_module_data_out[1] ;
 wire \sw_133_module_data_out[2] ;
 wire \sw_133_module_data_out[3] ;
 wire \sw_133_module_data_out[4] ;
 wire \sw_133_module_data_out[5] ;
 wire \sw_133_module_data_out[6] ;
 wire \sw_133_module_data_out[7] ;
 wire sw_133_scan_out;
 wire sw_134_clk_out;
 wire sw_134_data_out;
 wire sw_134_latch_out;
 wire \sw_134_module_data_in[0] ;
 wire \sw_134_module_data_in[1] ;
 wire \sw_134_module_data_in[2] ;
 wire \sw_134_module_data_in[3] ;
 wire \sw_134_module_data_in[4] ;
 wire \sw_134_module_data_in[5] ;
 wire \sw_134_module_data_in[6] ;
 wire \sw_134_module_data_in[7] ;
 wire \sw_134_module_data_out[0] ;
 wire \sw_134_module_data_out[1] ;
 wire \sw_134_module_data_out[2] ;
 wire \sw_134_module_data_out[3] ;
 wire \sw_134_module_data_out[4] ;
 wire \sw_134_module_data_out[5] ;
 wire \sw_134_module_data_out[6] ;
 wire \sw_134_module_data_out[7] ;
 wire sw_134_scan_out;
 wire sw_135_clk_out;
 wire sw_135_data_out;
 wire sw_135_latch_out;
 wire \sw_135_module_data_in[0] ;
 wire \sw_135_module_data_in[1] ;
 wire \sw_135_module_data_in[2] ;
 wire \sw_135_module_data_in[3] ;
 wire \sw_135_module_data_in[4] ;
 wire \sw_135_module_data_in[5] ;
 wire \sw_135_module_data_in[6] ;
 wire \sw_135_module_data_in[7] ;
 wire \sw_135_module_data_out[0] ;
 wire \sw_135_module_data_out[1] ;
 wire \sw_135_module_data_out[2] ;
 wire \sw_135_module_data_out[3] ;
 wire \sw_135_module_data_out[4] ;
 wire \sw_135_module_data_out[5] ;
 wire \sw_135_module_data_out[6] ;
 wire \sw_135_module_data_out[7] ;
 wire sw_135_scan_out;
 wire sw_136_clk_out;
 wire sw_136_data_out;
 wire sw_136_latch_out;
 wire \sw_136_module_data_in[0] ;
 wire \sw_136_module_data_in[1] ;
 wire \sw_136_module_data_in[2] ;
 wire \sw_136_module_data_in[3] ;
 wire \sw_136_module_data_in[4] ;
 wire \sw_136_module_data_in[5] ;
 wire \sw_136_module_data_in[6] ;
 wire \sw_136_module_data_in[7] ;
 wire \sw_136_module_data_out[0] ;
 wire \sw_136_module_data_out[1] ;
 wire \sw_136_module_data_out[2] ;
 wire \sw_136_module_data_out[3] ;
 wire \sw_136_module_data_out[4] ;
 wire \sw_136_module_data_out[5] ;
 wire \sw_136_module_data_out[6] ;
 wire \sw_136_module_data_out[7] ;
 wire sw_136_scan_out;
 wire sw_137_clk_out;
 wire sw_137_data_out;
 wire sw_137_latch_out;
 wire \sw_137_module_data_in[0] ;
 wire \sw_137_module_data_in[1] ;
 wire \sw_137_module_data_in[2] ;
 wire \sw_137_module_data_in[3] ;
 wire \sw_137_module_data_in[4] ;
 wire \sw_137_module_data_in[5] ;
 wire \sw_137_module_data_in[6] ;
 wire \sw_137_module_data_in[7] ;
 wire \sw_137_module_data_out[0] ;
 wire \sw_137_module_data_out[1] ;
 wire \sw_137_module_data_out[2] ;
 wire \sw_137_module_data_out[3] ;
 wire \sw_137_module_data_out[4] ;
 wire \sw_137_module_data_out[5] ;
 wire \sw_137_module_data_out[6] ;
 wire \sw_137_module_data_out[7] ;
 wire sw_137_scan_out;
 wire sw_138_clk_out;
 wire sw_138_data_out;
 wire sw_138_latch_out;
 wire \sw_138_module_data_in[0] ;
 wire \sw_138_module_data_in[1] ;
 wire \sw_138_module_data_in[2] ;
 wire \sw_138_module_data_in[3] ;
 wire \sw_138_module_data_in[4] ;
 wire \sw_138_module_data_in[5] ;
 wire \sw_138_module_data_in[6] ;
 wire \sw_138_module_data_in[7] ;
 wire \sw_138_module_data_out[0] ;
 wire \sw_138_module_data_out[1] ;
 wire \sw_138_module_data_out[2] ;
 wire \sw_138_module_data_out[3] ;
 wire \sw_138_module_data_out[4] ;
 wire \sw_138_module_data_out[5] ;
 wire \sw_138_module_data_out[6] ;
 wire \sw_138_module_data_out[7] ;
 wire sw_138_scan_out;
 wire sw_139_clk_out;
 wire sw_139_data_out;
 wire sw_139_latch_out;
 wire \sw_139_module_data_in[0] ;
 wire \sw_139_module_data_in[1] ;
 wire \sw_139_module_data_in[2] ;
 wire \sw_139_module_data_in[3] ;
 wire \sw_139_module_data_in[4] ;
 wire \sw_139_module_data_in[5] ;
 wire \sw_139_module_data_in[6] ;
 wire \sw_139_module_data_in[7] ;
 wire \sw_139_module_data_out[0] ;
 wire \sw_139_module_data_out[1] ;
 wire \sw_139_module_data_out[2] ;
 wire \sw_139_module_data_out[3] ;
 wire \sw_139_module_data_out[4] ;
 wire \sw_139_module_data_out[5] ;
 wire \sw_139_module_data_out[6] ;
 wire \sw_139_module_data_out[7] ;
 wire sw_139_scan_out;
 wire sw_140_clk_out;
 wire sw_140_data_out;
 wire sw_140_latch_out;
 wire \sw_140_module_data_in[0] ;
 wire \sw_140_module_data_in[1] ;
 wire \sw_140_module_data_in[2] ;
 wire \sw_140_module_data_in[3] ;
 wire \sw_140_module_data_in[4] ;
 wire \sw_140_module_data_in[5] ;
 wire \sw_140_module_data_in[6] ;
 wire \sw_140_module_data_in[7] ;
 wire \sw_140_module_data_out[0] ;
 wire \sw_140_module_data_out[1] ;
 wire \sw_140_module_data_out[2] ;
 wire \sw_140_module_data_out[3] ;
 wire \sw_140_module_data_out[4] ;
 wire \sw_140_module_data_out[5] ;
 wire \sw_140_module_data_out[6] ;
 wire \sw_140_module_data_out[7] ;
 wire sw_140_scan_out;
 wire sw_141_clk_out;
 wire sw_141_data_out;
 wire sw_141_latch_out;
 wire \sw_141_module_data_in[0] ;
 wire \sw_141_module_data_in[1] ;
 wire \sw_141_module_data_in[2] ;
 wire \sw_141_module_data_in[3] ;
 wire \sw_141_module_data_in[4] ;
 wire \sw_141_module_data_in[5] ;
 wire \sw_141_module_data_in[6] ;
 wire \sw_141_module_data_in[7] ;
 wire \sw_141_module_data_out[0] ;
 wire \sw_141_module_data_out[1] ;
 wire \sw_141_module_data_out[2] ;
 wire \sw_141_module_data_out[3] ;
 wire \sw_141_module_data_out[4] ;
 wire \sw_141_module_data_out[5] ;
 wire \sw_141_module_data_out[6] ;
 wire \sw_141_module_data_out[7] ;
 wire sw_141_scan_out;
 wire sw_142_clk_out;
 wire sw_142_data_out;
 wire sw_142_latch_out;
 wire \sw_142_module_data_in[0] ;
 wire \sw_142_module_data_in[1] ;
 wire \sw_142_module_data_in[2] ;
 wire \sw_142_module_data_in[3] ;
 wire \sw_142_module_data_in[4] ;
 wire \sw_142_module_data_in[5] ;
 wire \sw_142_module_data_in[6] ;
 wire \sw_142_module_data_in[7] ;
 wire \sw_142_module_data_out[0] ;
 wire \sw_142_module_data_out[1] ;
 wire \sw_142_module_data_out[2] ;
 wire \sw_142_module_data_out[3] ;
 wire \sw_142_module_data_out[4] ;
 wire \sw_142_module_data_out[5] ;
 wire \sw_142_module_data_out[6] ;
 wire \sw_142_module_data_out[7] ;
 wire sw_142_scan_out;
 wire sw_143_clk_out;
 wire sw_143_data_out;
 wire sw_143_latch_out;
 wire \sw_143_module_data_in[0] ;
 wire \sw_143_module_data_in[1] ;
 wire \sw_143_module_data_in[2] ;
 wire \sw_143_module_data_in[3] ;
 wire \sw_143_module_data_in[4] ;
 wire \sw_143_module_data_in[5] ;
 wire \sw_143_module_data_in[6] ;
 wire \sw_143_module_data_in[7] ;
 wire \sw_143_module_data_out[0] ;
 wire \sw_143_module_data_out[1] ;
 wire \sw_143_module_data_out[2] ;
 wire \sw_143_module_data_out[3] ;
 wire \sw_143_module_data_out[4] ;
 wire \sw_143_module_data_out[5] ;
 wire \sw_143_module_data_out[6] ;
 wire \sw_143_module_data_out[7] ;
 wire sw_143_scan_out;
 wire sw_144_clk_out;
 wire sw_144_data_out;
 wire sw_144_latch_out;
 wire \sw_144_module_data_in[0] ;
 wire \sw_144_module_data_in[1] ;
 wire \sw_144_module_data_in[2] ;
 wire \sw_144_module_data_in[3] ;
 wire \sw_144_module_data_in[4] ;
 wire \sw_144_module_data_in[5] ;
 wire \sw_144_module_data_in[6] ;
 wire \sw_144_module_data_in[7] ;
 wire \sw_144_module_data_out[0] ;
 wire \sw_144_module_data_out[1] ;
 wire \sw_144_module_data_out[2] ;
 wire \sw_144_module_data_out[3] ;
 wire \sw_144_module_data_out[4] ;
 wire \sw_144_module_data_out[5] ;
 wire \sw_144_module_data_out[6] ;
 wire \sw_144_module_data_out[7] ;
 wire sw_144_scan_out;
 wire sw_145_clk_out;
 wire sw_145_data_out;
 wire sw_145_latch_out;
 wire \sw_145_module_data_in[0] ;
 wire \sw_145_module_data_in[1] ;
 wire \sw_145_module_data_in[2] ;
 wire \sw_145_module_data_in[3] ;
 wire \sw_145_module_data_in[4] ;
 wire \sw_145_module_data_in[5] ;
 wire \sw_145_module_data_in[6] ;
 wire \sw_145_module_data_in[7] ;
 wire \sw_145_module_data_out[0] ;
 wire \sw_145_module_data_out[1] ;
 wire \sw_145_module_data_out[2] ;
 wire \sw_145_module_data_out[3] ;
 wire \sw_145_module_data_out[4] ;
 wire \sw_145_module_data_out[5] ;
 wire \sw_145_module_data_out[6] ;
 wire \sw_145_module_data_out[7] ;
 wire sw_145_scan_out;
 wire sw_146_clk_out;
 wire sw_146_data_out;
 wire sw_146_latch_out;
 wire \sw_146_module_data_in[0] ;
 wire \sw_146_module_data_in[1] ;
 wire \sw_146_module_data_in[2] ;
 wire \sw_146_module_data_in[3] ;
 wire \sw_146_module_data_in[4] ;
 wire \sw_146_module_data_in[5] ;
 wire \sw_146_module_data_in[6] ;
 wire \sw_146_module_data_in[7] ;
 wire \sw_146_module_data_out[0] ;
 wire \sw_146_module_data_out[1] ;
 wire \sw_146_module_data_out[2] ;
 wire \sw_146_module_data_out[3] ;
 wire \sw_146_module_data_out[4] ;
 wire \sw_146_module_data_out[5] ;
 wire \sw_146_module_data_out[6] ;
 wire \sw_146_module_data_out[7] ;
 wire sw_146_scan_out;
 wire sw_147_clk_out;
 wire sw_147_data_out;
 wire sw_147_latch_out;
 wire \sw_147_module_data_in[0] ;
 wire \sw_147_module_data_in[1] ;
 wire \sw_147_module_data_in[2] ;
 wire \sw_147_module_data_in[3] ;
 wire \sw_147_module_data_in[4] ;
 wire \sw_147_module_data_in[5] ;
 wire \sw_147_module_data_in[6] ;
 wire \sw_147_module_data_in[7] ;
 wire \sw_147_module_data_out[0] ;
 wire \sw_147_module_data_out[1] ;
 wire \sw_147_module_data_out[2] ;
 wire \sw_147_module_data_out[3] ;
 wire \sw_147_module_data_out[4] ;
 wire \sw_147_module_data_out[5] ;
 wire \sw_147_module_data_out[6] ;
 wire \sw_147_module_data_out[7] ;
 wire sw_147_scan_out;
 wire sw_148_clk_out;
 wire sw_148_data_out;
 wire sw_148_latch_out;
 wire \sw_148_module_data_in[0] ;
 wire \sw_148_module_data_in[1] ;
 wire \sw_148_module_data_in[2] ;
 wire \sw_148_module_data_in[3] ;
 wire \sw_148_module_data_in[4] ;
 wire \sw_148_module_data_in[5] ;
 wire \sw_148_module_data_in[6] ;
 wire \sw_148_module_data_in[7] ;
 wire \sw_148_module_data_out[0] ;
 wire \sw_148_module_data_out[1] ;
 wire \sw_148_module_data_out[2] ;
 wire \sw_148_module_data_out[3] ;
 wire \sw_148_module_data_out[4] ;
 wire \sw_148_module_data_out[5] ;
 wire \sw_148_module_data_out[6] ;
 wire \sw_148_module_data_out[7] ;
 wire sw_148_scan_out;
 wire sw_149_clk_out;
 wire sw_149_data_out;
 wire sw_149_latch_out;
 wire \sw_149_module_data_in[0] ;
 wire \sw_149_module_data_in[1] ;
 wire \sw_149_module_data_in[2] ;
 wire \sw_149_module_data_in[3] ;
 wire \sw_149_module_data_in[4] ;
 wire \sw_149_module_data_in[5] ;
 wire \sw_149_module_data_in[6] ;
 wire \sw_149_module_data_in[7] ;
 wire \sw_149_module_data_out[0] ;
 wire \sw_149_module_data_out[1] ;
 wire \sw_149_module_data_out[2] ;
 wire \sw_149_module_data_out[3] ;
 wire \sw_149_module_data_out[4] ;
 wire \sw_149_module_data_out[5] ;
 wire \sw_149_module_data_out[6] ;
 wire \sw_149_module_data_out[7] ;
 wire sw_149_scan_out;
 wire sw_150_clk_out;
 wire sw_150_data_out;
 wire sw_150_latch_out;
 wire \sw_150_module_data_in[0] ;
 wire \sw_150_module_data_in[1] ;
 wire \sw_150_module_data_in[2] ;
 wire \sw_150_module_data_in[3] ;
 wire \sw_150_module_data_in[4] ;
 wire \sw_150_module_data_in[5] ;
 wire \sw_150_module_data_in[6] ;
 wire \sw_150_module_data_in[7] ;
 wire \sw_150_module_data_out[0] ;
 wire \sw_150_module_data_out[1] ;
 wire \sw_150_module_data_out[2] ;
 wire \sw_150_module_data_out[3] ;
 wire \sw_150_module_data_out[4] ;
 wire \sw_150_module_data_out[5] ;
 wire \sw_150_module_data_out[6] ;
 wire \sw_150_module_data_out[7] ;
 wire sw_150_scan_out;
 wire sw_151_clk_out;
 wire sw_151_data_out;
 wire sw_151_latch_out;
 wire \sw_151_module_data_in[0] ;
 wire \sw_151_module_data_in[1] ;
 wire \sw_151_module_data_in[2] ;
 wire \sw_151_module_data_in[3] ;
 wire \sw_151_module_data_in[4] ;
 wire \sw_151_module_data_in[5] ;
 wire \sw_151_module_data_in[6] ;
 wire \sw_151_module_data_in[7] ;
 wire \sw_151_module_data_out[0] ;
 wire \sw_151_module_data_out[1] ;
 wire \sw_151_module_data_out[2] ;
 wire \sw_151_module_data_out[3] ;
 wire \sw_151_module_data_out[4] ;
 wire \sw_151_module_data_out[5] ;
 wire \sw_151_module_data_out[6] ;
 wire \sw_151_module_data_out[7] ;
 wire sw_151_scan_out;
 wire sw_152_clk_out;
 wire sw_152_data_out;
 wire sw_152_latch_out;
 wire \sw_152_module_data_in[0] ;
 wire \sw_152_module_data_in[1] ;
 wire \sw_152_module_data_in[2] ;
 wire \sw_152_module_data_in[3] ;
 wire \sw_152_module_data_in[4] ;
 wire \sw_152_module_data_in[5] ;
 wire \sw_152_module_data_in[6] ;
 wire \sw_152_module_data_in[7] ;
 wire \sw_152_module_data_out[0] ;
 wire \sw_152_module_data_out[1] ;
 wire \sw_152_module_data_out[2] ;
 wire \sw_152_module_data_out[3] ;
 wire \sw_152_module_data_out[4] ;
 wire \sw_152_module_data_out[5] ;
 wire \sw_152_module_data_out[6] ;
 wire \sw_152_module_data_out[7] ;
 wire sw_152_scan_out;
 wire sw_153_clk_out;
 wire sw_153_data_out;
 wire sw_153_latch_out;
 wire \sw_153_module_data_in[0] ;
 wire \sw_153_module_data_in[1] ;
 wire \sw_153_module_data_in[2] ;
 wire \sw_153_module_data_in[3] ;
 wire \sw_153_module_data_in[4] ;
 wire \sw_153_module_data_in[5] ;
 wire \sw_153_module_data_in[6] ;
 wire \sw_153_module_data_in[7] ;
 wire \sw_153_module_data_out[0] ;
 wire \sw_153_module_data_out[1] ;
 wire \sw_153_module_data_out[2] ;
 wire \sw_153_module_data_out[3] ;
 wire \sw_153_module_data_out[4] ;
 wire \sw_153_module_data_out[5] ;
 wire \sw_153_module_data_out[6] ;
 wire \sw_153_module_data_out[7] ;
 wire sw_153_scan_out;
 wire sw_154_clk_out;
 wire sw_154_data_out;
 wire sw_154_latch_out;
 wire \sw_154_module_data_in[0] ;
 wire \sw_154_module_data_in[1] ;
 wire \sw_154_module_data_in[2] ;
 wire \sw_154_module_data_in[3] ;
 wire \sw_154_module_data_in[4] ;
 wire \sw_154_module_data_in[5] ;
 wire \sw_154_module_data_in[6] ;
 wire \sw_154_module_data_in[7] ;
 wire \sw_154_module_data_out[0] ;
 wire \sw_154_module_data_out[1] ;
 wire \sw_154_module_data_out[2] ;
 wire \sw_154_module_data_out[3] ;
 wire \sw_154_module_data_out[4] ;
 wire \sw_154_module_data_out[5] ;
 wire \sw_154_module_data_out[6] ;
 wire \sw_154_module_data_out[7] ;
 wire sw_154_scan_out;
 wire sw_155_clk_out;
 wire sw_155_data_out;
 wire sw_155_latch_out;
 wire \sw_155_module_data_in[0] ;
 wire \sw_155_module_data_in[1] ;
 wire \sw_155_module_data_in[2] ;
 wire \sw_155_module_data_in[3] ;
 wire \sw_155_module_data_in[4] ;
 wire \sw_155_module_data_in[5] ;
 wire \sw_155_module_data_in[6] ;
 wire \sw_155_module_data_in[7] ;
 wire \sw_155_module_data_out[0] ;
 wire \sw_155_module_data_out[1] ;
 wire \sw_155_module_data_out[2] ;
 wire \sw_155_module_data_out[3] ;
 wire \sw_155_module_data_out[4] ;
 wire \sw_155_module_data_out[5] ;
 wire \sw_155_module_data_out[6] ;
 wire \sw_155_module_data_out[7] ;
 wire sw_155_scan_out;
 wire sw_156_clk_out;
 wire sw_156_data_out;
 wire sw_156_latch_out;
 wire \sw_156_module_data_in[0] ;
 wire \sw_156_module_data_in[1] ;
 wire \sw_156_module_data_in[2] ;
 wire \sw_156_module_data_in[3] ;
 wire \sw_156_module_data_in[4] ;
 wire \sw_156_module_data_in[5] ;
 wire \sw_156_module_data_in[6] ;
 wire \sw_156_module_data_in[7] ;
 wire \sw_156_module_data_out[0] ;
 wire \sw_156_module_data_out[1] ;
 wire \sw_156_module_data_out[2] ;
 wire \sw_156_module_data_out[3] ;
 wire \sw_156_module_data_out[4] ;
 wire \sw_156_module_data_out[5] ;
 wire \sw_156_module_data_out[6] ;
 wire \sw_156_module_data_out[7] ;
 wire sw_156_scan_out;
 wire sw_157_clk_out;
 wire sw_157_data_out;
 wire sw_157_latch_out;
 wire \sw_157_module_data_in[0] ;
 wire \sw_157_module_data_in[1] ;
 wire \sw_157_module_data_in[2] ;
 wire \sw_157_module_data_in[3] ;
 wire \sw_157_module_data_in[4] ;
 wire \sw_157_module_data_in[5] ;
 wire \sw_157_module_data_in[6] ;
 wire \sw_157_module_data_in[7] ;
 wire \sw_157_module_data_out[0] ;
 wire \sw_157_module_data_out[1] ;
 wire \sw_157_module_data_out[2] ;
 wire \sw_157_module_data_out[3] ;
 wire \sw_157_module_data_out[4] ;
 wire \sw_157_module_data_out[5] ;
 wire \sw_157_module_data_out[6] ;
 wire \sw_157_module_data_out[7] ;
 wire sw_157_scan_out;
 wire sw_158_clk_out;
 wire sw_158_data_out;
 wire sw_158_latch_out;
 wire \sw_158_module_data_in[0] ;
 wire \sw_158_module_data_in[1] ;
 wire \sw_158_module_data_in[2] ;
 wire \sw_158_module_data_in[3] ;
 wire \sw_158_module_data_in[4] ;
 wire \sw_158_module_data_in[5] ;
 wire \sw_158_module_data_in[6] ;
 wire \sw_158_module_data_in[7] ;
 wire \sw_158_module_data_out[0] ;
 wire \sw_158_module_data_out[1] ;
 wire \sw_158_module_data_out[2] ;
 wire \sw_158_module_data_out[3] ;
 wire \sw_158_module_data_out[4] ;
 wire \sw_158_module_data_out[5] ;
 wire \sw_158_module_data_out[6] ;
 wire \sw_158_module_data_out[7] ;
 wire sw_158_scan_out;
 wire sw_159_clk_out;
 wire sw_159_data_out;
 wire sw_159_latch_out;
 wire \sw_159_module_data_in[0] ;
 wire \sw_159_module_data_in[1] ;
 wire \sw_159_module_data_in[2] ;
 wire \sw_159_module_data_in[3] ;
 wire \sw_159_module_data_in[4] ;
 wire \sw_159_module_data_in[5] ;
 wire \sw_159_module_data_in[6] ;
 wire \sw_159_module_data_in[7] ;
 wire \sw_159_module_data_out[0] ;
 wire \sw_159_module_data_out[1] ;
 wire \sw_159_module_data_out[2] ;
 wire \sw_159_module_data_out[3] ;
 wire \sw_159_module_data_out[4] ;
 wire \sw_159_module_data_out[5] ;
 wire \sw_159_module_data_out[6] ;
 wire \sw_159_module_data_out[7] ;
 wire sw_159_scan_out;
 wire sw_160_clk_out;
 wire sw_160_data_out;
 wire sw_160_latch_out;
 wire \sw_160_module_data_in[0] ;
 wire \sw_160_module_data_in[1] ;
 wire \sw_160_module_data_in[2] ;
 wire \sw_160_module_data_in[3] ;
 wire \sw_160_module_data_in[4] ;
 wire \sw_160_module_data_in[5] ;
 wire \sw_160_module_data_in[6] ;
 wire \sw_160_module_data_in[7] ;
 wire \sw_160_module_data_out[0] ;
 wire \sw_160_module_data_out[1] ;
 wire \sw_160_module_data_out[2] ;
 wire \sw_160_module_data_out[3] ;
 wire \sw_160_module_data_out[4] ;
 wire \sw_160_module_data_out[5] ;
 wire \sw_160_module_data_out[6] ;
 wire \sw_160_module_data_out[7] ;
 wire sw_160_scan_out;
 wire sw_161_clk_out;
 wire sw_161_data_out;
 wire sw_161_latch_out;
 wire \sw_161_module_data_in[0] ;
 wire \sw_161_module_data_in[1] ;
 wire \sw_161_module_data_in[2] ;
 wire \sw_161_module_data_in[3] ;
 wire \sw_161_module_data_in[4] ;
 wire \sw_161_module_data_in[5] ;
 wire \sw_161_module_data_in[6] ;
 wire \sw_161_module_data_in[7] ;
 wire \sw_161_module_data_out[0] ;
 wire \sw_161_module_data_out[1] ;
 wire \sw_161_module_data_out[2] ;
 wire \sw_161_module_data_out[3] ;
 wire \sw_161_module_data_out[4] ;
 wire \sw_161_module_data_out[5] ;
 wire \sw_161_module_data_out[6] ;
 wire \sw_161_module_data_out[7] ;
 wire sw_161_scan_out;
 wire sw_162_clk_out;
 wire sw_162_data_out;
 wire sw_162_latch_out;
 wire \sw_162_module_data_in[0] ;
 wire \sw_162_module_data_in[1] ;
 wire \sw_162_module_data_in[2] ;
 wire \sw_162_module_data_in[3] ;
 wire \sw_162_module_data_in[4] ;
 wire \sw_162_module_data_in[5] ;
 wire \sw_162_module_data_in[6] ;
 wire \sw_162_module_data_in[7] ;
 wire \sw_162_module_data_out[0] ;
 wire \sw_162_module_data_out[1] ;
 wire \sw_162_module_data_out[2] ;
 wire \sw_162_module_data_out[3] ;
 wire \sw_162_module_data_out[4] ;
 wire \sw_162_module_data_out[5] ;
 wire \sw_162_module_data_out[6] ;
 wire \sw_162_module_data_out[7] ;
 wire sw_162_scan_out;
 wire sw_163_clk_out;
 wire sw_163_data_out;
 wire sw_163_latch_out;
 wire \sw_163_module_data_in[0] ;
 wire \sw_163_module_data_in[1] ;
 wire \sw_163_module_data_in[2] ;
 wire \sw_163_module_data_in[3] ;
 wire \sw_163_module_data_in[4] ;
 wire \sw_163_module_data_in[5] ;
 wire \sw_163_module_data_in[6] ;
 wire \sw_163_module_data_in[7] ;
 wire \sw_163_module_data_out[0] ;
 wire \sw_163_module_data_out[1] ;
 wire \sw_163_module_data_out[2] ;
 wire \sw_163_module_data_out[3] ;
 wire \sw_163_module_data_out[4] ;
 wire \sw_163_module_data_out[5] ;
 wire \sw_163_module_data_out[6] ;
 wire \sw_163_module_data_out[7] ;
 wire sw_163_scan_out;
 wire sw_164_clk_out;
 wire sw_164_data_out;
 wire sw_164_latch_out;
 wire \sw_164_module_data_in[0] ;
 wire \sw_164_module_data_in[1] ;
 wire \sw_164_module_data_in[2] ;
 wire \sw_164_module_data_in[3] ;
 wire \sw_164_module_data_in[4] ;
 wire \sw_164_module_data_in[5] ;
 wire \sw_164_module_data_in[6] ;
 wire \sw_164_module_data_in[7] ;
 wire \sw_164_module_data_out[0] ;
 wire \sw_164_module_data_out[1] ;
 wire \sw_164_module_data_out[2] ;
 wire \sw_164_module_data_out[3] ;
 wire \sw_164_module_data_out[4] ;
 wire \sw_164_module_data_out[5] ;
 wire \sw_164_module_data_out[6] ;
 wire \sw_164_module_data_out[7] ;
 wire sw_164_scan_out;
 wire sw_165_clk_out;
 wire sw_165_data_out;
 wire sw_165_latch_out;
 wire \sw_165_module_data_in[0] ;
 wire \sw_165_module_data_in[1] ;
 wire \sw_165_module_data_in[2] ;
 wire \sw_165_module_data_in[3] ;
 wire \sw_165_module_data_in[4] ;
 wire \sw_165_module_data_in[5] ;
 wire \sw_165_module_data_in[6] ;
 wire \sw_165_module_data_in[7] ;
 wire \sw_165_module_data_out[0] ;
 wire \sw_165_module_data_out[1] ;
 wire \sw_165_module_data_out[2] ;
 wire \sw_165_module_data_out[3] ;
 wire \sw_165_module_data_out[4] ;
 wire \sw_165_module_data_out[5] ;
 wire \sw_165_module_data_out[6] ;
 wire \sw_165_module_data_out[7] ;
 wire sw_165_scan_out;
 wire sw_166_clk_out;
 wire sw_166_data_out;
 wire sw_166_latch_out;
 wire \sw_166_module_data_in[0] ;
 wire \sw_166_module_data_in[1] ;
 wire \sw_166_module_data_in[2] ;
 wire \sw_166_module_data_in[3] ;
 wire \sw_166_module_data_in[4] ;
 wire \sw_166_module_data_in[5] ;
 wire \sw_166_module_data_in[6] ;
 wire \sw_166_module_data_in[7] ;
 wire \sw_166_module_data_out[0] ;
 wire \sw_166_module_data_out[1] ;
 wire \sw_166_module_data_out[2] ;
 wire \sw_166_module_data_out[3] ;
 wire \sw_166_module_data_out[4] ;
 wire \sw_166_module_data_out[5] ;
 wire \sw_166_module_data_out[6] ;
 wire \sw_166_module_data_out[7] ;
 wire sw_166_scan_out;
 wire sw_167_clk_out;
 wire sw_167_data_out;
 wire sw_167_latch_out;
 wire \sw_167_module_data_in[0] ;
 wire \sw_167_module_data_in[1] ;
 wire \sw_167_module_data_in[2] ;
 wire \sw_167_module_data_in[3] ;
 wire \sw_167_module_data_in[4] ;
 wire \sw_167_module_data_in[5] ;
 wire \sw_167_module_data_in[6] ;
 wire \sw_167_module_data_in[7] ;
 wire \sw_167_module_data_out[0] ;
 wire \sw_167_module_data_out[1] ;
 wire \sw_167_module_data_out[2] ;
 wire \sw_167_module_data_out[3] ;
 wire \sw_167_module_data_out[4] ;
 wire \sw_167_module_data_out[5] ;
 wire \sw_167_module_data_out[6] ;
 wire \sw_167_module_data_out[7] ;
 wire sw_167_scan_out;
 wire sw_168_clk_out;
 wire sw_168_data_out;
 wire sw_168_latch_out;
 wire \sw_168_module_data_in[0] ;
 wire \sw_168_module_data_in[1] ;
 wire \sw_168_module_data_in[2] ;
 wire \sw_168_module_data_in[3] ;
 wire \sw_168_module_data_in[4] ;
 wire \sw_168_module_data_in[5] ;
 wire \sw_168_module_data_in[6] ;
 wire \sw_168_module_data_in[7] ;
 wire \sw_168_module_data_out[0] ;
 wire \sw_168_module_data_out[1] ;
 wire \sw_168_module_data_out[2] ;
 wire \sw_168_module_data_out[3] ;
 wire \sw_168_module_data_out[4] ;
 wire \sw_168_module_data_out[5] ;
 wire \sw_168_module_data_out[6] ;
 wire \sw_168_module_data_out[7] ;
 wire sw_168_scan_out;
 wire sw_169_clk_out;
 wire sw_169_data_out;
 wire sw_169_latch_out;
 wire \sw_169_module_data_in[0] ;
 wire \sw_169_module_data_in[1] ;
 wire \sw_169_module_data_in[2] ;
 wire \sw_169_module_data_in[3] ;
 wire \sw_169_module_data_in[4] ;
 wire \sw_169_module_data_in[5] ;
 wire \sw_169_module_data_in[6] ;
 wire \sw_169_module_data_in[7] ;
 wire \sw_169_module_data_out[0] ;
 wire \sw_169_module_data_out[1] ;
 wire \sw_169_module_data_out[2] ;
 wire \sw_169_module_data_out[3] ;
 wire \sw_169_module_data_out[4] ;
 wire \sw_169_module_data_out[5] ;
 wire \sw_169_module_data_out[6] ;
 wire \sw_169_module_data_out[7] ;
 wire sw_169_scan_out;
 wire sw_170_clk_out;
 wire sw_170_data_out;
 wire sw_170_latch_out;
 wire \sw_170_module_data_in[0] ;
 wire \sw_170_module_data_in[1] ;
 wire \sw_170_module_data_in[2] ;
 wire \sw_170_module_data_in[3] ;
 wire \sw_170_module_data_in[4] ;
 wire \sw_170_module_data_in[5] ;
 wire \sw_170_module_data_in[6] ;
 wire \sw_170_module_data_in[7] ;
 wire \sw_170_module_data_out[0] ;
 wire \sw_170_module_data_out[1] ;
 wire \sw_170_module_data_out[2] ;
 wire \sw_170_module_data_out[3] ;
 wire \sw_170_module_data_out[4] ;
 wire \sw_170_module_data_out[5] ;
 wire \sw_170_module_data_out[6] ;
 wire \sw_170_module_data_out[7] ;
 wire sw_170_scan_out;
 wire sw_171_clk_out;
 wire sw_171_data_out;
 wire sw_171_latch_out;
 wire \sw_171_module_data_in[0] ;
 wire \sw_171_module_data_in[1] ;
 wire \sw_171_module_data_in[2] ;
 wire \sw_171_module_data_in[3] ;
 wire \sw_171_module_data_in[4] ;
 wire \sw_171_module_data_in[5] ;
 wire \sw_171_module_data_in[6] ;
 wire \sw_171_module_data_in[7] ;
 wire \sw_171_module_data_out[0] ;
 wire \sw_171_module_data_out[1] ;
 wire \sw_171_module_data_out[2] ;
 wire \sw_171_module_data_out[3] ;
 wire \sw_171_module_data_out[4] ;
 wire \sw_171_module_data_out[5] ;
 wire \sw_171_module_data_out[6] ;
 wire \sw_171_module_data_out[7] ;
 wire sw_171_scan_out;
 wire sw_172_clk_out;
 wire sw_172_data_out;
 wire sw_172_latch_out;
 wire \sw_172_module_data_in[0] ;
 wire \sw_172_module_data_in[1] ;
 wire \sw_172_module_data_in[2] ;
 wire \sw_172_module_data_in[3] ;
 wire \sw_172_module_data_in[4] ;
 wire \sw_172_module_data_in[5] ;
 wire \sw_172_module_data_in[6] ;
 wire \sw_172_module_data_in[7] ;
 wire \sw_172_module_data_out[0] ;
 wire \sw_172_module_data_out[1] ;
 wire \sw_172_module_data_out[2] ;
 wire \sw_172_module_data_out[3] ;
 wire \sw_172_module_data_out[4] ;
 wire \sw_172_module_data_out[5] ;
 wire \sw_172_module_data_out[6] ;
 wire \sw_172_module_data_out[7] ;
 wire sw_172_scan_out;
 wire sw_173_clk_out;
 wire sw_173_data_out;
 wire sw_173_latch_out;
 wire \sw_173_module_data_in[0] ;
 wire \sw_173_module_data_in[1] ;
 wire \sw_173_module_data_in[2] ;
 wire \sw_173_module_data_in[3] ;
 wire \sw_173_module_data_in[4] ;
 wire \sw_173_module_data_in[5] ;
 wire \sw_173_module_data_in[6] ;
 wire \sw_173_module_data_in[7] ;
 wire \sw_173_module_data_out[0] ;
 wire \sw_173_module_data_out[1] ;
 wire \sw_173_module_data_out[2] ;
 wire \sw_173_module_data_out[3] ;
 wire \sw_173_module_data_out[4] ;
 wire \sw_173_module_data_out[5] ;
 wire \sw_173_module_data_out[6] ;
 wire \sw_173_module_data_out[7] ;
 wire sw_173_scan_out;
 wire sw_174_clk_out;
 wire sw_174_data_out;
 wire sw_174_latch_out;
 wire \sw_174_module_data_in[0] ;
 wire \sw_174_module_data_in[1] ;
 wire \sw_174_module_data_in[2] ;
 wire \sw_174_module_data_in[3] ;
 wire \sw_174_module_data_in[4] ;
 wire \sw_174_module_data_in[5] ;
 wire \sw_174_module_data_in[6] ;
 wire \sw_174_module_data_in[7] ;
 wire \sw_174_module_data_out[0] ;
 wire \sw_174_module_data_out[1] ;
 wire \sw_174_module_data_out[2] ;
 wire \sw_174_module_data_out[3] ;
 wire \sw_174_module_data_out[4] ;
 wire \sw_174_module_data_out[5] ;
 wire \sw_174_module_data_out[6] ;
 wire \sw_174_module_data_out[7] ;
 wire sw_174_scan_out;
 wire sw_175_clk_out;
 wire sw_175_data_out;
 wire sw_175_latch_out;
 wire \sw_175_module_data_in[0] ;
 wire \sw_175_module_data_in[1] ;
 wire \sw_175_module_data_in[2] ;
 wire \sw_175_module_data_in[3] ;
 wire \sw_175_module_data_in[4] ;
 wire \sw_175_module_data_in[5] ;
 wire \sw_175_module_data_in[6] ;
 wire \sw_175_module_data_in[7] ;
 wire \sw_175_module_data_out[0] ;
 wire \sw_175_module_data_out[1] ;
 wire \sw_175_module_data_out[2] ;
 wire \sw_175_module_data_out[3] ;
 wire \sw_175_module_data_out[4] ;
 wire \sw_175_module_data_out[5] ;
 wire \sw_175_module_data_out[6] ;
 wire \sw_175_module_data_out[7] ;
 wire sw_175_scan_out;
 wire sw_176_clk_out;
 wire sw_176_data_out;
 wire sw_176_latch_out;
 wire \sw_176_module_data_in[0] ;
 wire \sw_176_module_data_in[1] ;
 wire \sw_176_module_data_in[2] ;
 wire \sw_176_module_data_in[3] ;
 wire \sw_176_module_data_in[4] ;
 wire \sw_176_module_data_in[5] ;
 wire \sw_176_module_data_in[6] ;
 wire \sw_176_module_data_in[7] ;
 wire \sw_176_module_data_out[0] ;
 wire \sw_176_module_data_out[1] ;
 wire \sw_176_module_data_out[2] ;
 wire \sw_176_module_data_out[3] ;
 wire \sw_176_module_data_out[4] ;
 wire \sw_176_module_data_out[5] ;
 wire \sw_176_module_data_out[6] ;
 wire \sw_176_module_data_out[7] ;
 wire sw_176_scan_out;
 wire sw_177_clk_out;
 wire sw_177_data_out;
 wire sw_177_latch_out;
 wire \sw_177_module_data_in[0] ;
 wire \sw_177_module_data_in[1] ;
 wire \sw_177_module_data_in[2] ;
 wire \sw_177_module_data_in[3] ;
 wire \sw_177_module_data_in[4] ;
 wire \sw_177_module_data_in[5] ;
 wire \sw_177_module_data_in[6] ;
 wire \sw_177_module_data_in[7] ;
 wire \sw_177_module_data_out[0] ;
 wire \sw_177_module_data_out[1] ;
 wire \sw_177_module_data_out[2] ;
 wire \sw_177_module_data_out[3] ;
 wire \sw_177_module_data_out[4] ;
 wire \sw_177_module_data_out[5] ;
 wire \sw_177_module_data_out[6] ;
 wire \sw_177_module_data_out[7] ;
 wire sw_177_scan_out;
 wire sw_178_clk_out;
 wire sw_178_data_out;
 wire sw_178_latch_out;
 wire \sw_178_module_data_in[0] ;
 wire \sw_178_module_data_in[1] ;
 wire \sw_178_module_data_in[2] ;
 wire \sw_178_module_data_in[3] ;
 wire \sw_178_module_data_in[4] ;
 wire \sw_178_module_data_in[5] ;
 wire \sw_178_module_data_in[6] ;
 wire \sw_178_module_data_in[7] ;
 wire \sw_178_module_data_out[0] ;
 wire \sw_178_module_data_out[1] ;
 wire \sw_178_module_data_out[2] ;
 wire \sw_178_module_data_out[3] ;
 wire \sw_178_module_data_out[4] ;
 wire \sw_178_module_data_out[5] ;
 wire \sw_178_module_data_out[6] ;
 wire \sw_178_module_data_out[7] ;
 wire sw_178_scan_out;
 wire sw_179_clk_out;
 wire sw_179_data_out;
 wire sw_179_latch_out;
 wire \sw_179_module_data_in[0] ;
 wire \sw_179_module_data_in[1] ;
 wire \sw_179_module_data_in[2] ;
 wire \sw_179_module_data_in[3] ;
 wire \sw_179_module_data_in[4] ;
 wire \sw_179_module_data_in[5] ;
 wire \sw_179_module_data_in[6] ;
 wire \sw_179_module_data_in[7] ;
 wire \sw_179_module_data_out[0] ;
 wire \sw_179_module_data_out[1] ;
 wire \sw_179_module_data_out[2] ;
 wire \sw_179_module_data_out[3] ;
 wire \sw_179_module_data_out[4] ;
 wire \sw_179_module_data_out[5] ;
 wire \sw_179_module_data_out[6] ;
 wire \sw_179_module_data_out[7] ;
 wire sw_179_scan_out;
 wire sw_180_clk_out;
 wire sw_180_data_out;
 wire sw_180_latch_out;
 wire \sw_180_module_data_in[0] ;
 wire \sw_180_module_data_in[1] ;
 wire \sw_180_module_data_in[2] ;
 wire \sw_180_module_data_in[3] ;
 wire \sw_180_module_data_in[4] ;
 wire \sw_180_module_data_in[5] ;
 wire \sw_180_module_data_in[6] ;
 wire \sw_180_module_data_in[7] ;
 wire \sw_180_module_data_out[0] ;
 wire \sw_180_module_data_out[1] ;
 wire \sw_180_module_data_out[2] ;
 wire \sw_180_module_data_out[3] ;
 wire \sw_180_module_data_out[4] ;
 wire \sw_180_module_data_out[5] ;
 wire \sw_180_module_data_out[6] ;
 wire \sw_180_module_data_out[7] ;
 wire sw_180_scan_out;
 wire sw_181_clk_out;
 wire sw_181_data_out;
 wire sw_181_latch_out;
 wire \sw_181_module_data_in[0] ;
 wire \sw_181_module_data_in[1] ;
 wire \sw_181_module_data_in[2] ;
 wire \sw_181_module_data_in[3] ;
 wire \sw_181_module_data_in[4] ;
 wire \sw_181_module_data_in[5] ;
 wire \sw_181_module_data_in[6] ;
 wire \sw_181_module_data_in[7] ;
 wire \sw_181_module_data_out[0] ;
 wire \sw_181_module_data_out[1] ;
 wire \sw_181_module_data_out[2] ;
 wire \sw_181_module_data_out[3] ;
 wire \sw_181_module_data_out[4] ;
 wire \sw_181_module_data_out[5] ;
 wire \sw_181_module_data_out[6] ;
 wire \sw_181_module_data_out[7] ;
 wire sw_181_scan_out;
 wire sw_182_clk_out;
 wire sw_182_data_out;
 wire sw_182_latch_out;
 wire \sw_182_module_data_in[0] ;
 wire \sw_182_module_data_in[1] ;
 wire \sw_182_module_data_in[2] ;
 wire \sw_182_module_data_in[3] ;
 wire \sw_182_module_data_in[4] ;
 wire \sw_182_module_data_in[5] ;
 wire \sw_182_module_data_in[6] ;
 wire \sw_182_module_data_in[7] ;
 wire \sw_182_module_data_out[0] ;
 wire \sw_182_module_data_out[1] ;
 wire \sw_182_module_data_out[2] ;
 wire \sw_182_module_data_out[3] ;
 wire \sw_182_module_data_out[4] ;
 wire \sw_182_module_data_out[5] ;
 wire \sw_182_module_data_out[6] ;
 wire \sw_182_module_data_out[7] ;
 wire sw_182_scan_out;
 wire sw_183_clk_out;
 wire sw_183_data_out;
 wire sw_183_latch_out;
 wire \sw_183_module_data_in[0] ;
 wire \sw_183_module_data_in[1] ;
 wire \sw_183_module_data_in[2] ;
 wire \sw_183_module_data_in[3] ;
 wire \sw_183_module_data_in[4] ;
 wire \sw_183_module_data_in[5] ;
 wire \sw_183_module_data_in[6] ;
 wire \sw_183_module_data_in[7] ;
 wire \sw_183_module_data_out[0] ;
 wire \sw_183_module_data_out[1] ;
 wire \sw_183_module_data_out[2] ;
 wire \sw_183_module_data_out[3] ;
 wire \sw_183_module_data_out[4] ;
 wire \sw_183_module_data_out[5] ;
 wire \sw_183_module_data_out[6] ;
 wire \sw_183_module_data_out[7] ;
 wire sw_183_scan_out;
 wire sw_184_clk_out;
 wire sw_184_data_out;
 wire sw_184_latch_out;
 wire \sw_184_module_data_in[0] ;
 wire \sw_184_module_data_in[1] ;
 wire \sw_184_module_data_in[2] ;
 wire \sw_184_module_data_in[3] ;
 wire \sw_184_module_data_in[4] ;
 wire \sw_184_module_data_in[5] ;
 wire \sw_184_module_data_in[6] ;
 wire \sw_184_module_data_in[7] ;
 wire \sw_184_module_data_out[0] ;
 wire \sw_184_module_data_out[1] ;
 wire \sw_184_module_data_out[2] ;
 wire \sw_184_module_data_out[3] ;
 wire \sw_184_module_data_out[4] ;
 wire \sw_184_module_data_out[5] ;
 wire \sw_184_module_data_out[6] ;
 wire \sw_184_module_data_out[7] ;
 wire sw_184_scan_out;
 wire sw_185_clk_out;
 wire sw_185_data_out;
 wire sw_185_latch_out;
 wire \sw_185_module_data_in[0] ;
 wire \sw_185_module_data_in[1] ;
 wire \sw_185_module_data_in[2] ;
 wire \sw_185_module_data_in[3] ;
 wire \sw_185_module_data_in[4] ;
 wire \sw_185_module_data_in[5] ;
 wire \sw_185_module_data_in[6] ;
 wire \sw_185_module_data_in[7] ;
 wire \sw_185_module_data_out[0] ;
 wire \sw_185_module_data_out[1] ;
 wire \sw_185_module_data_out[2] ;
 wire \sw_185_module_data_out[3] ;
 wire \sw_185_module_data_out[4] ;
 wire \sw_185_module_data_out[5] ;
 wire \sw_185_module_data_out[6] ;
 wire \sw_185_module_data_out[7] ;
 wire sw_185_scan_out;
 wire sw_186_clk_out;
 wire sw_186_data_out;
 wire sw_186_latch_out;
 wire \sw_186_module_data_in[0] ;
 wire \sw_186_module_data_in[1] ;
 wire \sw_186_module_data_in[2] ;
 wire \sw_186_module_data_in[3] ;
 wire \sw_186_module_data_in[4] ;
 wire \sw_186_module_data_in[5] ;
 wire \sw_186_module_data_in[6] ;
 wire \sw_186_module_data_in[7] ;
 wire \sw_186_module_data_out[0] ;
 wire \sw_186_module_data_out[1] ;
 wire \sw_186_module_data_out[2] ;
 wire \sw_186_module_data_out[3] ;
 wire \sw_186_module_data_out[4] ;
 wire \sw_186_module_data_out[5] ;
 wire \sw_186_module_data_out[6] ;
 wire \sw_186_module_data_out[7] ;
 wire sw_186_scan_out;
 wire sw_187_clk_out;
 wire sw_187_data_out;
 wire sw_187_latch_out;
 wire \sw_187_module_data_in[0] ;
 wire \sw_187_module_data_in[1] ;
 wire \sw_187_module_data_in[2] ;
 wire \sw_187_module_data_in[3] ;
 wire \sw_187_module_data_in[4] ;
 wire \sw_187_module_data_in[5] ;
 wire \sw_187_module_data_in[6] ;
 wire \sw_187_module_data_in[7] ;
 wire \sw_187_module_data_out[0] ;
 wire \sw_187_module_data_out[1] ;
 wire \sw_187_module_data_out[2] ;
 wire \sw_187_module_data_out[3] ;
 wire \sw_187_module_data_out[4] ;
 wire \sw_187_module_data_out[5] ;
 wire \sw_187_module_data_out[6] ;
 wire \sw_187_module_data_out[7] ;
 wire sw_187_scan_out;
 wire sw_188_clk_out;
 wire sw_188_data_out;
 wire sw_188_latch_out;
 wire \sw_188_module_data_in[0] ;
 wire \sw_188_module_data_in[1] ;
 wire \sw_188_module_data_in[2] ;
 wire \sw_188_module_data_in[3] ;
 wire \sw_188_module_data_in[4] ;
 wire \sw_188_module_data_in[5] ;
 wire \sw_188_module_data_in[6] ;
 wire \sw_188_module_data_in[7] ;
 wire \sw_188_module_data_out[0] ;
 wire \sw_188_module_data_out[1] ;
 wire \sw_188_module_data_out[2] ;
 wire \sw_188_module_data_out[3] ;
 wire \sw_188_module_data_out[4] ;
 wire \sw_188_module_data_out[5] ;
 wire \sw_188_module_data_out[6] ;
 wire \sw_188_module_data_out[7] ;
 wire sw_188_scan_out;
 wire sw_189_clk_out;
 wire sw_189_data_out;
 wire sw_189_latch_out;
 wire \sw_189_module_data_in[0] ;
 wire \sw_189_module_data_in[1] ;
 wire \sw_189_module_data_in[2] ;
 wire \sw_189_module_data_in[3] ;
 wire \sw_189_module_data_in[4] ;
 wire \sw_189_module_data_in[5] ;
 wire \sw_189_module_data_in[6] ;
 wire \sw_189_module_data_in[7] ;
 wire \sw_189_module_data_out[0] ;
 wire \sw_189_module_data_out[1] ;
 wire \sw_189_module_data_out[2] ;
 wire \sw_189_module_data_out[3] ;
 wire \sw_189_module_data_out[4] ;
 wire \sw_189_module_data_out[5] ;
 wire \sw_189_module_data_out[6] ;
 wire \sw_189_module_data_out[7] ;
 wire sw_189_scan_out;
 wire sw_190_clk_out;
 wire sw_190_data_out;
 wire sw_190_latch_out;
 wire \sw_190_module_data_in[0] ;
 wire \sw_190_module_data_in[1] ;
 wire \sw_190_module_data_in[2] ;
 wire \sw_190_module_data_in[3] ;
 wire \sw_190_module_data_in[4] ;
 wire \sw_190_module_data_in[5] ;
 wire \sw_190_module_data_in[6] ;
 wire \sw_190_module_data_in[7] ;
 wire \sw_190_module_data_out[0] ;
 wire \sw_190_module_data_out[1] ;
 wire \sw_190_module_data_out[2] ;
 wire \sw_190_module_data_out[3] ;
 wire \sw_190_module_data_out[4] ;
 wire \sw_190_module_data_out[5] ;
 wire \sw_190_module_data_out[6] ;
 wire \sw_190_module_data_out[7] ;
 wire sw_190_scan_out;
 wire sw_191_clk_out;
 wire sw_191_data_out;
 wire sw_191_latch_out;
 wire \sw_191_module_data_in[0] ;
 wire \sw_191_module_data_in[1] ;
 wire \sw_191_module_data_in[2] ;
 wire \sw_191_module_data_in[3] ;
 wire \sw_191_module_data_in[4] ;
 wire \sw_191_module_data_in[5] ;
 wire \sw_191_module_data_in[6] ;
 wire \sw_191_module_data_in[7] ;
 wire \sw_191_module_data_out[0] ;
 wire \sw_191_module_data_out[1] ;
 wire \sw_191_module_data_out[2] ;
 wire \sw_191_module_data_out[3] ;
 wire \sw_191_module_data_out[4] ;
 wire \sw_191_module_data_out[5] ;
 wire \sw_191_module_data_out[6] ;
 wire \sw_191_module_data_out[7] ;
 wire sw_191_scan_out;
 wire sw_192_clk_out;
 wire sw_192_data_out;
 wire sw_192_latch_out;
 wire \sw_192_module_data_in[0] ;
 wire \sw_192_module_data_in[1] ;
 wire \sw_192_module_data_in[2] ;
 wire \sw_192_module_data_in[3] ;
 wire \sw_192_module_data_in[4] ;
 wire \sw_192_module_data_in[5] ;
 wire \sw_192_module_data_in[6] ;
 wire \sw_192_module_data_in[7] ;
 wire \sw_192_module_data_out[0] ;
 wire \sw_192_module_data_out[1] ;
 wire \sw_192_module_data_out[2] ;
 wire \sw_192_module_data_out[3] ;
 wire \sw_192_module_data_out[4] ;
 wire \sw_192_module_data_out[5] ;
 wire \sw_192_module_data_out[6] ;
 wire \sw_192_module_data_out[7] ;
 wire sw_192_scan_out;
 wire sw_193_clk_out;
 wire sw_193_data_out;
 wire sw_193_latch_out;
 wire \sw_193_module_data_in[0] ;
 wire \sw_193_module_data_in[1] ;
 wire \sw_193_module_data_in[2] ;
 wire \sw_193_module_data_in[3] ;
 wire \sw_193_module_data_in[4] ;
 wire \sw_193_module_data_in[5] ;
 wire \sw_193_module_data_in[6] ;
 wire \sw_193_module_data_in[7] ;
 wire \sw_193_module_data_out[0] ;
 wire \sw_193_module_data_out[1] ;
 wire \sw_193_module_data_out[2] ;
 wire \sw_193_module_data_out[3] ;
 wire \sw_193_module_data_out[4] ;
 wire \sw_193_module_data_out[5] ;
 wire \sw_193_module_data_out[6] ;
 wire \sw_193_module_data_out[7] ;
 wire sw_193_scan_out;
 wire sw_194_clk_out;
 wire sw_194_data_out;
 wire sw_194_latch_out;
 wire \sw_194_module_data_in[0] ;
 wire \sw_194_module_data_in[1] ;
 wire \sw_194_module_data_in[2] ;
 wire \sw_194_module_data_in[3] ;
 wire \sw_194_module_data_in[4] ;
 wire \sw_194_module_data_in[5] ;
 wire \sw_194_module_data_in[6] ;
 wire \sw_194_module_data_in[7] ;
 wire \sw_194_module_data_out[0] ;
 wire \sw_194_module_data_out[1] ;
 wire \sw_194_module_data_out[2] ;
 wire \sw_194_module_data_out[3] ;
 wire \sw_194_module_data_out[4] ;
 wire \sw_194_module_data_out[5] ;
 wire \sw_194_module_data_out[6] ;
 wire \sw_194_module_data_out[7] ;
 wire sw_194_scan_out;
 wire sw_195_clk_out;
 wire sw_195_data_out;
 wire sw_195_latch_out;
 wire \sw_195_module_data_in[0] ;
 wire \sw_195_module_data_in[1] ;
 wire \sw_195_module_data_in[2] ;
 wire \sw_195_module_data_in[3] ;
 wire \sw_195_module_data_in[4] ;
 wire \sw_195_module_data_in[5] ;
 wire \sw_195_module_data_in[6] ;
 wire \sw_195_module_data_in[7] ;
 wire \sw_195_module_data_out[0] ;
 wire \sw_195_module_data_out[1] ;
 wire \sw_195_module_data_out[2] ;
 wire \sw_195_module_data_out[3] ;
 wire \sw_195_module_data_out[4] ;
 wire \sw_195_module_data_out[5] ;
 wire \sw_195_module_data_out[6] ;
 wire \sw_195_module_data_out[7] ;
 wire sw_195_scan_out;
 wire sw_196_clk_out;
 wire sw_196_data_out;
 wire sw_196_latch_out;
 wire \sw_196_module_data_in[0] ;
 wire \sw_196_module_data_in[1] ;
 wire \sw_196_module_data_in[2] ;
 wire \sw_196_module_data_in[3] ;
 wire \sw_196_module_data_in[4] ;
 wire \sw_196_module_data_in[5] ;
 wire \sw_196_module_data_in[6] ;
 wire \sw_196_module_data_in[7] ;
 wire \sw_196_module_data_out[0] ;
 wire \sw_196_module_data_out[1] ;
 wire \sw_196_module_data_out[2] ;
 wire \sw_196_module_data_out[3] ;
 wire \sw_196_module_data_out[4] ;
 wire \sw_196_module_data_out[5] ;
 wire \sw_196_module_data_out[6] ;
 wire \sw_196_module_data_out[7] ;
 wire sw_196_scan_out;
 wire sw_197_clk_out;
 wire sw_197_data_out;
 wire sw_197_latch_out;
 wire \sw_197_module_data_in[0] ;
 wire \sw_197_module_data_in[1] ;
 wire \sw_197_module_data_in[2] ;
 wire \sw_197_module_data_in[3] ;
 wire \sw_197_module_data_in[4] ;
 wire \sw_197_module_data_in[5] ;
 wire \sw_197_module_data_in[6] ;
 wire \sw_197_module_data_in[7] ;
 wire \sw_197_module_data_out[0] ;
 wire \sw_197_module_data_out[1] ;
 wire \sw_197_module_data_out[2] ;
 wire \sw_197_module_data_out[3] ;
 wire \sw_197_module_data_out[4] ;
 wire \sw_197_module_data_out[5] ;
 wire \sw_197_module_data_out[6] ;
 wire \sw_197_module_data_out[7] ;
 wire sw_197_scan_out;
 wire sw_198_clk_out;
 wire sw_198_data_out;
 wire sw_198_latch_out;
 wire \sw_198_module_data_in[0] ;
 wire \sw_198_module_data_in[1] ;
 wire \sw_198_module_data_in[2] ;
 wire \sw_198_module_data_in[3] ;
 wire \sw_198_module_data_in[4] ;
 wire \sw_198_module_data_in[5] ;
 wire \sw_198_module_data_in[6] ;
 wire \sw_198_module_data_in[7] ;
 wire \sw_198_module_data_out[0] ;
 wire \sw_198_module_data_out[1] ;
 wire \sw_198_module_data_out[2] ;
 wire \sw_198_module_data_out[3] ;
 wire \sw_198_module_data_out[4] ;
 wire \sw_198_module_data_out[5] ;
 wire \sw_198_module_data_out[6] ;
 wire \sw_198_module_data_out[7] ;
 wire sw_198_scan_out;
 wire sw_199_clk_out;
 wire sw_199_data_out;
 wire sw_199_latch_out;
 wire \sw_199_module_data_in[0] ;
 wire \sw_199_module_data_in[1] ;
 wire \sw_199_module_data_in[2] ;
 wire \sw_199_module_data_in[3] ;
 wire \sw_199_module_data_in[4] ;
 wire \sw_199_module_data_in[5] ;
 wire \sw_199_module_data_in[6] ;
 wire \sw_199_module_data_in[7] ;
 wire \sw_199_module_data_out[0] ;
 wire \sw_199_module_data_out[1] ;
 wire \sw_199_module_data_out[2] ;
 wire \sw_199_module_data_out[3] ;
 wire \sw_199_module_data_out[4] ;
 wire \sw_199_module_data_out[5] ;
 wire \sw_199_module_data_out[6] ;
 wire \sw_199_module_data_out[7] ;
 wire sw_199_scan_out;
 wire sw_200_clk_out;
 wire sw_200_data_out;
 wire sw_200_latch_out;
 wire \sw_200_module_data_in[0] ;
 wire \sw_200_module_data_in[1] ;
 wire \sw_200_module_data_in[2] ;
 wire \sw_200_module_data_in[3] ;
 wire \sw_200_module_data_in[4] ;
 wire \sw_200_module_data_in[5] ;
 wire \sw_200_module_data_in[6] ;
 wire \sw_200_module_data_in[7] ;
 wire \sw_200_module_data_out[0] ;
 wire \sw_200_module_data_out[1] ;
 wire \sw_200_module_data_out[2] ;
 wire \sw_200_module_data_out[3] ;
 wire \sw_200_module_data_out[4] ;
 wire \sw_200_module_data_out[5] ;
 wire \sw_200_module_data_out[6] ;
 wire \sw_200_module_data_out[7] ;
 wire sw_200_scan_out;
 wire sw_201_clk_out;
 wire sw_201_data_out;
 wire sw_201_latch_out;
 wire \sw_201_module_data_in[0] ;
 wire \sw_201_module_data_in[1] ;
 wire \sw_201_module_data_in[2] ;
 wire \sw_201_module_data_in[3] ;
 wire \sw_201_module_data_in[4] ;
 wire \sw_201_module_data_in[5] ;
 wire \sw_201_module_data_in[6] ;
 wire \sw_201_module_data_in[7] ;
 wire \sw_201_module_data_out[0] ;
 wire \sw_201_module_data_out[1] ;
 wire \sw_201_module_data_out[2] ;
 wire \sw_201_module_data_out[3] ;
 wire \sw_201_module_data_out[4] ;
 wire \sw_201_module_data_out[5] ;
 wire \sw_201_module_data_out[6] ;
 wire \sw_201_module_data_out[7] ;
 wire sw_201_scan_out;
 wire sw_202_clk_out;
 wire sw_202_data_out;
 wire sw_202_latch_out;
 wire \sw_202_module_data_in[0] ;
 wire \sw_202_module_data_in[1] ;
 wire \sw_202_module_data_in[2] ;
 wire \sw_202_module_data_in[3] ;
 wire \sw_202_module_data_in[4] ;
 wire \sw_202_module_data_in[5] ;
 wire \sw_202_module_data_in[6] ;
 wire \sw_202_module_data_in[7] ;
 wire \sw_202_module_data_out[0] ;
 wire \sw_202_module_data_out[1] ;
 wire \sw_202_module_data_out[2] ;
 wire \sw_202_module_data_out[3] ;
 wire \sw_202_module_data_out[4] ;
 wire \sw_202_module_data_out[5] ;
 wire \sw_202_module_data_out[6] ;
 wire \sw_202_module_data_out[7] ;
 wire sw_202_scan_out;
 wire sw_203_clk_out;
 wire sw_203_data_out;
 wire sw_203_latch_out;
 wire \sw_203_module_data_in[0] ;
 wire \sw_203_module_data_in[1] ;
 wire \sw_203_module_data_in[2] ;
 wire \sw_203_module_data_in[3] ;
 wire \sw_203_module_data_in[4] ;
 wire \sw_203_module_data_in[5] ;
 wire \sw_203_module_data_in[6] ;
 wire \sw_203_module_data_in[7] ;
 wire \sw_203_module_data_out[0] ;
 wire \sw_203_module_data_out[1] ;
 wire \sw_203_module_data_out[2] ;
 wire \sw_203_module_data_out[3] ;
 wire \sw_203_module_data_out[4] ;
 wire \sw_203_module_data_out[5] ;
 wire \sw_203_module_data_out[6] ;
 wire \sw_203_module_data_out[7] ;
 wire sw_203_scan_out;
 wire sw_204_clk_out;
 wire sw_204_data_out;
 wire sw_204_latch_out;
 wire \sw_204_module_data_in[0] ;
 wire \sw_204_module_data_in[1] ;
 wire \sw_204_module_data_in[2] ;
 wire \sw_204_module_data_in[3] ;
 wire \sw_204_module_data_in[4] ;
 wire \sw_204_module_data_in[5] ;
 wire \sw_204_module_data_in[6] ;
 wire \sw_204_module_data_in[7] ;
 wire \sw_204_module_data_out[0] ;
 wire \sw_204_module_data_out[1] ;
 wire \sw_204_module_data_out[2] ;
 wire \sw_204_module_data_out[3] ;
 wire \sw_204_module_data_out[4] ;
 wire \sw_204_module_data_out[5] ;
 wire \sw_204_module_data_out[6] ;
 wire \sw_204_module_data_out[7] ;
 wire sw_204_scan_out;
 wire sw_205_clk_out;
 wire sw_205_data_out;
 wire sw_205_latch_out;
 wire \sw_205_module_data_in[0] ;
 wire \sw_205_module_data_in[1] ;
 wire \sw_205_module_data_in[2] ;
 wire \sw_205_module_data_in[3] ;
 wire \sw_205_module_data_in[4] ;
 wire \sw_205_module_data_in[5] ;
 wire \sw_205_module_data_in[6] ;
 wire \sw_205_module_data_in[7] ;
 wire \sw_205_module_data_out[0] ;
 wire \sw_205_module_data_out[1] ;
 wire \sw_205_module_data_out[2] ;
 wire \sw_205_module_data_out[3] ;
 wire \sw_205_module_data_out[4] ;
 wire \sw_205_module_data_out[5] ;
 wire \sw_205_module_data_out[6] ;
 wire \sw_205_module_data_out[7] ;
 wire sw_205_scan_out;
 wire sw_206_clk_out;
 wire sw_206_data_out;
 wire sw_206_latch_out;
 wire \sw_206_module_data_in[0] ;
 wire \sw_206_module_data_in[1] ;
 wire \sw_206_module_data_in[2] ;
 wire \sw_206_module_data_in[3] ;
 wire \sw_206_module_data_in[4] ;
 wire \sw_206_module_data_in[5] ;
 wire \sw_206_module_data_in[6] ;
 wire \sw_206_module_data_in[7] ;
 wire \sw_206_module_data_out[0] ;
 wire \sw_206_module_data_out[1] ;
 wire \sw_206_module_data_out[2] ;
 wire \sw_206_module_data_out[3] ;
 wire \sw_206_module_data_out[4] ;
 wire \sw_206_module_data_out[5] ;
 wire \sw_206_module_data_out[6] ;
 wire \sw_206_module_data_out[7] ;
 wire sw_206_scan_out;
 wire sw_207_clk_out;
 wire sw_207_data_out;
 wire sw_207_latch_out;
 wire \sw_207_module_data_in[0] ;
 wire \sw_207_module_data_in[1] ;
 wire \sw_207_module_data_in[2] ;
 wire \sw_207_module_data_in[3] ;
 wire \sw_207_module_data_in[4] ;
 wire \sw_207_module_data_in[5] ;
 wire \sw_207_module_data_in[6] ;
 wire \sw_207_module_data_in[7] ;
 wire \sw_207_module_data_out[0] ;
 wire \sw_207_module_data_out[1] ;
 wire \sw_207_module_data_out[2] ;
 wire \sw_207_module_data_out[3] ;
 wire \sw_207_module_data_out[4] ;
 wire \sw_207_module_data_out[5] ;
 wire \sw_207_module_data_out[6] ;
 wire \sw_207_module_data_out[7] ;
 wire sw_207_scan_out;
 wire sw_208_clk_out;
 wire sw_208_data_out;
 wire sw_208_latch_out;
 wire \sw_208_module_data_in[0] ;
 wire \sw_208_module_data_in[1] ;
 wire \sw_208_module_data_in[2] ;
 wire \sw_208_module_data_in[3] ;
 wire \sw_208_module_data_in[4] ;
 wire \sw_208_module_data_in[5] ;
 wire \sw_208_module_data_in[6] ;
 wire \sw_208_module_data_in[7] ;
 wire \sw_208_module_data_out[0] ;
 wire \sw_208_module_data_out[1] ;
 wire \sw_208_module_data_out[2] ;
 wire \sw_208_module_data_out[3] ;
 wire \sw_208_module_data_out[4] ;
 wire \sw_208_module_data_out[5] ;
 wire \sw_208_module_data_out[6] ;
 wire \sw_208_module_data_out[7] ;
 wire sw_208_scan_out;
 wire sw_209_clk_out;
 wire sw_209_data_out;
 wire sw_209_latch_out;
 wire \sw_209_module_data_in[0] ;
 wire \sw_209_module_data_in[1] ;
 wire \sw_209_module_data_in[2] ;
 wire \sw_209_module_data_in[3] ;
 wire \sw_209_module_data_in[4] ;
 wire \sw_209_module_data_in[5] ;
 wire \sw_209_module_data_in[6] ;
 wire \sw_209_module_data_in[7] ;
 wire \sw_209_module_data_out[0] ;
 wire \sw_209_module_data_out[1] ;
 wire \sw_209_module_data_out[2] ;
 wire \sw_209_module_data_out[3] ;
 wire \sw_209_module_data_out[4] ;
 wire \sw_209_module_data_out[5] ;
 wire \sw_209_module_data_out[6] ;
 wire \sw_209_module_data_out[7] ;
 wire sw_209_scan_out;
 wire sw_210_clk_out;
 wire sw_210_data_out;
 wire sw_210_latch_out;
 wire \sw_210_module_data_in[0] ;
 wire \sw_210_module_data_in[1] ;
 wire \sw_210_module_data_in[2] ;
 wire \sw_210_module_data_in[3] ;
 wire \sw_210_module_data_in[4] ;
 wire \sw_210_module_data_in[5] ;
 wire \sw_210_module_data_in[6] ;
 wire \sw_210_module_data_in[7] ;
 wire \sw_210_module_data_out[0] ;
 wire \sw_210_module_data_out[1] ;
 wire \sw_210_module_data_out[2] ;
 wire \sw_210_module_data_out[3] ;
 wire \sw_210_module_data_out[4] ;
 wire \sw_210_module_data_out[5] ;
 wire \sw_210_module_data_out[6] ;
 wire \sw_210_module_data_out[7] ;
 wire sw_210_scan_out;
 wire sw_211_clk_out;
 wire sw_211_data_out;
 wire sw_211_latch_out;
 wire \sw_211_module_data_in[0] ;
 wire \sw_211_module_data_in[1] ;
 wire \sw_211_module_data_in[2] ;
 wire \sw_211_module_data_in[3] ;
 wire \sw_211_module_data_in[4] ;
 wire \sw_211_module_data_in[5] ;
 wire \sw_211_module_data_in[6] ;
 wire \sw_211_module_data_in[7] ;
 wire \sw_211_module_data_out[0] ;
 wire \sw_211_module_data_out[1] ;
 wire \sw_211_module_data_out[2] ;
 wire \sw_211_module_data_out[3] ;
 wire \sw_211_module_data_out[4] ;
 wire \sw_211_module_data_out[5] ;
 wire \sw_211_module_data_out[6] ;
 wire \sw_211_module_data_out[7] ;
 wire sw_211_scan_out;
 wire sw_212_clk_out;
 wire sw_212_data_out;
 wire sw_212_latch_out;
 wire \sw_212_module_data_in[0] ;
 wire \sw_212_module_data_in[1] ;
 wire \sw_212_module_data_in[2] ;
 wire \sw_212_module_data_in[3] ;
 wire \sw_212_module_data_in[4] ;
 wire \sw_212_module_data_in[5] ;
 wire \sw_212_module_data_in[6] ;
 wire \sw_212_module_data_in[7] ;
 wire \sw_212_module_data_out[0] ;
 wire \sw_212_module_data_out[1] ;
 wire \sw_212_module_data_out[2] ;
 wire \sw_212_module_data_out[3] ;
 wire \sw_212_module_data_out[4] ;
 wire \sw_212_module_data_out[5] ;
 wire \sw_212_module_data_out[6] ;
 wire \sw_212_module_data_out[7] ;
 wire sw_212_scan_out;
 wire sw_213_clk_out;
 wire sw_213_data_out;
 wire sw_213_latch_out;
 wire \sw_213_module_data_in[0] ;
 wire \sw_213_module_data_in[1] ;
 wire \sw_213_module_data_in[2] ;
 wire \sw_213_module_data_in[3] ;
 wire \sw_213_module_data_in[4] ;
 wire \sw_213_module_data_in[5] ;
 wire \sw_213_module_data_in[6] ;
 wire \sw_213_module_data_in[7] ;
 wire \sw_213_module_data_out[0] ;
 wire \sw_213_module_data_out[1] ;
 wire \sw_213_module_data_out[2] ;
 wire \sw_213_module_data_out[3] ;
 wire \sw_213_module_data_out[4] ;
 wire \sw_213_module_data_out[5] ;
 wire \sw_213_module_data_out[6] ;
 wire \sw_213_module_data_out[7] ;
 wire sw_213_scan_out;
 wire sw_214_clk_out;
 wire sw_214_data_out;
 wire sw_214_latch_out;
 wire \sw_214_module_data_in[0] ;
 wire \sw_214_module_data_in[1] ;
 wire \sw_214_module_data_in[2] ;
 wire \sw_214_module_data_in[3] ;
 wire \sw_214_module_data_in[4] ;
 wire \sw_214_module_data_in[5] ;
 wire \sw_214_module_data_in[6] ;
 wire \sw_214_module_data_in[7] ;
 wire \sw_214_module_data_out[0] ;
 wire \sw_214_module_data_out[1] ;
 wire \sw_214_module_data_out[2] ;
 wire \sw_214_module_data_out[3] ;
 wire \sw_214_module_data_out[4] ;
 wire \sw_214_module_data_out[5] ;
 wire \sw_214_module_data_out[6] ;
 wire \sw_214_module_data_out[7] ;
 wire sw_214_scan_out;
 wire sw_215_clk_out;
 wire sw_215_data_out;
 wire sw_215_latch_out;
 wire \sw_215_module_data_in[0] ;
 wire \sw_215_module_data_in[1] ;
 wire \sw_215_module_data_in[2] ;
 wire \sw_215_module_data_in[3] ;
 wire \sw_215_module_data_in[4] ;
 wire \sw_215_module_data_in[5] ;
 wire \sw_215_module_data_in[6] ;
 wire \sw_215_module_data_in[7] ;
 wire \sw_215_module_data_out[0] ;
 wire \sw_215_module_data_out[1] ;
 wire \sw_215_module_data_out[2] ;
 wire \sw_215_module_data_out[3] ;
 wire \sw_215_module_data_out[4] ;
 wire \sw_215_module_data_out[5] ;
 wire \sw_215_module_data_out[6] ;
 wire \sw_215_module_data_out[7] ;
 wire sw_215_scan_out;
 wire sw_216_clk_out;
 wire sw_216_data_out;
 wire sw_216_latch_out;
 wire \sw_216_module_data_in[0] ;
 wire \sw_216_module_data_in[1] ;
 wire \sw_216_module_data_in[2] ;
 wire \sw_216_module_data_in[3] ;
 wire \sw_216_module_data_in[4] ;
 wire \sw_216_module_data_in[5] ;
 wire \sw_216_module_data_in[6] ;
 wire \sw_216_module_data_in[7] ;
 wire \sw_216_module_data_out[0] ;
 wire \sw_216_module_data_out[1] ;
 wire \sw_216_module_data_out[2] ;
 wire \sw_216_module_data_out[3] ;
 wire \sw_216_module_data_out[4] ;
 wire \sw_216_module_data_out[5] ;
 wire \sw_216_module_data_out[6] ;
 wire \sw_216_module_data_out[7] ;
 wire sw_216_scan_out;
 wire sw_217_clk_out;
 wire sw_217_data_out;
 wire sw_217_latch_out;
 wire \sw_217_module_data_in[0] ;
 wire \sw_217_module_data_in[1] ;
 wire \sw_217_module_data_in[2] ;
 wire \sw_217_module_data_in[3] ;
 wire \sw_217_module_data_in[4] ;
 wire \sw_217_module_data_in[5] ;
 wire \sw_217_module_data_in[6] ;
 wire \sw_217_module_data_in[7] ;
 wire \sw_217_module_data_out[0] ;
 wire \sw_217_module_data_out[1] ;
 wire \sw_217_module_data_out[2] ;
 wire \sw_217_module_data_out[3] ;
 wire \sw_217_module_data_out[4] ;
 wire \sw_217_module_data_out[5] ;
 wire \sw_217_module_data_out[6] ;
 wire \sw_217_module_data_out[7] ;
 wire sw_217_scan_out;
 wire sw_218_clk_out;
 wire sw_218_data_out;
 wire sw_218_latch_out;
 wire \sw_218_module_data_in[0] ;
 wire \sw_218_module_data_in[1] ;
 wire \sw_218_module_data_in[2] ;
 wire \sw_218_module_data_in[3] ;
 wire \sw_218_module_data_in[4] ;
 wire \sw_218_module_data_in[5] ;
 wire \sw_218_module_data_in[6] ;
 wire \sw_218_module_data_in[7] ;
 wire \sw_218_module_data_out[0] ;
 wire \sw_218_module_data_out[1] ;
 wire \sw_218_module_data_out[2] ;
 wire \sw_218_module_data_out[3] ;
 wire \sw_218_module_data_out[4] ;
 wire \sw_218_module_data_out[5] ;
 wire \sw_218_module_data_out[6] ;
 wire \sw_218_module_data_out[7] ;
 wire sw_218_scan_out;
 wire sw_219_clk_out;
 wire sw_219_data_out;
 wire sw_219_latch_out;
 wire \sw_219_module_data_in[0] ;
 wire \sw_219_module_data_in[1] ;
 wire \sw_219_module_data_in[2] ;
 wire \sw_219_module_data_in[3] ;
 wire \sw_219_module_data_in[4] ;
 wire \sw_219_module_data_in[5] ;
 wire \sw_219_module_data_in[6] ;
 wire \sw_219_module_data_in[7] ;
 wire \sw_219_module_data_out[0] ;
 wire \sw_219_module_data_out[1] ;
 wire \sw_219_module_data_out[2] ;
 wire \sw_219_module_data_out[3] ;
 wire \sw_219_module_data_out[4] ;
 wire \sw_219_module_data_out[5] ;
 wire \sw_219_module_data_out[6] ;
 wire \sw_219_module_data_out[7] ;
 wire sw_219_scan_out;
 wire sw_220_clk_out;
 wire sw_220_data_out;
 wire sw_220_latch_out;
 wire \sw_220_module_data_in[0] ;
 wire \sw_220_module_data_in[1] ;
 wire \sw_220_module_data_in[2] ;
 wire \sw_220_module_data_in[3] ;
 wire \sw_220_module_data_in[4] ;
 wire \sw_220_module_data_in[5] ;
 wire \sw_220_module_data_in[6] ;
 wire \sw_220_module_data_in[7] ;
 wire \sw_220_module_data_out[0] ;
 wire \sw_220_module_data_out[1] ;
 wire \sw_220_module_data_out[2] ;
 wire \sw_220_module_data_out[3] ;
 wire \sw_220_module_data_out[4] ;
 wire \sw_220_module_data_out[5] ;
 wire \sw_220_module_data_out[6] ;
 wire \sw_220_module_data_out[7] ;
 wire sw_220_scan_out;
 wire sw_221_clk_out;
 wire sw_221_data_out;
 wire sw_221_latch_out;
 wire \sw_221_module_data_in[0] ;
 wire \sw_221_module_data_in[1] ;
 wire \sw_221_module_data_in[2] ;
 wire \sw_221_module_data_in[3] ;
 wire \sw_221_module_data_in[4] ;
 wire \sw_221_module_data_in[5] ;
 wire \sw_221_module_data_in[6] ;
 wire \sw_221_module_data_in[7] ;
 wire \sw_221_module_data_out[0] ;
 wire \sw_221_module_data_out[1] ;
 wire \sw_221_module_data_out[2] ;
 wire \sw_221_module_data_out[3] ;
 wire \sw_221_module_data_out[4] ;
 wire \sw_221_module_data_out[5] ;
 wire \sw_221_module_data_out[6] ;
 wire \sw_221_module_data_out[7] ;
 wire sw_221_scan_out;
 wire sw_222_clk_out;
 wire sw_222_data_out;
 wire sw_222_latch_out;
 wire \sw_222_module_data_in[0] ;
 wire \sw_222_module_data_in[1] ;
 wire \sw_222_module_data_in[2] ;
 wire \sw_222_module_data_in[3] ;
 wire \sw_222_module_data_in[4] ;
 wire \sw_222_module_data_in[5] ;
 wire \sw_222_module_data_in[6] ;
 wire \sw_222_module_data_in[7] ;
 wire \sw_222_module_data_out[0] ;
 wire \sw_222_module_data_out[1] ;
 wire \sw_222_module_data_out[2] ;
 wire \sw_222_module_data_out[3] ;
 wire \sw_222_module_data_out[4] ;
 wire \sw_222_module_data_out[5] ;
 wire \sw_222_module_data_out[6] ;
 wire \sw_222_module_data_out[7] ;
 wire sw_222_scan_out;
 wire sw_223_clk_out;
 wire sw_223_data_out;
 wire sw_223_latch_out;
 wire \sw_223_module_data_in[0] ;
 wire \sw_223_module_data_in[1] ;
 wire \sw_223_module_data_in[2] ;
 wire \sw_223_module_data_in[3] ;
 wire \sw_223_module_data_in[4] ;
 wire \sw_223_module_data_in[5] ;
 wire \sw_223_module_data_in[6] ;
 wire \sw_223_module_data_in[7] ;
 wire \sw_223_module_data_out[0] ;
 wire \sw_223_module_data_out[1] ;
 wire \sw_223_module_data_out[2] ;
 wire \sw_223_module_data_out[3] ;
 wire \sw_223_module_data_out[4] ;
 wire \sw_223_module_data_out[5] ;
 wire \sw_223_module_data_out[6] ;
 wire \sw_223_module_data_out[7] ;
 wire sw_223_scan_out;
 wire sw_224_clk_out;
 wire sw_224_data_out;
 wire sw_224_latch_out;
 wire \sw_224_module_data_in[0] ;
 wire \sw_224_module_data_in[1] ;
 wire \sw_224_module_data_in[2] ;
 wire \sw_224_module_data_in[3] ;
 wire \sw_224_module_data_in[4] ;
 wire \sw_224_module_data_in[5] ;
 wire \sw_224_module_data_in[6] ;
 wire \sw_224_module_data_in[7] ;
 wire \sw_224_module_data_out[0] ;
 wire \sw_224_module_data_out[1] ;
 wire \sw_224_module_data_out[2] ;
 wire \sw_224_module_data_out[3] ;
 wire \sw_224_module_data_out[4] ;
 wire \sw_224_module_data_out[5] ;
 wire \sw_224_module_data_out[6] ;
 wire \sw_224_module_data_out[7] ;
 wire sw_224_scan_out;
 wire sw_225_clk_out;
 wire sw_225_data_out;
 wire sw_225_latch_out;
 wire \sw_225_module_data_in[0] ;
 wire \sw_225_module_data_in[1] ;
 wire \sw_225_module_data_in[2] ;
 wire \sw_225_module_data_in[3] ;
 wire \sw_225_module_data_in[4] ;
 wire \sw_225_module_data_in[5] ;
 wire \sw_225_module_data_in[6] ;
 wire \sw_225_module_data_in[7] ;
 wire \sw_225_module_data_out[0] ;
 wire \sw_225_module_data_out[1] ;
 wire \sw_225_module_data_out[2] ;
 wire \sw_225_module_data_out[3] ;
 wire \sw_225_module_data_out[4] ;
 wire \sw_225_module_data_out[5] ;
 wire \sw_225_module_data_out[6] ;
 wire \sw_225_module_data_out[7] ;
 wire sw_225_scan_out;
 wire sw_226_clk_out;
 wire sw_226_data_out;
 wire sw_226_latch_out;
 wire \sw_226_module_data_in[0] ;
 wire \sw_226_module_data_in[1] ;
 wire \sw_226_module_data_in[2] ;
 wire \sw_226_module_data_in[3] ;
 wire \sw_226_module_data_in[4] ;
 wire \sw_226_module_data_in[5] ;
 wire \sw_226_module_data_in[6] ;
 wire \sw_226_module_data_in[7] ;
 wire \sw_226_module_data_out[0] ;
 wire \sw_226_module_data_out[1] ;
 wire \sw_226_module_data_out[2] ;
 wire \sw_226_module_data_out[3] ;
 wire \sw_226_module_data_out[4] ;
 wire \sw_226_module_data_out[5] ;
 wire \sw_226_module_data_out[6] ;
 wire \sw_226_module_data_out[7] ;
 wire sw_226_scan_out;
 wire sw_227_clk_out;
 wire sw_227_data_out;
 wire sw_227_latch_out;
 wire \sw_227_module_data_in[0] ;
 wire \sw_227_module_data_in[1] ;
 wire \sw_227_module_data_in[2] ;
 wire \sw_227_module_data_in[3] ;
 wire \sw_227_module_data_in[4] ;
 wire \sw_227_module_data_in[5] ;
 wire \sw_227_module_data_in[6] ;
 wire \sw_227_module_data_in[7] ;
 wire \sw_227_module_data_out[0] ;
 wire \sw_227_module_data_out[1] ;
 wire \sw_227_module_data_out[2] ;
 wire \sw_227_module_data_out[3] ;
 wire \sw_227_module_data_out[4] ;
 wire \sw_227_module_data_out[5] ;
 wire \sw_227_module_data_out[6] ;
 wire \sw_227_module_data_out[7] ;
 wire sw_227_scan_out;
 wire sw_228_clk_out;
 wire sw_228_data_out;
 wire sw_228_latch_out;
 wire \sw_228_module_data_in[0] ;
 wire \sw_228_module_data_in[1] ;
 wire \sw_228_module_data_in[2] ;
 wire \sw_228_module_data_in[3] ;
 wire \sw_228_module_data_in[4] ;
 wire \sw_228_module_data_in[5] ;
 wire \sw_228_module_data_in[6] ;
 wire \sw_228_module_data_in[7] ;
 wire \sw_228_module_data_out[0] ;
 wire \sw_228_module_data_out[1] ;
 wire \sw_228_module_data_out[2] ;
 wire \sw_228_module_data_out[3] ;
 wire \sw_228_module_data_out[4] ;
 wire \sw_228_module_data_out[5] ;
 wire \sw_228_module_data_out[6] ;
 wire \sw_228_module_data_out[7] ;
 wire sw_228_scan_out;
 wire sw_229_clk_out;
 wire sw_229_data_out;
 wire sw_229_latch_out;
 wire \sw_229_module_data_in[0] ;
 wire \sw_229_module_data_in[1] ;
 wire \sw_229_module_data_in[2] ;
 wire \sw_229_module_data_in[3] ;
 wire \sw_229_module_data_in[4] ;
 wire \sw_229_module_data_in[5] ;
 wire \sw_229_module_data_in[6] ;
 wire \sw_229_module_data_in[7] ;
 wire \sw_229_module_data_out[0] ;
 wire \sw_229_module_data_out[1] ;
 wire \sw_229_module_data_out[2] ;
 wire \sw_229_module_data_out[3] ;
 wire \sw_229_module_data_out[4] ;
 wire \sw_229_module_data_out[5] ;
 wire \sw_229_module_data_out[6] ;
 wire \sw_229_module_data_out[7] ;
 wire sw_229_scan_out;
 wire sw_230_clk_out;
 wire sw_230_data_out;
 wire sw_230_latch_out;
 wire \sw_230_module_data_in[0] ;
 wire \sw_230_module_data_in[1] ;
 wire \sw_230_module_data_in[2] ;
 wire \sw_230_module_data_in[3] ;
 wire \sw_230_module_data_in[4] ;
 wire \sw_230_module_data_in[5] ;
 wire \sw_230_module_data_in[6] ;
 wire \sw_230_module_data_in[7] ;
 wire \sw_230_module_data_out[0] ;
 wire \sw_230_module_data_out[1] ;
 wire \sw_230_module_data_out[2] ;
 wire \sw_230_module_data_out[3] ;
 wire \sw_230_module_data_out[4] ;
 wire \sw_230_module_data_out[5] ;
 wire \sw_230_module_data_out[6] ;
 wire \sw_230_module_data_out[7] ;
 wire sw_230_scan_out;
 wire sw_231_clk_out;
 wire sw_231_data_out;
 wire sw_231_latch_out;
 wire \sw_231_module_data_in[0] ;
 wire \sw_231_module_data_in[1] ;
 wire \sw_231_module_data_in[2] ;
 wire \sw_231_module_data_in[3] ;
 wire \sw_231_module_data_in[4] ;
 wire \sw_231_module_data_in[5] ;
 wire \sw_231_module_data_in[6] ;
 wire \sw_231_module_data_in[7] ;
 wire \sw_231_module_data_out[0] ;
 wire \sw_231_module_data_out[1] ;
 wire \sw_231_module_data_out[2] ;
 wire \sw_231_module_data_out[3] ;
 wire \sw_231_module_data_out[4] ;
 wire \sw_231_module_data_out[5] ;
 wire \sw_231_module_data_out[6] ;
 wire \sw_231_module_data_out[7] ;
 wire sw_231_scan_out;
 wire sw_232_clk_out;
 wire sw_232_data_out;
 wire sw_232_latch_out;
 wire \sw_232_module_data_in[0] ;
 wire \sw_232_module_data_in[1] ;
 wire \sw_232_module_data_in[2] ;
 wire \sw_232_module_data_in[3] ;
 wire \sw_232_module_data_in[4] ;
 wire \sw_232_module_data_in[5] ;
 wire \sw_232_module_data_in[6] ;
 wire \sw_232_module_data_in[7] ;
 wire \sw_232_module_data_out[0] ;
 wire \sw_232_module_data_out[1] ;
 wire \sw_232_module_data_out[2] ;
 wire \sw_232_module_data_out[3] ;
 wire \sw_232_module_data_out[4] ;
 wire \sw_232_module_data_out[5] ;
 wire \sw_232_module_data_out[6] ;
 wire \sw_232_module_data_out[7] ;
 wire sw_232_scan_out;
 wire sw_233_clk_out;
 wire sw_233_data_out;
 wire sw_233_latch_out;
 wire \sw_233_module_data_in[0] ;
 wire \sw_233_module_data_in[1] ;
 wire \sw_233_module_data_in[2] ;
 wire \sw_233_module_data_in[3] ;
 wire \sw_233_module_data_in[4] ;
 wire \sw_233_module_data_in[5] ;
 wire \sw_233_module_data_in[6] ;
 wire \sw_233_module_data_in[7] ;
 wire \sw_233_module_data_out[0] ;
 wire \sw_233_module_data_out[1] ;
 wire \sw_233_module_data_out[2] ;
 wire \sw_233_module_data_out[3] ;
 wire \sw_233_module_data_out[4] ;
 wire \sw_233_module_data_out[5] ;
 wire \sw_233_module_data_out[6] ;
 wire \sw_233_module_data_out[7] ;
 wire sw_233_scan_out;
 wire sw_234_clk_out;
 wire sw_234_data_out;
 wire sw_234_latch_out;
 wire \sw_234_module_data_in[0] ;
 wire \sw_234_module_data_in[1] ;
 wire \sw_234_module_data_in[2] ;
 wire \sw_234_module_data_in[3] ;
 wire \sw_234_module_data_in[4] ;
 wire \sw_234_module_data_in[5] ;
 wire \sw_234_module_data_in[6] ;
 wire \sw_234_module_data_in[7] ;
 wire \sw_234_module_data_out[0] ;
 wire \sw_234_module_data_out[1] ;
 wire \sw_234_module_data_out[2] ;
 wire \sw_234_module_data_out[3] ;
 wire \sw_234_module_data_out[4] ;
 wire \sw_234_module_data_out[5] ;
 wire \sw_234_module_data_out[6] ;
 wire \sw_234_module_data_out[7] ;
 wire sw_234_scan_out;
 wire sw_235_clk_out;
 wire sw_235_data_out;
 wire sw_235_latch_out;
 wire \sw_235_module_data_in[0] ;
 wire \sw_235_module_data_in[1] ;
 wire \sw_235_module_data_in[2] ;
 wire \sw_235_module_data_in[3] ;
 wire \sw_235_module_data_in[4] ;
 wire \sw_235_module_data_in[5] ;
 wire \sw_235_module_data_in[6] ;
 wire \sw_235_module_data_in[7] ;
 wire \sw_235_module_data_out[0] ;
 wire \sw_235_module_data_out[1] ;
 wire \sw_235_module_data_out[2] ;
 wire \sw_235_module_data_out[3] ;
 wire \sw_235_module_data_out[4] ;
 wire \sw_235_module_data_out[5] ;
 wire \sw_235_module_data_out[6] ;
 wire \sw_235_module_data_out[7] ;
 wire sw_235_scan_out;
 wire sw_236_clk_out;
 wire sw_236_data_out;
 wire sw_236_latch_out;
 wire \sw_236_module_data_in[0] ;
 wire \sw_236_module_data_in[1] ;
 wire \sw_236_module_data_in[2] ;
 wire \sw_236_module_data_in[3] ;
 wire \sw_236_module_data_in[4] ;
 wire \sw_236_module_data_in[5] ;
 wire \sw_236_module_data_in[6] ;
 wire \sw_236_module_data_in[7] ;
 wire \sw_236_module_data_out[0] ;
 wire \sw_236_module_data_out[1] ;
 wire \sw_236_module_data_out[2] ;
 wire \sw_236_module_data_out[3] ;
 wire \sw_236_module_data_out[4] ;
 wire \sw_236_module_data_out[5] ;
 wire \sw_236_module_data_out[6] ;
 wire \sw_236_module_data_out[7] ;
 wire sw_236_scan_out;
 wire sw_237_clk_out;
 wire sw_237_data_out;
 wire sw_237_latch_out;
 wire \sw_237_module_data_in[0] ;
 wire \sw_237_module_data_in[1] ;
 wire \sw_237_module_data_in[2] ;
 wire \sw_237_module_data_in[3] ;
 wire \sw_237_module_data_in[4] ;
 wire \sw_237_module_data_in[5] ;
 wire \sw_237_module_data_in[6] ;
 wire \sw_237_module_data_in[7] ;
 wire \sw_237_module_data_out[0] ;
 wire \sw_237_module_data_out[1] ;
 wire \sw_237_module_data_out[2] ;
 wire \sw_237_module_data_out[3] ;
 wire \sw_237_module_data_out[4] ;
 wire \sw_237_module_data_out[5] ;
 wire \sw_237_module_data_out[6] ;
 wire \sw_237_module_data_out[7] ;
 wire sw_237_scan_out;
 wire sw_238_clk_out;
 wire sw_238_data_out;
 wire sw_238_latch_out;
 wire \sw_238_module_data_in[0] ;
 wire \sw_238_module_data_in[1] ;
 wire \sw_238_module_data_in[2] ;
 wire \sw_238_module_data_in[3] ;
 wire \sw_238_module_data_in[4] ;
 wire \sw_238_module_data_in[5] ;
 wire \sw_238_module_data_in[6] ;
 wire \sw_238_module_data_in[7] ;
 wire \sw_238_module_data_out[0] ;
 wire \sw_238_module_data_out[1] ;
 wire \sw_238_module_data_out[2] ;
 wire \sw_238_module_data_out[3] ;
 wire \sw_238_module_data_out[4] ;
 wire \sw_238_module_data_out[5] ;
 wire \sw_238_module_data_out[6] ;
 wire \sw_238_module_data_out[7] ;
 wire sw_238_scan_out;
 wire sw_239_clk_out;
 wire sw_239_data_out;
 wire sw_239_latch_out;
 wire \sw_239_module_data_in[0] ;
 wire \sw_239_module_data_in[1] ;
 wire \sw_239_module_data_in[2] ;
 wire \sw_239_module_data_in[3] ;
 wire \sw_239_module_data_in[4] ;
 wire \sw_239_module_data_in[5] ;
 wire \sw_239_module_data_in[6] ;
 wire \sw_239_module_data_in[7] ;
 wire \sw_239_module_data_out[0] ;
 wire \sw_239_module_data_out[1] ;
 wire \sw_239_module_data_out[2] ;
 wire \sw_239_module_data_out[3] ;
 wire \sw_239_module_data_out[4] ;
 wire \sw_239_module_data_out[5] ;
 wire \sw_239_module_data_out[6] ;
 wire \sw_239_module_data_out[7] ;
 wire sw_239_scan_out;
 wire sw_240_clk_out;
 wire sw_240_data_out;
 wire sw_240_latch_out;
 wire \sw_240_module_data_in[0] ;
 wire \sw_240_module_data_in[1] ;
 wire \sw_240_module_data_in[2] ;
 wire \sw_240_module_data_in[3] ;
 wire \sw_240_module_data_in[4] ;
 wire \sw_240_module_data_in[5] ;
 wire \sw_240_module_data_in[6] ;
 wire \sw_240_module_data_in[7] ;
 wire \sw_240_module_data_out[0] ;
 wire \sw_240_module_data_out[1] ;
 wire \sw_240_module_data_out[2] ;
 wire \sw_240_module_data_out[3] ;
 wire \sw_240_module_data_out[4] ;
 wire \sw_240_module_data_out[5] ;
 wire \sw_240_module_data_out[6] ;
 wire \sw_240_module_data_out[7] ;
 wire sw_240_scan_out;
 wire sw_241_clk_out;
 wire sw_241_data_out;
 wire sw_241_latch_out;
 wire \sw_241_module_data_in[0] ;
 wire \sw_241_module_data_in[1] ;
 wire \sw_241_module_data_in[2] ;
 wire \sw_241_module_data_in[3] ;
 wire \sw_241_module_data_in[4] ;
 wire \sw_241_module_data_in[5] ;
 wire \sw_241_module_data_in[6] ;
 wire \sw_241_module_data_in[7] ;
 wire \sw_241_module_data_out[0] ;
 wire \sw_241_module_data_out[1] ;
 wire \sw_241_module_data_out[2] ;
 wire \sw_241_module_data_out[3] ;
 wire \sw_241_module_data_out[4] ;
 wire \sw_241_module_data_out[5] ;
 wire \sw_241_module_data_out[6] ;
 wire \sw_241_module_data_out[7] ;
 wire sw_241_scan_out;
 wire sw_242_clk_out;
 wire sw_242_data_out;
 wire sw_242_latch_out;
 wire \sw_242_module_data_in[0] ;
 wire \sw_242_module_data_in[1] ;
 wire \sw_242_module_data_in[2] ;
 wire \sw_242_module_data_in[3] ;
 wire \sw_242_module_data_in[4] ;
 wire \sw_242_module_data_in[5] ;
 wire \sw_242_module_data_in[6] ;
 wire \sw_242_module_data_in[7] ;
 wire \sw_242_module_data_out[0] ;
 wire \sw_242_module_data_out[1] ;
 wire \sw_242_module_data_out[2] ;
 wire \sw_242_module_data_out[3] ;
 wire \sw_242_module_data_out[4] ;
 wire \sw_242_module_data_out[5] ;
 wire \sw_242_module_data_out[6] ;
 wire \sw_242_module_data_out[7] ;
 wire sw_242_scan_out;
 wire sw_243_clk_out;
 wire sw_243_data_out;
 wire sw_243_latch_out;
 wire \sw_243_module_data_in[0] ;
 wire \sw_243_module_data_in[1] ;
 wire \sw_243_module_data_in[2] ;
 wire \sw_243_module_data_in[3] ;
 wire \sw_243_module_data_in[4] ;
 wire \sw_243_module_data_in[5] ;
 wire \sw_243_module_data_in[6] ;
 wire \sw_243_module_data_in[7] ;
 wire \sw_243_module_data_out[0] ;
 wire \sw_243_module_data_out[1] ;
 wire \sw_243_module_data_out[2] ;
 wire \sw_243_module_data_out[3] ;
 wire \sw_243_module_data_out[4] ;
 wire \sw_243_module_data_out[5] ;
 wire \sw_243_module_data_out[6] ;
 wire \sw_243_module_data_out[7] ;
 wire sw_243_scan_out;
 wire sw_244_clk_out;
 wire sw_244_data_out;
 wire sw_244_latch_out;
 wire \sw_244_module_data_in[0] ;
 wire \sw_244_module_data_in[1] ;
 wire \sw_244_module_data_in[2] ;
 wire \sw_244_module_data_in[3] ;
 wire \sw_244_module_data_in[4] ;
 wire \sw_244_module_data_in[5] ;
 wire \sw_244_module_data_in[6] ;
 wire \sw_244_module_data_in[7] ;
 wire \sw_244_module_data_out[0] ;
 wire \sw_244_module_data_out[1] ;
 wire \sw_244_module_data_out[2] ;
 wire \sw_244_module_data_out[3] ;
 wire \sw_244_module_data_out[4] ;
 wire \sw_244_module_data_out[5] ;
 wire \sw_244_module_data_out[6] ;
 wire \sw_244_module_data_out[7] ;
 wire sw_244_scan_out;
 wire sw_245_clk_out;
 wire sw_245_data_out;
 wire sw_245_latch_out;
 wire \sw_245_module_data_in[0] ;
 wire \sw_245_module_data_in[1] ;
 wire \sw_245_module_data_in[2] ;
 wire \sw_245_module_data_in[3] ;
 wire \sw_245_module_data_in[4] ;
 wire \sw_245_module_data_in[5] ;
 wire \sw_245_module_data_in[6] ;
 wire \sw_245_module_data_in[7] ;
 wire \sw_245_module_data_out[0] ;
 wire \sw_245_module_data_out[1] ;
 wire \sw_245_module_data_out[2] ;
 wire \sw_245_module_data_out[3] ;
 wire \sw_245_module_data_out[4] ;
 wire \sw_245_module_data_out[5] ;
 wire \sw_245_module_data_out[6] ;
 wire \sw_245_module_data_out[7] ;
 wire sw_245_scan_out;
 wire sw_246_clk_out;
 wire sw_246_data_out;
 wire sw_246_latch_out;
 wire \sw_246_module_data_in[0] ;
 wire \sw_246_module_data_in[1] ;
 wire \sw_246_module_data_in[2] ;
 wire \sw_246_module_data_in[3] ;
 wire \sw_246_module_data_in[4] ;
 wire \sw_246_module_data_in[5] ;
 wire \sw_246_module_data_in[6] ;
 wire \sw_246_module_data_in[7] ;
 wire \sw_246_module_data_out[0] ;
 wire \sw_246_module_data_out[1] ;
 wire \sw_246_module_data_out[2] ;
 wire \sw_246_module_data_out[3] ;
 wire \sw_246_module_data_out[4] ;
 wire \sw_246_module_data_out[5] ;
 wire \sw_246_module_data_out[6] ;
 wire \sw_246_module_data_out[7] ;
 wire sw_246_scan_out;
 wire sw_247_clk_out;
 wire sw_247_data_out;
 wire sw_247_latch_out;
 wire \sw_247_module_data_in[0] ;
 wire \sw_247_module_data_in[1] ;
 wire \sw_247_module_data_in[2] ;
 wire \sw_247_module_data_in[3] ;
 wire \sw_247_module_data_in[4] ;
 wire \sw_247_module_data_in[5] ;
 wire \sw_247_module_data_in[6] ;
 wire \sw_247_module_data_in[7] ;
 wire \sw_247_module_data_out[0] ;
 wire \sw_247_module_data_out[1] ;
 wire \sw_247_module_data_out[2] ;
 wire \sw_247_module_data_out[3] ;
 wire \sw_247_module_data_out[4] ;
 wire \sw_247_module_data_out[5] ;
 wire \sw_247_module_data_out[6] ;
 wire \sw_247_module_data_out[7] ;
 wire sw_247_scan_out;
 wire sw_248_clk_out;
 wire sw_248_data_out;
 wire sw_248_latch_out;
 wire \sw_248_module_data_in[0] ;
 wire \sw_248_module_data_in[1] ;
 wire \sw_248_module_data_in[2] ;
 wire \sw_248_module_data_in[3] ;
 wire \sw_248_module_data_in[4] ;
 wire \sw_248_module_data_in[5] ;
 wire \sw_248_module_data_in[6] ;
 wire \sw_248_module_data_in[7] ;
 wire \sw_248_module_data_out[0] ;
 wire \sw_248_module_data_out[1] ;
 wire \sw_248_module_data_out[2] ;
 wire \sw_248_module_data_out[3] ;
 wire \sw_248_module_data_out[4] ;
 wire \sw_248_module_data_out[5] ;
 wire \sw_248_module_data_out[6] ;
 wire \sw_248_module_data_out[7] ;
 wire sw_248_scan_out;
 wire sw_249_clk_out;
 wire sw_249_data_out;
 wire sw_249_latch_out;
 wire \sw_249_module_data_in[0] ;
 wire \sw_249_module_data_in[1] ;
 wire \sw_249_module_data_in[2] ;
 wire \sw_249_module_data_in[3] ;
 wire \sw_249_module_data_in[4] ;
 wire \sw_249_module_data_in[5] ;
 wire \sw_249_module_data_in[6] ;
 wire \sw_249_module_data_in[7] ;
 wire \sw_249_module_data_out[0] ;
 wire \sw_249_module_data_out[1] ;
 wire \sw_249_module_data_out[2] ;
 wire \sw_249_module_data_out[3] ;
 wire \sw_249_module_data_out[4] ;
 wire \sw_249_module_data_out[5] ;
 wire \sw_249_module_data_out[6] ;
 wire \sw_249_module_data_out[7] ;
 wire sw_249_scan_out;
 wire sw_250_clk_out;
 wire sw_250_data_out;
 wire sw_250_latch_out;
 wire \sw_250_module_data_in[0] ;
 wire \sw_250_module_data_in[1] ;
 wire \sw_250_module_data_in[2] ;
 wire \sw_250_module_data_in[3] ;
 wire \sw_250_module_data_in[4] ;
 wire \sw_250_module_data_in[5] ;
 wire \sw_250_module_data_in[6] ;
 wire \sw_250_module_data_in[7] ;
 wire \sw_250_module_data_out[0] ;
 wire \sw_250_module_data_out[1] ;
 wire \sw_250_module_data_out[2] ;
 wire \sw_250_module_data_out[3] ;
 wire \sw_250_module_data_out[4] ;
 wire \sw_250_module_data_out[5] ;
 wire \sw_250_module_data_out[6] ;
 wire \sw_250_module_data_out[7] ;
 wire sw_250_scan_out;
 wire sw_251_clk_out;
 wire sw_251_data_out;
 wire sw_251_latch_out;
 wire \sw_251_module_data_in[0] ;
 wire \sw_251_module_data_in[1] ;
 wire \sw_251_module_data_in[2] ;
 wire \sw_251_module_data_in[3] ;
 wire \sw_251_module_data_in[4] ;
 wire \sw_251_module_data_in[5] ;
 wire \sw_251_module_data_in[6] ;
 wire \sw_251_module_data_in[7] ;
 wire \sw_251_module_data_out[0] ;
 wire \sw_251_module_data_out[1] ;
 wire \sw_251_module_data_out[2] ;
 wire \sw_251_module_data_out[3] ;
 wire \sw_251_module_data_out[4] ;
 wire \sw_251_module_data_out[5] ;
 wire \sw_251_module_data_out[6] ;
 wire \sw_251_module_data_out[7] ;
 wire sw_251_scan_out;
 wire sw_252_clk_out;
 wire sw_252_data_out;
 wire sw_252_latch_out;
 wire \sw_252_module_data_in[0] ;
 wire \sw_252_module_data_in[1] ;
 wire \sw_252_module_data_in[2] ;
 wire \sw_252_module_data_in[3] ;
 wire \sw_252_module_data_in[4] ;
 wire \sw_252_module_data_in[5] ;
 wire \sw_252_module_data_in[6] ;
 wire \sw_252_module_data_in[7] ;
 wire \sw_252_module_data_out[0] ;
 wire \sw_252_module_data_out[1] ;
 wire \sw_252_module_data_out[2] ;
 wire \sw_252_module_data_out[3] ;
 wire \sw_252_module_data_out[4] ;
 wire \sw_252_module_data_out[5] ;
 wire \sw_252_module_data_out[6] ;
 wire \sw_252_module_data_out[7] ;
 wire sw_252_scan_out;
 wire sw_253_clk_out;
 wire sw_253_data_out;
 wire sw_253_latch_out;
 wire \sw_253_module_data_in[0] ;
 wire \sw_253_module_data_in[1] ;
 wire \sw_253_module_data_in[2] ;
 wire \sw_253_module_data_in[3] ;
 wire \sw_253_module_data_in[4] ;
 wire \sw_253_module_data_in[5] ;
 wire \sw_253_module_data_in[6] ;
 wire \sw_253_module_data_in[7] ;
 wire \sw_253_module_data_out[0] ;
 wire \sw_253_module_data_out[1] ;
 wire \sw_253_module_data_out[2] ;
 wire \sw_253_module_data_out[3] ;
 wire \sw_253_module_data_out[4] ;
 wire \sw_253_module_data_out[5] ;
 wire \sw_253_module_data_out[6] ;
 wire \sw_253_module_data_out[7] ;
 wire sw_253_scan_out;
 wire sw_254_clk_out;
 wire sw_254_data_out;
 wire sw_254_latch_out;
 wire \sw_254_module_data_in[0] ;
 wire \sw_254_module_data_in[1] ;
 wire \sw_254_module_data_in[2] ;
 wire \sw_254_module_data_in[3] ;
 wire \sw_254_module_data_in[4] ;
 wire \sw_254_module_data_in[5] ;
 wire \sw_254_module_data_in[6] ;
 wire \sw_254_module_data_in[7] ;
 wire \sw_254_module_data_out[0] ;
 wire \sw_254_module_data_out[1] ;
 wire \sw_254_module_data_out[2] ;
 wire \sw_254_module_data_out[3] ;
 wire \sw_254_module_data_out[4] ;
 wire \sw_254_module_data_out[5] ;
 wire \sw_254_module_data_out[6] ;
 wire \sw_254_module_data_out[7] ;
 wire sw_254_scan_out;
 wire sw_255_clk_out;
 wire sw_255_data_out;
 wire sw_255_latch_out;
 wire \sw_255_module_data_in[0] ;
 wire \sw_255_module_data_in[1] ;
 wire \sw_255_module_data_in[2] ;
 wire \sw_255_module_data_in[3] ;
 wire \sw_255_module_data_in[4] ;
 wire \sw_255_module_data_in[5] ;
 wire \sw_255_module_data_in[6] ;
 wire \sw_255_module_data_in[7] ;
 wire \sw_255_module_data_out[0] ;
 wire \sw_255_module_data_out[1] ;
 wire \sw_255_module_data_out[2] ;
 wire \sw_255_module_data_out[3] ;
 wire \sw_255_module_data_out[4] ;
 wire \sw_255_module_data_out[5] ;
 wire \sw_255_module_data_out[6] ;
 wire \sw_255_module_data_out[7] ;
 wire sw_255_scan_out;
 wire sw_256_clk_out;
 wire sw_256_data_out;
 wire sw_256_latch_out;
 wire \sw_256_module_data_in[0] ;
 wire \sw_256_module_data_in[1] ;
 wire \sw_256_module_data_in[2] ;
 wire \sw_256_module_data_in[3] ;
 wire \sw_256_module_data_in[4] ;
 wire \sw_256_module_data_in[5] ;
 wire \sw_256_module_data_in[6] ;
 wire \sw_256_module_data_in[7] ;
 wire \sw_256_module_data_out[0] ;
 wire \sw_256_module_data_out[1] ;
 wire \sw_256_module_data_out[2] ;
 wire \sw_256_module_data_out[3] ;
 wire \sw_256_module_data_out[4] ;
 wire \sw_256_module_data_out[5] ;
 wire \sw_256_module_data_out[6] ;
 wire \sw_256_module_data_out[7] ;
 wire sw_256_scan_out;
 wire sw_257_clk_out;
 wire sw_257_data_out;
 wire sw_257_latch_out;
 wire \sw_257_module_data_in[0] ;
 wire \sw_257_module_data_in[1] ;
 wire \sw_257_module_data_in[2] ;
 wire \sw_257_module_data_in[3] ;
 wire \sw_257_module_data_in[4] ;
 wire \sw_257_module_data_in[5] ;
 wire \sw_257_module_data_in[6] ;
 wire \sw_257_module_data_in[7] ;
 wire \sw_257_module_data_out[0] ;
 wire \sw_257_module_data_out[1] ;
 wire \sw_257_module_data_out[2] ;
 wire \sw_257_module_data_out[3] ;
 wire \sw_257_module_data_out[4] ;
 wire \sw_257_module_data_out[5] ;
 wire \sw_257_module_data_out[6] ;
 wire \sw_257_module_data_out[7] ;
 wire sw_257_scan_out;
 wire sw_258_clk_out;
 wire sw_258_data_out;
 wire sw_258_latch_out;
 wire \sw_258_module_data_in[0] ;
 wire \sw_258_module_data_in[1] ;
 wire \sw_258_module_data_in[2] ;
 wire \sw_258_module_data_in[3] ;
 wire \sw_258_module_data_in[4] ;
 wire \sw_258_module_data_in[5] ;
 wire \sw_258_module_data_in[6] ;
 wire \sw_258_module_data_in[7] ;
 wire \sw_258_module_data_out[0] ;
 wire \sw_258_module_data_out[1] ;
 wire \sw_258_module_data_out[2] ;
 wire \sw_258_module_data_out[3] ;
 wire \sw_258_module_data_out[4] ;
 wire \sw_258_module_data_out[5] ;
 wire \sw_258_module_data_out[6] ;
 wire \sw_258_module_data_out[7] ;
 wire sw_258_scan_out;
 wire sw_259_clk_out;
 wire sw_259_data_out;
 wire sw_259_latch_out;
 wire \sw_259_module_data_in[0] ;
 wire \sw_259_module_data_in[1] ;
 wire \sw_259_module_data_in[2] ;
 wire \sw_259_module_data_in[3] ;
 wire \sw_259_module_data_in[4] ;
 wire \sw_259_module_data_in[5] ;
 wire \sw_259_module_data_in[6] ;
 wire \sw_259_module_data_in[7] ;
 wire \sw_259_module_data_out[0] ;
 wire \sw_259_module_data_out[1] ;
 wire \sw_259_module_data_out[2] ;
 wire \sw_259_module_data_out[3] ;
 wire \sw_259_module_data_out[4] ;
 wire \sw_259_module_data_out[5] ;
 wire \sw_259_module_data_out[6] ;
 wire \sw_259_module_data_out[7] ;
 wire sw_259_scan_out;
 wire sw_260_clk_out;
 wire sw_260_data_out;
 wire sw_260_latch_out;
 wire \sw_260_module_data_in[0] ;
 wire \sw_260_module_data_in[1] ;
 wire \sw_260_module_data_in[2] ;
 wire \sw_260_module_data_in[3] ;
 wire \sw_260_module_data_in[4] ;
 wire \sw_260_module_data_in[5] ;
 wire \sw_260_module_data_in[6] ;
 wire \sw_260_module_data_in[7] ;
 wire \sw_260_module_data_out[0] ;
 wire \sw_260_module_data_out[1] ;
 wire \sw_260_module_data_out[2] ;
 wire \sw_260_module_data_out[3] ;
 wire \sw_260_module_data_out[4] ;
 wire \sw_260_module_data_out[5] ;
 wire \sw_260_module_data_out[6] ;
 wire \sw_260_module_data_out[7] ;
 wire sw_260_scan_out;
 wire sw_261_clk_out;
 wire sw_261_data_out;
 wire sw_261_latch_out;
 wire \sw_261_module_data_in[0] ;
 wire \sw_261_module_data_in[1] ;
 wire \sw_261_module_data_in[2] ;
 wire \sw_261_module_data_in[3] ;
 wire \sw_261_module_data_in[4] ;
 wire \sw_261_module_data_in[5] ;
 wire \sw_261_module_data_in[6] ;
 wire \sw_261_module_data_in[7] ;
 wire \sw_261_module_data_out[0] ;
 wire \sw_261_module_data_out[1] ;
 wire \sw_261_module_data_out[2] ;
 wire \sw_261_module_data_out[3] ;
 wire \sw_261_module_data_out[4] ;
 wire \sw_261_module_data_out[5] ;
 wire \sw_261_module_data_out[6] ;
 wire \sw_261_module_data_out[7] ;
 wire sw_261_scan_out;
 wire sw_262_clk_out;
 wire sw_262_data_out;
 wire sw_262_latch_out;
 wire \sw_262_module_data_in[0] ;
 wire \sw_262_module_data_in[1] ;
 wire \sw_262_module_data_in[2] ;
 wire \sw_262_module_data_in[3] ;
 wire \sw_262_module_data_in[4] ;
 wire \sw_262_module_data_in[5] ;
 wire \sw_262_module_data_in[6] ;
 wire \sw_262_module_data_in[7] ;
 wire \sw_262_module_data_out[0] ;
 wire \sw_262_module_data_out[1] ;
 wire \sw_262_module_data_out[2] ;
 wire \sw_262_module_data_out[3] ;
 wire \sw_262_module_data_out[4] ;
 wire \sw_262_module_data_out[5] ;
 wire \sw_262_module_data_out[6] ;
 wire \sw_262_module_data_out[7] ;
 wire sw_262_scan_out;
 wire sw_263_clk_out;
 wire sw_263_data_out;
 wire sw_263_latch_out;
 wire \sw_263_module_data_in[0] ;
 wire \sw_263_module_data_in[1] ;
 wire \sw_263_module_data_in[2] ;
 wire \sw_263_module_data_in[3] ;
 wire \sw_263_module_data_in[4] ;
 wire \sw_263_module_data_in[5] ;
 wire \sw_263_module_data_in[6] ;
 wire \sw_263_module_data_in[7] ;
 wire \sw_263_module_data_out[0] ;
 wire \sw_263_module_data_out[1] ;
 wire \sw_263_module_data_out[2] ;
 wire \sw_263_module_data_out[3] ;
 wire \sw_263_module_data_out[4] ;
 wire \sw_263_module_data_out[5] ;
 wire \sw_263_module_data_out[6] ;
 wire \sw_263_module_data_out[7] ;
 wire sw_263_scan_out;
 wire sw_264_clk_out;
 wire sw_264_data_out;
 wire sw_264_latch_out;
 wire \sw_264_module_data_in[0] ;
 wire \sw_264_module_data_in[1] ;
 wire \sw_264_module_data_in[2] ;
 wire \sw_264_module_data_in[3] ;
 wire \sw_264_module_data_in[4] ;
 wire \sw_264_module_data_in[5] ;
 wire \sw_264_module_data_in[6] ;
 wire \sw_264_module_data_in[7] ;
 wire \sw_264_module_data_out[0] ;
 wire \sw_264_module_data_out[1] ;
 wire \sw_264_module_data_out[2] ;
 wire \sw_264_module_data_out[3] ;
 wire \sw_264_module_data_out[4] ;
 wire \sw_264_module_data_out[5] ;
 wire \sw_264_module_data_out[6] ;
 wire \sw_264_module_data_out[7] ;
 wire sw_264_scan_out;
 wire sw_265_clk_out;
 wire sw_265_data_out;
 wire sw_265_latch_out;
 wire \sw_265_module_data_in[0] ;
 wire \sw_265_module_data_in[1] ;
 wire \sw_265_module_data_in[2] ;
 wire \sw_265_module_data_in[3] ;
 wire \sw_265_module_data_in[4] ;
 wire \sw_265_module_data_in[5] ;
 wire \sw_265_module_data_in[6] ;
 wire \sw_265_module_data_in[7] ;
 wire \sw_265_module_data_out[0] ;
 wire \sw_265_module_data_out[1] ;
 wire \sw_265_module_data_out[2] ;
 wire \sw_265_module_data_out[3] ;
 wire \sw_265_module_data_out[4] ;
 wire \sw_265_module_data_out[5] ;
 wire \sw_265_module_data_out[6] ;
 wire \sw_265_module_data_out[7] ;
 wire sw_265_scan_out;
 wire sw_266_clk_out;
 wire sw_266_data_out;
 wire sw_266_latch_out;
 wire \sw_266_module_data_in[0] ;
 wire \sw_266_module_data_in[1] ;
 wire \sw_266_module_data_in[2] ;
 wire \sw_266_module_data_in[3] ;
 wire \sw_266_module_data_in[4] ;
 wire \sw_266_module_data_in[5] ;
 wire \sw_266_module_data_in[6] ;
 wire \sw_266_module_data_in[7] ;
 wire \sw_266_module_data_out[0] ;
 wire \sw_266_module_data_out[1] ;
 wire \sw_266_module_data_out[2] ;
 wire \sw_266_module_data_out[3] ;
 wire \sw_266_module_data_out[4] ;
 wire \sw_266_module_data_out[5] ;
 wire \sw_266_module_data_out[6] ;
 wire \sw_266_module_data_out[7] ;
 wire sw_266_scan_out;
 wire sw_267_clk_out;
 wire sw_267_data_out;
 wire sw_267_latch_out;
 wire \sw_267_module_data_in[0] ;
 wire \sw_267_module_data_in[1] ;
 wire \sw_267_module_data_in[2] ;
 wire \sw_267_module_data_in[3] ;
 wire \sw_267_module_data_in[4] ;
 wire \sw_267_module_data_in[5] ;
 wire \sw_267_module_data_in[6] ;
 wire \sw_267_module_data_in[7] ;
 wire \sw_267_module_data_out[0] ;
 wire \sw_267_module_data_out[1] ;
 wire \sw_267_module_data_out[2] ;
 wire \sw_267_module_data_out[3] ;
 wire \sw_267_module_data_out[4] ;
 wire \sw_267_module_data_out[5] ;
 wire \sw_267_module_data_out[6] ;
 wire \sw_267_module_data_out[7] ;
 wire sw_267_scan_out;
 wire sw_268_clk_out;
 wire sw_268_data_out;
 wire sw_268_latch_out;
 wire \sw_268_module_data_in[0] ;
 wire \sw_268_module_data_in[1] ;
 wire \sw_268_module_data_in[2] ;
 wire \sw_268_module_data_in[3] ;
 wire \sw_268_module_data_in[4] ;
 wire \sw_268_module_data_in[5] ;
 wire \sw_268_module_data_in[6] ;
 wire \sw_268_module_data_in[7] ;
 wire \sw_268_module_data_out[0] ;
 wire \sw_268_module_data_out[1] ;
 wire \sw_268_module_data_out[2] ;
 wire \sw_268_module_data_out[3] ;
 wire \sw_268_module_data_out[4] ;
 wire \sw_268_module_data_out[5] ;
 wire \sw_268_module_data_out[6] ;
 wire \sw_268_module_data_out[7] ;
 wire sw_268_scan_out;
 wire sw_269_clk_out;
 wire sw_269_data_out;
 wire sw_269_latch_out;
 wire \sw_269_module_data_in[0] ;
 wire \sw_269_module_data_in[1] ;
 wire \sw_269_module_data_in[2] ;
 wire \sw_269_module_data_in[3] ;
 wire \sw_269_module_data_in[4] ;
 wire \sw_269_module_data_in[5] ;
 wire \sw_269_module_data_in[6] ;
 wire \sw_269_module_data_in[7] ;
 wire \sw_269_module_data_out[0] ;
 wire \sw_269_module_data_out[1] ;
 wire \sw_269_module_data_out[2] ;
 wire \sw_269_module_data_out[3] ;
 wire \sw_269_module_data_out[4] ;
 wire \sw_269_module_data_out[5] ;
 wire \sw_269_module_data_out[6] ;
 wire \sw_269_module_data_out[7] ;
 wire sw_269_scan_out;
 wire sw_270_clk_out;
 wire sw_270_data_out;
 wire sw_270_latch_out;
 wire \sw_270_module_data_in[0] ;
 wire \sw_270_module_data_in[1] ;
 wire \sw_270_module_data_in[2] ;
 wire \sw_270_module_data_in[3] ;
 wire \sw_270_module_data_in[4] ;
 wire \sw_270_module_data_in[5] ;
 wire \sw_270_module_data_in[6] ;
 wire \sw_270_module_data_in[7] ;
 wire \sw_270_module_data_out[0] ;
 wire \sw_270_module_data_out[1] ;
 wire \sw_270_module_data_out[2] ;
 wire \sw_270_module_data_out[3] ;
 wire \sw_270_module_data_out[4] ;
 wire \sw_270_module_data_out[5] ;
 wire \sw_270_module_data_out[6] ;
 wire \sw_270_module_data_out[7] ;
 wire sw_270_scan_out;
 wire sw_271_clk_out;
 wire sw_271_data_out;
 wire sw_271_latch_out;
 wire \sw_271_module_data_in[0] ;
 wire \sw_271_module_data_in[1] ;
 wire \sw_271_module_data_in[2] ;
 wire \sw_271_module_data_in[3] ;
 wire \sw_271_module_data_in[4] ;
 wire \sw_271_module_data_in[5] ;
 wire \sw_271_module_data_in[6] ;
 wire \sw_271_module_data_in[7] ;
 wire \sw_271_module_data_out[0] ;
 wire \sw_271_module_data_out[1] ;
 wire \sw_271_module_data_out[2] ;
 wire \sw_271_module_data_out[3] ;
 wire \sw_271_module_data_out[4] ;
 wire \sw_271_module_data_out[5] ;
 wire \sw_271_module_data_out[6] ;
 wire \sw_271_module_data_out[7] ;
 wire sw_271_scan_out;
 wire sw_272_clk_out;
 wire sw_272_data_out;
 wire sw_272_latch_out;
 wire \sw_272_module_data_in[0] ;
 wire \sw_272_module_data_in[1] ;
 wire \sw_272_module_data_in[2] ;
 wire \sw_272_module_data_in[3] ;
 wire \sw_272_module_data_in[4] ;
 wire \sw_272_module_data_in[5] ;
 wire \sw_272_module_data_in[6] ;
 wire \sw_272_module_data_in[7] ;
 wire \sw_272_module_data_out[0] ;
 wire \sw_272_module_data_out[1] ;
 wire \sw_272_module_data_out[2] ;
 wire \sw_272_module_data_out[3] ;
 wire \sw_272_module_data_out[4] ;
 wire \sw_272_module_data_out[5] ;
 wire \sw_272_module_data_out[6] ;
 wire \sw_272_module_data_out[7] ;
 wire sw_272_scan_out;
 wire sw_273_clk_out;
 wire sw_273_data_out;
 wire sw_273_latch_out;
 wire \sw_273_module_data_in[0] ;
 wire \sw_273_module_data_in[1] ;
 wire \sw_273_module_data_in[2] ;
 wire \sw_273_module_data_in[3] ;
 wire \sw_273_module_data_in[4] ;
 wire \sw_273_module_data_in[5] ;
 wire \sw_273_module_data_in[6] ;
 wire \sw_273_module_data_in[7] ;
 wire \sw_273_module_data_out[0] ;
 wire \sw_273_module_data_out[1] ;
 wire \sw_273_module_data_out[2] ;
 wire \sw_273_module_data_out[3] ;
 wire \sw_273_module_data_out[4] ;
 wire \sw_273_module_data_out[5] ;
 wire \sw_273_module_data_out[6] ;
 wire \sw_273_module_data_out[7] ;
 wire sw_273_scan_out;
 wire sw_274_clk_out;
 wire sw_274_data_out;
 wire sw_274_latch_out;
 wire \sw_274_module_data_in[0] ;
 wire \sw_274_module_data_in[1] ;
 wire \sw_274_module_data_in[2] ;
 wire \sw_274_module_data_in[3] ;
 wire \sw_274_module_data_in[4] ;
 wire \sw_274_module_data_in[5] ;
 wire \sw_274_module_data_in[6] ;
 wire \sw_274_module_data_in[7] ;
 wire \sw_274_module_data_out[0] ;
 wire \sw_274_module_data_out[1] ;
 wire \sw_274_module_data_out[2] ;
 wire \sw_274_module_data_out[3] ;
 wire \sw_274_module_data_out[4] ;
 wire \sw_274_module_data_out[5] ;
 wire \sw_274_module_data_out[6] ;
 wire \sw_274_module_data_out[7] ;
 wire sw_274_scan_out;
 wire sw_275_clk_out;
 wire sw_275_data_out;
 wire sw_275_latch_out;
 wire \sw_275_module_data_in[0] ;
 wire \sw_275_module_data_in[1] ;
 wire \sw_275_module_data_in[2] ;
 wire \sw_275_module_data_in[3] ;
 wire \sw_275_module_data_in[4] ;
 wire \sw_275_module_data_in[5] ;
 wire \sw_275_module_data_in[6] ;
 wire \sw_275_module_data_in[7] ;
 wire \sw_275_module_data_out[0] ;
 wire \sw_275_module_data_out[1] ;
 wire \sw_275_module_data_out[2] ;
 wire \sw_275_module_data_out[3] ;
 wire \sw_275_module_data_out[4] ;
 wire \sw_275_module_data_out[5] ;
 wire \sw_275_module_data_out[6] ;
 wire \sw_275_module_data_out[7] ;
 wire sw_275_scan_out;
 wire sw_276_clk_out;
 wire sw_276_data_out;
 wire sw_276_latch_out;
 wire \sw_276_module_data_in[0] ;
 wire \sw_276_module_data_in[1] ;
 wire \sw_276_module_data_in[2] ;
 wire \sw_276_module_data_in[3] ;
 wire \sw_276_module_data_in[4] ;
 wire \sw_276_module_data_in[5] ;
 wire \sw_276_module_data_in[6] ;
 wire \sw_276_module_data_in[7] ;
 wire \sw_276_module_data_out[0] ;
 wire \sw_276_module_data_out[1] ;
 wire \sw_276_module_data_out[2] ;
 wire \sw_276_module_data_out[3] ;
 wire \sw_276_module_data_out[4] ;
 wire \sw_276_module_data_out[5] ;
 wire \sw_276_module_data_out[6] ;
 wire \sw_276_module_data_out[7] ;
 wire sw_276_scan_out;
 wire sw_277_clk_out;
 wire sw_277_data_out;
 wire sw_277_latch_out;
 wire \sw_277_module_data_in[0] ;
 wire \sw_277_module_data_in[1] ;
 wire \sw_277_module_data_in[2] ;
 wire \sw_277_module_data_in[3] ;
 wire \sw_277_module_data_in[4] ;
 wire \sw_277_module_data_in[5] ;
 wire \sw_277_module_data_in[6] ;
 wire \sw_277_module_data_in[7] ;
 wire \sw_277_module_data_out[0] ;
 wire \sw_277_module_data_out[1] ;
 wire \sw_277_module_data_out[2] ;
 wire \sw_277_module_data_out[3] ;
 wire \sw_277_module_data_out[4] ;
 wire \sw_277_module_data_out[5] ;
 wire \sw_277_module_data_out[6] ;
 wire \sw_277_module_data_out[7] ;
 wire sw_277_scan_out;
 wire sw_278_clk_out;
 wire sw_278_data_out;
 wire sw_278_latch_out;
 wire \sw_278_module_data_in[0] ;
 wire \sw_278_module_data_in[1] ;
 wire \sw_278_module_data_in[2] ;
 wire \sw_278_module_data_in[3] ;
 wire \sw_278_module_data_in[4] ;
 wire \sw_278_module_data_in[5] ;
 wire \sw_278_module_data_in[6] ;
 wire \sw_278_module_data_in[7] ;
 wire \sw_278_module_data_out[0] ;
 wire \sw_278_module_data_out[1] ;
 wire \sw_278_module_data_out[2] ;
 wire \sw_278_module_data_out[3] ;
 wire \sw_278_module_data_out[4] ;
 wire \sw_278_module_data_out[5] ;
 wire \sw_278_module_data_out[6] ;
 wire \sw_278_module_data_out[7] ;
 wire sw_278_scan_out;
 wire sw_279_clk_out;
 wire sw_279_data_out;
 wire sw_279_latch_out;
 wire \sw_279_module_data_in[0] ;
 wire \sw_279_module_data_in[1] ;
 wire \sw_279_module_data_in[2] ;
 wire \sw_279_module_data_in[3] ;
 wire \sw_279_module_data_in[4] ;
 wire \sw_279_module_data_in[5] ;
 wire \sw_279_module_data_in[6] ;
 wire \sw_279_module_data_in[7] ;
 wire \sw_279_module_data_out[0] ;
 wire \sw_279_module_data_out[1] ;
 wire \sw_279_module_data_out[2] ;
 wire \sw_279_module_data_out[3] ;
 wire \sw_279_module_data_out[4] ;
 wire \sw_279_module_data_out[5] ;
 wire \sw_279_module_data_out[6] ;
 wire \sw_279_module_data_out[7] ;
 wire sw_279_scan_out;
 wire sw_280_clk_out;
 wire sw_280_data_out;
 wire sw_280_latch_out;
 wire \sw_280_module_data_in[0] ;
 wire \sw_280_module_data_in[1] ;
 wire \sw_280_module_data_in[2] ;
 wire \sw_280_module_data_in[3] ;
 wire \sw_280_module_data_in[4] ;
 wire \sw_280_module_data_in[5] ;
 wire \sw_280_module_data_in[6] ;
 wire \sw_280_module_data_in[7] ;
 wire \sw_280_module_data_out[0] ;
 wire \sw_280_module_data_out[1] ;
 wire \sw_280_module_data_out[2] ;
 wire \sw_280_module_data_out[3] ;
 wire \sw_280_module_data_out[4] ;
 wire \sw_280_module_data_out[5] ;
 wire \sw_280_module_data_out[6] ;
 wire \sw_280_module_data_out[7] ;
 wire sw_280_scan_out;
 wire sw_281_clk_out;
 wire sw_281_data_out;
 wire sw_281_latch_out;
 wire \sw_281_module_data_in[0] ;
 wire \sw_281_module_data_in[1] ;
 wire \sw_281_module_data_in[2] ;
 wire \sw_281_module_data_in[3] ;
 wire \sw_281_module_data_in[4] ;
 wire \sw_281_module_data_in[5] ;
 wire \sw_281_module_data_in[6] ;
 wire \sw_281_module_data_in[7] ;
 wire \sw_281_module_data_out[0] ;
 wire \sw_281_module_data_out[1] ;
 wire \sw_281_module_data_out[2] ;
 wire \sw_281_module_data_out[3] ;
 wire \sw_281_module_data_out[4] ;
 wire \sw_281_module_data_out[5] ;
 wire \sw_281_module_data_out[6] ;
 wire \sw_281_module_data_out[7] ;
 wire sw_281_scan_out;
 wire sw_282_clk_out;
 wire sw_282_data_out;
 wire sw_282_latch_out;
 wire \sw_282_module_data_in[0] ;
 wire \sw_282_module_data_in[1] ;
 wire \sw_282_module_data_in[2] ;
 wire \sw_282_module_data_in[3] ;
 wire \sw_282_module_data_in[4] ;
 wire \sw_282_module_data_in[5] ;
 wire \sw_282_module_data_in[6] ;
 wire \sw_282_module_data_in[7] ;
 wire \sw_282_module_data_out[0] ;
 wire \sw_282_module_data_out[1] ;
 wire \sw_282_module_data_out[2] ;
 wire \sw_282_module_data_out[3] ;
 wire \sw_282_module_data_out[4] ;
 wire \sw_282_module_data_out[5] ;
 wire \sw_282_module_data_out[6] ;
 wire \sw_282_module_data_out[7] ;
 wire sw_282_scan_out;
 wire sw_283_clk_out;
 wire sw_283_data_out;
 wire sw_283_latch_out;
 wire \sw_283_module_data_in[0] ;
 wire \sw_283_module_data_in[1] ;
 wire \sw_283_module_data_in[2] ;
 wire \sw_283_module_data_in[3] ;
 wire \sw_283_module_data_in[4] ;
 wire \sw_283_module_data_in[5] ;
 wire \sw_283_module_data_in[6] ;
 wire \sw_283_module_data_in[7] ;
 wire \sw_283_module_data_out[0] ;
 wire \sw_283_module_data_out[1] ;
 wire \sw_283_module_data_out[2] ;
 wire \sw_283_module_data_out[3] ;
 wire \sw_283_module_data_out[4] ;
 wire \sw_283_module_data_out[5] ;
 wire \sw_283_module_data_out[6] ;
 wire \sw_283_module_data_out[7] ;
 wire sw_283_scan_out;
 wire sw_284_clk_out;
 wire sw_284_data_out;
 wire sw_284_latch_out;
 wire \sw_284_module_data_in[0] ;
 wire \sw_284_module_data_in[1] ;
 wire \sw_284_module_data_in[2] ;
 wire \sw_284_module_data_in[3] ;
 wire \sw_284_module_data_in[4] ;
 wire \sw_284_module_data_in[5] ;
 wire \sw_284_module_data_in[6] ;
 wire \sw_284_module_data_in[7] ;
 wire \sw_284_module_data_out[0] ;
 wire \sw_284_module_data_out[1] ;
 wire \sw_284_module_data_out[2] ;
 wire \sw_284_module_data_out[3] ;
 wire \sw_284_module_data_out[4] ;
 wire \sw_284_module_data_out[5] ;
 wire \sw_284_module_data_out[6] ;
 wire \sw_284_module_data_out[7] ;
 wire sw_284_scan_out;
 wire sw_285_clk_out;
 wire sw_285_data_out;
 wire sw_285_latch_out;
 wire \sw_285_module_data_in[0] ;
 wire \sw_285_module_data_in[1] ;
 wire \sw_285_module_data_in[2] ;
 wire \sw_285_module_data_in[3] ;
 wire \sw_285_module_data_in[4] ;
 wire \sw_285_module_data_in[5] ;
 wire \sw_285_module_data_in[6] ;
 wire \sw_285_module_data_in[7] ;
 wire \sw_285_module_data_out[0] ;
 wire \sw_285_module_data_out[1] ;
 wire \sw_285_module_data_out[2] ;
 wire \sw_285_module_data_out[3] ;
 wire \sw_285_module_data_out[4] ;
 wire \sw_285_module_data_out[5] ;
 wire \sw_285_module_data_out[6] ;
 wire \sw_285_module_data_out[7] ;
 wire sw_285_scan_out;
 wire sw_286_clk_out;
 wire sw_286_data_out;
 wire sw_286_latch_out;
 wire \sw_286_module_data_in[0] ;
 wire \sw_286_module_data_in[1] ;
 wire \sw_286_module_data_in[2] ;
 wire \sw_286_module_data_in[3] ;
 wire \sw_286_module_data_in[4] ;
 wire \sw_286_module_data_in[5] ;
 wire \sw_286_module_data_in[6] ;
 wire \sw_286_module_data_in[7] ;
 wire \sw_286_module_data_out[0] ;
 wire \sw_286_module_data_out[1] ;
 wire \sw_286_module_data_out[2] ;
 wire \sw_286_module_data_out[3] ;
 wire \sw_286_module_data_out[4] ;
 wire \sw_286_module_data_out[5] ;
 wire \sw_286_module_data_out[6] ;
 wire \sw_286_module_data_out[7] ;
 wire sw_286_scan_out;
 wire sw_287_clk_out;
 wire sw_287_data_out;
 wire sw_287_latch_out;
 wire \sw_287_module_data_in[0] ;
 wire \sw_287_module_data_in[1] ;
 wire \sw_287_module_data_in[2] ;
 wire \sw_287_module_data_in[3] ;
 wire \sw_287_module_data_in[4] ;
 wire \sw_287_module_data_in[5] ;
 wire \sw_287_module_data_in[6] ;
 wire \sw_287_module_data_in[7] ;
 wire \sw_287_module_data_out[0] ;
 wire \sw_287_module_data_out[1] ;
 wire \sw_287_module_data_out[2] ;
 wire \sw_287_module_data_out[3] ;
 wire \sw_287_module_data_out[4] ;
 wire \sw_287_module_data_out[5] ;
 wire \sw_287_module_data_out[6] ;
 wire \sw_287_module_data_out[7] ;
 wire sw_287_scan_out;
 wire sw_288_clk_out;
 wire sw_288_data_out;
 wire sw_288_latch_out;
 wire \sw_288_module_data_in[0] ;
 wire \sw_288_module_data_in[1] ;
 wire \sw_288_module_data_in[2] ;
 wire \sw_288_module_data_in[3] ;
 wire \sw_288_module_data_in[4] ;
 wire \sw_288_module_data_in[5] ;
 wire \sw_288_module_data_in[6] ;
 wire \sw_288_module_data_in[7] ;
 wire \sw_288_module_data_out[0] ;
 wire \sw_288_module_data_out[1] ;
 wire \sw_288_module_data_out[2] ;
 wire \sw_288_module_data_out[3] ;
 wire \sw_288_module_data_out[4] ;
 wire \sw_288_module_data_out[5] ;
 wire \sw_288_module_data_out[6] ;
 wire \sw_288_module_data_out[7] ;
 wire sw_288_scan_out;
 wire sw_289_clk_out;
 wire sw_289_data_out;
 wire sw_289_latch_out;
 wire \sw_289_module_data_in[0] ;
 wire \sw_289_module_data_in[1] ;
 wire \sw_289_module_data_in[2] ;
 wire \sw_289_module_data_in[3] ;
 wire \sw_289_module_data_in[4] ;
 wire \sw_289_module_data_in[5] ;
 wire \sw_289_module_data_in[6] ;
 wire \sw_289_module_data_in[7] ;
 wire \sw_289_module_data_out[0] ;
 wire \sw_289_module_data_out[1] ;
 wire \sw_289_module_data_out[2] ;
 wire \sw_289_module_data_out[3] ;
 wire \sw_289_module_data_out[4] ;
 wire \sw_289_module_data_out[5] ;
 wire \sw_289_module_data_out[6] ;
 wire \sw_289_module_data_out[7] ;
 wire sw_289_scan_out;
 wire sw_290_clk_out;
 wire sw_290_data_out;
 wire sw_290_latch_out;
 wire \sw_290_module_data_in[0] ;
 wire \sw_290_module_data_in[1] ;
 wire \sw_290_module_data_in[2] ;
 wire \sw_290_module_data_in[3] ;
 wire \sw_290_module_data_in[4] ;
 wire \sw_290_module_data_in[5] ;
 wire \sw_290_module_data_in[6] ;
 wire \sw_290_module_data_in[7] ;
 wire \sw_290_module_data_out[0] ;
 wire \sw_290_module_data_out[1] ;
 wire \sw_290_module_data_out[2] ;
 wire \sw_290_module_data_out[3] ;
 wire \sw_290_module_data_out[4] ;
 wire \sw_290_module_data_out[5] ;
 wire \sw_290_module_data_out[6] ;
 wire \sw_290_module_data_out[7] ;
 wire sw_290_scan_out;
 wire sw_291_clk_out;
 wire sw_291_data_out;
 wire sw_291_latch_out;
 wire \sw_291_module_data_in[0] ;
 wire \sw_291_module_data_in[1] ;
 wire \sw_291_module_data_in[2] ;
 wire \sw_291_module_data_in[3] ;
 wire \sw_291_module_data_in[4] ;
 wire \sw_291_module_data_in[5] ;
 wire \sw_291_module_data_in[6] ;
 wire \sw_291_module_data_in[7] ;
 wire \sw_291_module_data_out[0] ;
 wire \sw_291_module_data_out[1] ;
 wire \sw_291_module_data_out[2] ;
 wire \sw_291_module_data_out[3] ;
 wire \sw_291_module_data_out[4] ;
 wire \sw_291_module_data_out[5] ;
 wire \sw_291_module_data_out[6] ;
 wire \sw_291_module_data_out[7] ;
 wire sw_291_scan_out;
 wire sw_292_clk_out;
 wire sw_292_data_out;
 wire sw_292_latch_out;
 wire \sw_292_module_data_in[0] ;
 wire \sw_292_module_data_in[1] ;
 wire \sw_292_module_data_in[2] ;
 wire \sw_292_module_data_in[3] ;
 wire \sw_292_module_data_in[4] ;
 wire \sw_292_module_data_in[5] ;
 wire \sw_292_module_data_in[6] ;
 wire \sw_292_module_data_in[7] ;
 wire \sw_292_module_data_out[0] ;
 wire \sw_292_module_data_out[1] ;
 wire \sw_292_module_data_out[2] ;
 wire \sw_292_module_data_out[3] ;
 wire \sw_292_module_data_out[4] ;
 wire \sw_292_module_data_out[5] ;
 wire \sw_292_module_data_out[6] ;
 wire \sw_292_module_data_out[7] ;
 wire sw_292_scan_out;
 wire sw_293_clk_out;
 wire sw_293_data_out;
 wire sw_293_latch_out;
 wire \sw_293_module_data_in[0] ;
 wire \sw_293_module_data_in[1] ;
 wire \sw_293_module_data_in[2] ;
 wire \sw_293_module_data_in[3] ;
 wire \sw_293_module_data_in[4] ;
 wire \sw_293_module_data_in[5] ;
 wire \sw_293_module_data_in[6] ;
 wire \sw_293_module_data_in[7] ;
 wire \sw_293_module_data_out[0] ;
 wire \sw_293_module_data_out[1] ;
 wire \sw_293_module_data_out[2] ;
 wire \sw_293_module_data_out[3] ;
 wire \sw_293_module_data_out[4] ;
 wire \sw_293_module_data_out[5] ;
 wire \sw_293_module_data_out[6] ;
 wire \sw_293_module_data_out[7] ;
 wire sw_293_scan_out;
 wire sw_294_clk_out;
 wire sw_294_data_out;
 wire sw_294_latch_out;
 wire \sw_294_module_data_in[0] ;
 wire \sw_294_module_data_in[1] ;
 wire \sw_294_module_data_in[2] ;
 wire \sw_294_module_data_in[3] ;
 wire \sw_294_module_data_in[4] ;
 wire \sw_294_module_data_in[5] ;
 wire \sw_294_module_data_in[6] ;
 wire \sw_294_module_data_in[7] ;
 wire \sw_294_module_data_out[0] ;
 wire \sw_294_module_data_out[1] ;
 wire \sw_294_module_data_out[2] ;
 wire \sw_294_module_data_out[3] ;
 wire \sw_294_module_data_out[4] ;
 wire \sw_294_module_data_out[5] ;
 wire \sw_294_module_data_out[6] ;
 wire \sw_294_module_data_out[7] ;
 wire sw_294_scan_out;
 wire sw_295_clk_out;
 wire sw_295_data_out;
 wire sw_295_latch_out;
 wire \sw_295_module_data_in[0] ;
 wire \sw_295_module_data_in[1] ;
 wire \sw_295_module_data_in[2] ;
 wire \sw_295_module_data_in[3] ;
 wire \sw_295_module_data_in[4] ;
 wire \sw_295_module_data_in[5] ;
 wire \sw_295_module_data_in[6] ;
 wire \sw_295_module_data_in[7] ;
 wire \sw_295_module_data_out[0] ;
 wire \sw_295_module_data_out[1] ;
 wire \sw_295_module_data_out[2] ;
 wire \sw_295_module_data_out[3] ;
 wire \sw_295_module_data_out[4] ;
 wire \sw_295_module_data_out[5] ;
 wire \sw_295_module_data_out[6] ;
 wire \sw_295_module_data_out[7] ;
 wire sw_295_scan_out;
 wire sw_296_clk_out;
 wire sw_296_data_out;
 wire sw_296_latch_out;
 wire \sw_296_module_data_in[0] ;
 wire \sw_296_module_data_in[1] ;
 wire \sw_296_module_data_in[2] ;
 wire \sw_296_module_data_in[3] ;
 wire \sw_296_module_data_in[4] ;
 wire \sw_296_module_data_in[5] ;
 wire \sw_296_module_data_in[6] ;
 wire \sw_296_module_data_in[7] ;
 wire \sw_296_module_data_out[0] ;
 wire \sw_296_module_data_out[1] ;
 wire \sw_296_module_data_out[2] ;
 wire \sw_296_module_data_out[3] ;
 wire \sw_296_module_data_out[4] ;
 wire \sw_296_module_data_out[5] ;
 wire \sw_296_module_data_out[6] ;
 wire \sw_296_module_data_out[7] ;
 wire sw_296_scan_out;
 wire sw_297_clk_out;
 wire sw_297_data_out;
 wire sw_297_latch_out;
 wire \sw_297_module_data_in[0] ;
 wire \sw_297_module_data_in[1] ;
 wire \sw_297_module_data_in[2] ;
 wire \sw_297_module_data_in[3] ;
 wire \sw_297_module_data_in[4] ;
 wire \sw_297_module_data_in[5] ;
 wire \sw_297_module_data_in[6] ;
 wire \sw_297_module_data_in[7] ;
 wire \sw_297_module_data_out[0] ;
 wire \sw_297_module_data_out[1] ;
 wire \sw_297_module_data_out[2] ;
 wire \sw_297_module_data_out[3] ;
 wire \sw_297_module_data_out[4] ;
 wire \sw_297_module_data_out[5] ;
 wire \sw_297_module_data_out[6] ;
 wire \sw_297_module_data_out[7] ;
 wire sw_297_scan_out;
 wire sw_298_clk_out;
 wire sw_298_data_out;
 wire sw_298_latch_out;
 wire \sw_298_module_data_in[0] ;
 wire \sw_298_module_data_in[1] ;
 wire \sw_298_module_data_in[2] ;
 wire \sw_298_module_data_in[3] ;
 wire \sw_298_module_data_in[4] ;
 wire \sw_298_module_data_in[5] ;
 wire \sw_298_module_data_in[6] ;
 wire \sw_298_module_data_in[7] ;
 wire \sw_298_module_data_out[0] ;
 wire \sw_298_module_data_out[1] ;
 wire \sw_298_module_data_out[2] ;
 wire \sw_298_module_data_out[3] ;
 wire \sw_298_module_data_out[4] ;
 wire \sw_298_module_data_out[5] ;
 wire \sw_298_module_data_out[6] ;
 wire \sw_298_module_data_out[7] ;
 wire sw_298_scan_out;
 wire sw_299_clk_out;
 wire sw_299_data_out;
 wire sw_299_latch_out;
 wire \sw_299_module_data_in[0] ;
 wire \sw_299_module_data_in[1] ;
 wire \sw_299_module_data_in[2] ;
 wire \sw_299_module_data_in[3] ;
 wire \sw_299_module_data_in[4] ;
 wire \sw_299_module_data_in[5] ;
 wire \sw_299_module_data_in[6] ;
 wire \sw_299_module_data_in[7] ;
 wire \sw_299_module_data_out[0] ;
 wire \sw_299_module_data_out[1] ;
 wire \sw_299_module_data_out[2] ;
 wire \sw_299_module_data_out[3] ;
 wire \sw_299_module_data_out[4] ;
 wire \sw_299_module_data_out[5] ;
 wire \sw_299_module_data_out[6] ;
 wire \sw_299_module_data_out[7] ;
 wire sw_299_scan_out;
 wire sw_300_clk_out;
 wire sw_300_data_out;
 wire sw_300_latch_out;
 wire \sw_300_module_data_in[0] ;
 wire \sw_300_module_data_in[1] ;
 wire \sw_300_module_data_in[2] ;
 wire \sw_300_module_data_in[3] ;
 wire \sw_300_module_data_in[4] ;
 wire \sw_300_module_data_in[5] ;
 wire \sw_300_module_data_in[6] ;
 wire \sw_300_module_data_in[7] ;
 wire \sw_300_module_data_out[0] ;
 wire \sw_300_module_data_out[1] ;
 wire \sw_300_module_data_out[2] ;
 wire \sw_300_module_data_out[3] ;
 wire \sw_300_module_data_out[4] ;
 wire \sw_300_module_data_out[5] ;
 wire \sw_300_module_data_out[6] ;
 wire \sw_300_module_data_out[7] ;
 wire sw_300_scan_out;
 wire sw_301_clk_out;
 wire sw_301_data_out;
 wire sw_301_latch_out;
 wire \sw_301_module_data_in[0] ;
 wire \sw_301_module_data_in[1] ;
 wire \sw_301_module_data_in[2] ;
 wire \sw_301_module_data_in[3] ;
 wire \sw_301_module_data_in[4] ;
 wire \sw_301_module_data_in[5] ;
 wire \sw_301_module_data_in[6] ;
 wire \sw_301_module_data_in[7] ;
 wire \sw_301_module_data_out[0] ;
 wire \sw_301_module_data_out[1] ;
 wire \sw_301_module_data_out[2] ;
 wire \sw_301_module_data_out[3] ;
 wire \sw_301_module_data_out[4] ;
 wire \sw_301_module_data_out[5] ;
 wire \sw_301_module_data_out[6] ;
 wire \sw_301_module_data_out[7] ;
 wire sw_301_scan_out;
 wire sw_302_clk_out;
 wire sw_302_data_out;
 wire sw_302_latch_out;
 wire \sw_302_module_data_in[0] ;
 wire \sw_302_module_data_in[1] ;
 wire \sw_302_module_data_in[2] ;
 wire \sw_302_module_data_in[3] ;
 wire \sw_302_module_data_in[4] ;
 wire \sw_302_module_data_in[5] ;
 wire \sw_302_module_data_in[6] ;
 wire \sw_302_module_data_in[7] ;
 wire \sw_302_module_data_out[0] ;
 wire \sw_302_module_data_out[1] ;
 wire \sw_302_module_data_out[2] ;
 wire \sw_302_module_data_out[3] ;
 wire \sw_302_module_data_out[4] ;
 wire \sw_302_module_data_out[5] ;
 wire \sw_302_module_data_out[6] ;
 wire \sw_302_module_data_out[7] ;
 wire sw_302_scan_out;
 wire sw_303_clk_out;
 wire sw_303_data_out;
 wire sw_303_latch_out;
 wire \sw_303_module_data_in[0] ;
 wire \sw_303_module_data_in[1] ;
 wire \sw_303_module_data_in[2] ;
 wire \sw_303_module_data_in[3] ;
 wire \sw_303_module_data_in[4] ;
 wire \sw_303_module_data_in[5] ;
 wire \sw_303_module_data_in[6] ;
 wire \sw_303_module_data_in[7] ;
 wire \sw_303_module_data_out[0] ;
 wire \sw_303_module_data_out[1] ;
 wire \sw_303_module_data_out[2] ;
 wire \sw_303_module_data_out[3] ;
 wire \sw_303_module_data_out[4] ;
 wire \sw_303_module_data_out[5] ;
 wire \sw_303_module_data_out[6] ;
 wire \sw_303_module_data_out[7] ;
 wire sw_303_scan_out;
 wire sw_304_clk_out;
 wire sw_304_data_out;
 wire sw_304_latch_out;
 wire \sw_304_module_data_in[0] ;
 wire \sw_304_module_data_in[1] ;
 wire \sw_304_module_data_in[2] ;
 wire \sw_304_module_data_in[3] ;
 wire \sw_304_module_data_in[4] ;
 wire \sw_304_module_data_in[5] ;
 wire \sw_304_module_data_in[6] ;
 wire \sw_304_module_data_in[7] ;
 wire \sw_304_module_data_out[0] ;
 wire \sw_304_module_data_out[1] ;
 wire \sw_304_module_data_out[2] ;
 wire \sw_304_module_data_out[3] ;
 wire \sw_304_module_data_out[4] ;
 wire \sw_304_module_data_out[5] ;
 wire \sw_304_module_data_out[6] ;
 wire \sw_304_module_data_out[7] ;
 wire sw_304_scan_out;
 wire sw_305_clk_out;
 wire sw_305_data_out;
 wire sw_305_latch_out;
 wire \sw_305_module_data_in[0] ;
 wire \sw_305_module_data_in[1] ;
 wire \sw_305_module_data_in[2] ;
 wire \sw_305_module_data_in[3] ;
 wire \sw_305_module_data_in[4] ;
 wire \sw_305_module_data_in[5] ;
 wire \sw_305_module_data_in[6] ;
 wire \sw_305_module_data_in[7] ;
 wire \sw_305_module_data_out[0] ;
 wire \sw_305_module_data_out[1] ;
 wire \sw_305_module_data_out[2] ;
 wire \sw_305_module_data_out[3] ;
 wire \sw_305_module_data_out[4] ;
 wire \sw_305_module_data_out[5] ;
 wire \sw_305_module_data_out[6] ;
 wire \sw_305_module_data_out[7] ;
 wire sw_305_scan_out;
 wire sw_306_clk_out;
 wire sw_306_data_out;
 wire sw_306_latch_out;
 wire \sw_306_module_data_in[0] ;
 wire \sw_306_module_data_in[1] ;
 wire \sw_306_module_data_in[2] ;
 wire \sw_306_module_data_in[3] ;
 wire \sw_306_module_data_in[4] ;
 wire \sw_306_module_data_in[5] ;
 wire \sw_306_module_data_in[6] ;
 wire \sw_306_module_data_in[7] ;
 wire \sw_306_module_data_out[0] ;
 wire \sw_306_module_data_out[1] ;
 wire \sw_306_module_data_out[2] ;
 wire \sw_306_module_data_out[3] ;
 wire \sw_306_module_data_out[4] ;
 wire \sw_306_module_data_out[5] ;
 wire \sw_306_module_data_out[6] ;
 wire \sw_306_module_data_out[7] ;
 wire sw_306_scan_out;
 wire sw_307_clk_out;
 wire sw_307_data_out;
 wire sw_307_latch_out;
 wire \sw_307_module_data_in[0] ;
 wire \sw_307_module_data_in[1] ;
 wire \sw_307_module_data_in[2] ;
 wire \sw_307_module_data_in[3] ;
 wire \sw_307_module_data_in[4] ;
 wire \sw_307_module_data_in[5] ;
 wire \sw_307_module_data_in[6] ;
 wire \sw_307_module_data_in[7] ;
 wire \sw_307_module_data_out[0] ;
 wire \sw_307_module_data_out[1] ;
 wire \sw_307_module_data_out[2] ;
 wire \sw_307_module_data_out[3] ;
 wire \sw_307_module_data_out[4] ;
 wire \sw_307_module_data_out[5] ;
 wire \sw_307_module_data_out[6] ;
 wire \sw_307_module_data_out[7] ;
 wire sw_307_scan_out;
 wire sw_308_clk_out;
 wire sw_308_data_out;
 wire sw_308_latch_out;
 wire \sw_308_module_data_in[0] ;
 wire \sw_308_module_data_in[1] ;
 wire \sw_308_module_data_in[2] ;
 wire \sw_308_module_data_in[3] ;
 wire \sw_308_module_data_in[4] ;
 wire \sw_308_module_data_in[5] ;
 wire \sw_308_module_data_in[6] ;
 wire \sw_308_module_data_in[7] ;
 wire \sw_308_module_data_out[0] ;
 wire \sw_308_module_data_out[1] ;
 wire \sw_308_module_data_out[2] ;
 wire \sw_308_module_data_out[3] ;
 wire \sw_308_module_data_out[4] ;
 wire \sw_308_module_data_out[5] ;
 wire \sw_308_module_data_out[6] ;
 wire \sw_308_module_data_out[7] ;
 wire sw_308_scan_out;
 wire sw_309_clk_out;
 wire sw_309_data_out;
 wire sw_309_latch_out;
 wire \sw_309_module_data_in[0] ;
 wire \sw_309_module_data_in[1] ;
 wire \sw_309_module_data_in[2] ;
 wire \sw_309_module_data_in[3] ;
 wire \sw_309_module_data_in[4] ;
 wire \sw_309_module_data_in[5] ;
 wire \sw_309_module_data_in[6] ;
 wire \sw_309_module_data_in[7] ;
 wire \sw_309_module_data_out[0] ;
 wire \sw_309_module_data_out[1] ;
 wire \sw_309_module_data_out[2] ;
 wire \sw_309_module_data_out[3] ;
 wire \sw_309_module_data_out[4] ;
 wire \sw_309_module_data_out[5] ;
 wire \sw_309_module_data_out[6] ;
 wire \sw_309_module_data_out[7] ;
 wire sw_309_scan_out;
 wire sw_310_clk_out;
 wire sw_310_data_out;
 wire sw_310_latch_out;
 wire \sw_310_module_data_in[0] ;
 wire \sw_310_module_data_in[1] ;
 wire \sw_310_module_data_in[2] ;
 wire \sw_310_module_data_in[3] ;
 wire \sw_310_module_data_in[4] ;
 wire \sw_310_module_data_in[5] ;
 wire \sw_310_module_data_in[6] ;
 wire \sw_310_module_data_in[7] ;
 wire \sw_310_module_data_out[0] ;
 wire \sw_310_module_data_out[1] ;
 wire \sw_310_module_data_out[2] ;
 wire \sw_310_module_data_out[3] ;
 wire \sw_310_module_data_out[4] ;
 wire \sw_310_module_data_out[5] ;
 wire \sw_310_module_data_out[6] ;
 wire \sw_310_module_data_out[7] ;
 wire sw_310_scan_out;
 wire sw_311_clk_out;
 wire sw_311_data_out;
 wire sw_311_latch_out;
 wire \sw_311_module_data_in[0] ;
 wire \sw_311_module_data_in[1] ;
 wire \sw_311_module_data_in[2] ;
 wire \sw_311_module_data_in[3] ;
 wire \sw_311_module_data_in[4] ;
 wire \sw_311_module_data_in[5] ;
 wire \sw_311_module_data_in[6] ;
 wire \sw_311_module_data_in[7] ;
 wire \sw_311_module_data_out[0] ;
 wire \sw_311_module_data_out[1] ;
 wire \sw_311_module_data_out[2] ;
 wire \sw_311_module_data_out[3] ;
 wire \sw_311_module_data_out[4] ;
 wire \sw_311_module_data_out[5] ;
 wire \sw_311_module_data_out[6] ;
 wire \sw_311_module_data_out[7] ;
 wire sw_311_scan_out;
 wire sw_312_clk_out;
 wire sw_312_data_out;
 wire sw_312_latch_out;
 wire \sw_312_module_data_in[0] ;
 wire \sw_312_module_data_in[1] ;
 wire \sw_312_module_data_in[2] ;
 wire \sw_312_module_data_in[3] ;
 wire \sw_312_module_data_in[4] ;
 wire \sw_312_module_data_in[5] ;
 wire \sw_312_module_data_in[6] ;
 wire \sw_312_module_data_in[7] ;
 wire \sw_312_module_data_out[0] ;
 wire \sw_312_module_data_out[1] ;
 wire \sw_312_module_data_out[2] ;
 wire \sw_312_module_data_out[3] ;
 wire \sw_312_module_data_out[4] ;
 wire \sw_312_module_data_out[5] ;
 wire \sw_312_module_data_out[6] ;
 wire \sw_312_module_data_out[7] ;
 wire sw_312_scan_out;
 wire sw_313_clk_out;
 wire sw_313_data_out;
 wire sw_313_latch_out;
 wire \sw_313_module_data_in[0] ;
 wire \sw_313_module_data_in[1] ;
 wire \sw_313_module_data_in[2] ;
 wire \sw_313_module_data_in[3] ;
 wire \sw_313_module_data_in[4] ;
 wire \sw_313_module_data_in[5] ;
 wire \sw_313_module_data_in[6] ;
 wire \sw_313_module_data_in[7] ;
 wire \sw_313_module_data_out[0] ;
 wire \sw_313_module_data_out[1] ;
 wire \sw_313_module_data_out[2] ;
 wire \sw_313_module_data_out[3] ;
 wire \sw_313_module_data_out[4] ;
 wire \sw_313_module_data_out[5] ;
 wire \sw_313_module_data_out[6] ;
 wire \sw_313_module_data_out[7] ;
 wire sw_313_scan_out;
 wire sw_314_clk_out;
 wire sw_314_data_out;
 wire sw_314_latch_out;
 wire \sw_314_module_data_in[0] ;
 wire \sw_314_module_data_in[1] ;
 wire \sw_314_module_data_in[2] ;
 wire \sw_314_module_data_in[3] ;
 wire \sw_314_module_data_in[4] ;
 wire \sw_314_module_data_in[5] ;
 wire \sw_314_module_data_in[6] ;
 wire \sw_314_module_data_in[7] ;
 wire \sw_314_module_data_out[0] ;
 wire \sw_314_module_data_out[1] ;
 wire \sw_314_module_data_out[2] ;
 wire \sw_314_module_data_out[3] ;
 wire \sw_314_module_data_out[4] ;
 wire \sw_314_module_data_out[5] ;
 wire \sw_314_module_data_out[6] ;
 wire \sw_314_module_data_out[7] ;
 wire sw_314_scan_out;
 wire sw_315_clk_out;
 wire sw_315_data_out;
 wire sw_315_latch_out;
 wire \sw_315_module_data_in[0] ;
 wire \sw_315_module_data_in[1] ;
 wire \sw_315_module_data_in[2] ;
 wire \sw_315_module_data_in[3] ;
 wire \sw_315_module_data_in[4] ;
 wire \sw_315_module_data_in[5] ;
 wire \sw_315_module_data_in[6] ;
 wire \sw_315_module_data_in[7] ;
 wire \sw_315_module_data_out[0] ;
 wire \sw_315_module_data_out[1] ;
 wire \sw_315_module_data_out[2] ;
 wire \sw_315_module_data_out[3] ;
 wire \sw_315_module_data_out[4] ;
 wire \sw_315_module_data_out[5] ;
 wire \sw_315_module_data_out[6] ;
 wire \sw_315_module_data_out[7] ;
 wire sw_315_scan_out;
 wire sw_316_clk_out;
 wire sw_316_data_out;
 wire sw_316_latch_out;
 wire \sw_316_module_data_in[0] ;
 wire \sw_316_module_data_in[1] ;
 wire \sw_316_module_data_in[2] ;
 wire \sw_316_module_data_in[3] ;
 wire \sw_316_module_data_in[4] ;
 wire \sw_316_module_data_in[5] ;
 wire \sw_316_module_data_in[6] ;
 wire \sw_316_module_data_in[7] ;
 wire \sw_316_module_data_out[0] ;
 wire \sw_316_module_data_out[1] ;
 wire \sw_316_module_data_out[2] ;
 wire \sw_316_module_data_out[3] ;
 wire \sw_316_module_data_out[4] ;
 wire \sw_316_module_data_out[5] ;
 wire \sw_316_module_data_out[6] ;
 wire \sw_316_module_data_out[7] ;
 wire sw_316_scan_out;
 wire sw_317_clk_out;
 wire sw_317_data_out;
 wire sw_317_latch_out;
 wire \sw_317_module_data_in[0] ;
 wire \sw_317_module_data_in[1] ;
 wire \sw_317_module_data_in[2] ;
 wire \sw_317_module_data_in[3] ;
 wire \sw_317_module_data_in[4] ;
 wire \sw_317_module_data_in[5] ;
 wire \sw_317_module_data_in[6] ;
 wire \sw_317_module_data_in[7] ;
 wire \sw_317_module_data_out[0] ;
 wire \sw_317_module_data_out[1] ;
 wire \sw_317_module_data_out[2] ;
 wire \sw_317_module_data_out[3] ;
 wire \sw_317_module_data_out[4] ;
 wire \sw_317_module_data_out[5] ;
 wire \sw_317_module_data_out[6] ;
 wire \sw_317_module_data_out[7] ;
 wire sw_317_scan_out;
 wire sw_318_clk_out;
 wire sw_318_data_out;
 wire sw_318_latch_out;
 wire \sw_318_module_data_in[0] ;
 wire \sw_318_module_data_in[1] ;
 wire \sw_318_module_data_in[2] ;
 wire \sw_318_module_data_in[3] ;
 wire \sw_318_module_data_in[4] ;
 wire \sw_318_module_data_in[5] ;
 wire \sw_318_module_data_in[6] ;
 wire \sw_318_module_data_in[7] ;
 wire \sw_318_module_data_out[0] ;
 wire \sw_318_module_data_out[1] ;
 wire \sw_318_module_data_out[2] ;
 wire \sw_318_module_data_out[3] ;
 wire \sw_318_module_data_out[4] ;
 wire \sw_318_module_data_out[5] ;
 wire \sw_318_module_data_out[6] ;
 wire \sw_318_module_data_out[7] ;
 wire sw_318_scan_out;
 wire sw_319_clk_out;
 wire sw_319_data_out;
 wire sw_319_latch_out;
 wire \sw_319_module_data_in[0] ;
 wire \sw_319_module_data_in[1] ;
 wire \sw_319_module_data_in[2] ;
 wire \sw_319_module_data_in[3] ;
 wire \sw_319_module_data_in[4] ;
 wire \sw_319_module_data_in[5] ;
 wire \sw_319_module_data_in[6] ;
 wire \sw_319_module_data_in[7] ;
 wire \sw_319_module_data_out[0] ;
 wire \sw_319_module_data_out[1] ;
 wire \sw_319_module_data_out[2] ;
 wire \sw_319_module_data_out[3] ;
 wire \sw_319_module_data_out[4] ;
 wire \sw_319_module_data_out[5] ;
 wire \sw_319_module_data_out[6] ;
 wire \sw_319_module_data_out[7] ;
 wire sw_319_scan_out;
 wire sw_320_clk_out;
 wire sw_320_data_out;
 wire sw_320_latch_out;
 wire \sw_320_module_data_in[0] ;
 wire \sw_320_module_data_in[1] ;
 wire \sw_320_module_data_in[2] ;
 wire \sw_320_module_data_in[3] ;
 wire \sw_320_module_data_in[4] ;
 wire \sw_320_module_data_in[5] ;
 wire \sw_320_module_data_in[6] ;
 wire \sw_320_module_data_in[7] ;
 wire \sw_320_module_data_out[0] ;
 wire \sw_320_module_data_out[1] ;
 wire \sw_320_module_data_out[2] ;
 wire \sw_320_module_data_out[3] ;
 wire \sw_320_module_data_out[4] ;
 wire \sw_320_module_data_out[5] ;
 wire \sw_320_module_data_out[6] ;
 wire \sw_320_module_data_out[7] ;
 wire sw_320_scan_out;
 wire sw_321_clk_out;
 wire sw_321_data_out;
 wire sw_321_latch_out;
 wire \sw_321_module_data_in[0] ;
 wire \sw_321_module_data_in[1] ;
 wire \sw_321_module_data_in[2] ;
 wire \sw_321_module_data_in[3] ;
 wire \sw_321_module_data_in[4] ;
 wire \sw_321_module_data_in[5] ;
 wire \sw_321_module_data_in[6] ;
 wire \sw_321_module_data_in[7] ;
 wire \sw_321_module_data_out[0] ;
 wire \sw_321_module_data_out[1] ;
 wire \sw_321_module_data_out[2] ;
 wire \sw_321_module_data_out[3] ;
 wire \sw_321_module_data_out[4] ;
 wire \sw_321_module_data_out[5] ;
 wire \sw_321_module_data_out[6] ;
 wire \sw_321_module_data_out[7] ;
 wire sw_321_scan_out;
 wire sw_322_clk_out;
 wire sw_322_data_out;
 wire sw_322_latch_out;
 wire \sw_322_module_data_in[0] ;
 wire \sw_322_module_data_in[1] ;
 wire \sw_322_module_data_in[2] ;
 wire \sw_322_module_data_in[3] ;
 wire \sw_322_module_data_in[4] ;
 wire \sw_322_module_data_in[5] ;
 wire \sw_322_module_data_in[6] ;
 wire \sw_322_module_data_in[7] ;
 wire \sw_322_module_data_out[0] ;
 wire \sw_322_module_data_out[1] ;
 wire \sw_322_module_data_out[2] ;
 wire \sw_322_module_data_out[3] ;
 wire \sw_322_module_data_out[4] ;
 wire \sw_322_module_data_out[5] ;
 wire \sw_322_module_data_out[6] ;
 wire \sw_322_module_data_out[7] ;
 wire sw_322_scan_out;
 wire sw_323_clk_out;
 wire sw_323_data_out;
 wire sw_323_latch_out;
 wire \sw_323_module_data_in[0] ;
 wire \sw_323_module_data_in[1] ;
 wire \sw_323_module_data_in[2] ;
 wire \sw_323_module_data_in[3] ;
 wire \sw_323_module_data_in[4] ;
 wire \sw_323_module_data_in[5] ;
 wire \sw_323_module_data_in[6] ;
 wire \sw_323_module_data_in[7] ;
 wire \sw_323_module_data_out[0] ;
 wire \sw_323_module_data_out[1] ;
 wire \sw_323_module_data_out[2] ;
 wire \sw_323_module_data_out[3] ;
 wire \sw_323_module_data_out[4] ;
 wire \sw_323_module_data_out[5] ;
 wire \sw_323_module_data_out[6] ;
 wire \sw_323_module_data_out[7] ;
 wire sw_323_scan_out;
 wire sw_324_clk_out;
 wire sw_324_data_out;
 wire sw_324_latch_out;
 wire \sw_324_module_data_in[0] ;
 wire \sw_324_module_data_in[1] ;
 wire \sw_324_module_data_in[2] ;
 wire \sw_324_module_data_in[3] ;
 wire \sw_324_module_data_in[4] ;
 wire \sw_324_module_data_in[5] ;
 wire \sw_324_module_data_in[6] ;
 wire \sw_324_module_data_in[7] ;
 wire \sw_324_module_data_out[0] ;
 wire \sw_324_module_data_out[1] ;
 wire \sw_324_module_data_out[2] ;
 wire \sw_324_module_data_out[3] ;
 wire \sw_324_module_data_out[4] ;
 wire \sw_324_module_data_out[5] ;
 wire \sw_324_module_data_out[6] ;
 wire \sw_324_module_data_out[7] ;
 wire sw_324_scan_out;
 wire sw_325_clk_out;
 wire sw_325_data_out;
 wire sw_325_latch_out;
 wire \sw_325_module_data_in[0] ;
 wire \sw_325_module_data_in[1] ;
 wire \sw_325_module_data_in[2] ;
 wire \sw_325_module_data_in[3] ;
 wire \sw_325_module_data_in[4] ;
 wire \sw_325_module_data_in[5] ;
 wire \sw_325_module_data_in[6] ;
 wire \sw_325_module_data_in[7] ;
 wire \sw_325_module_data_out[0] ;
 wire \sw_325_module_data_out[1] ;
 wire \sw_325_module_data_out[2] ;
 wire \sw_325_module_data_out[3] ;
 wire \sw_325_module_data_out[4] ;
 wire \sw_325_module_data_out[5] ;
 wire \sw_325_module_data_out[6] ;
 wire \sw_325_module_data_out[7] ;
 wire sw_325_scan_out;
 wire sw_326_clk_out;
 wire sw_326_data_out;
 wire sw_326_latch_out;
 wire \sw_326_module_data_in[0] ;
 wire \sw_326_module_data_in[1] ;
 wire \sw_326_module_data_in[2] ;
 wire \sw_326_module_data_in[3] ;
 wire \sw_326_module_data_in[4] ;
 wire \sw_326_module_data_in[5] ;
 wire \sw_326_module_data_in[6] ;
 wire \sw_326_module_data_in[7] ;
 wire \sw_326_module_data_out[0] ;
 wire \sw_326_module_data_out[1] ;
 wire \sw_326_module_data_out[2] ;
 wire \sw_326_module_data_out[3] ;
 wire \sw_326_module_data_out[4] ;
 wire \sw_326_module_data_out[5] ;
 wire \sw_326_module_data_out[6] ;
 wire \sw_326_module_data_out[7] ;
 wire sw_326_scan_out;
 wire sw_327_clk_out;
 wire sw_327_data_out;
 wire sw_327_latch_out;
 wire \sw_327_module_data_in[0] ;
 wire \sw_327_module_data_in[1] ;
 wire \sw_327_module_data_in[2] ;
 wire \sw_327_module_data_in[3] ;
 wire \sw_327_module_data_in[4] ;
 wire \sw_327_module_data_in[5] ;
 wire \sw_327_module_data_in[6] ;
 wire \sw_327_module_data_in[7] ;
 wire \sw_327_module_data_out[0] ;
 wire \sw_327_module_data_out[1] ;
 wire \sw_327_module_data_out[2] ;
 wire \sw_327_module_data_out[3] ;
 wire \sw_327_module_data_out[4] ;
 wire \sw_327_module_data_out[5] ;
 wire \sw_327_module_data_out[6] ;
 wire \sw_327_module_data_out[7] ;
 wire sw_327_scan_out;
 wire sw_328_clk_out;
 wire sw_328_data_out;
 wire sw_328_latch_out;
 wire \sw_328_module_data_in[0] ;
 wire \sw_328_module_data_in[1] ;
 wire \sw_328_module_data_in[2] ;
 wire \sw_328_module_data_in[3] ;
 wire \sw_328_module_data_in[4] ;
 wire \sw_328_module_data_in[5] ;
 wire \sw_328_module_data_in[6] ;
 wire \sw_328_module_data_in[7] ;
 wire \sw_328_module_data_out[0] ;
 wire \sw_328_module_data_out[1] ;
 wire \sw_328_module_data_out[2] ;
 wire \sw_328_module_data_out[3] ;
 wire \sw_328_module_data_out[4] ;
 wire \sw_328_module_data_out[5] ;
 wire \sw_328_module_data_out[6] ;
 wire \sw_328_module_data_out[7] ;
 wire sw_328_scan_out;
 wire sw_329_clk_out;
 wire sw_329_data_out;
 wire sw_329_latch_out;
 wire \sw_329_module_data_in[0] ;
 wire \sw_329_module_data_in[1] ;
 wire \sw_329_module_data_in[2] ;
 wire \sw_329_module_data_in[3] ;
 wire \sw_329_module_data_in[4] ;
 wire \sw_329_module_data_in[5] ;
 wire \sw_329_module_data_in[6] ;
 wire \sw_329_module_data_in[7] ;
 wire \sw_329_module_data_out[0] ;
 wire \sw_329_module_data_out[1] ;
 wire \sw_329_module_data_out[2] ;
 wire \sw_329_module_data_out[3] ;
 wire \sw_329_module_data_out[4] ;
 wire \sw_329_module_data_out[5] ;
 wire \sw_329_module_data_out[6] ;
 wire \sw_329_module_data_out[7] ;
 wire sw_329_scan_out;
 wire sw_330_clk_out;
 wire sw_330_data_out;
 wire sw_330_latch_out;
 wire \sw_330_module_data_in[0] ;
 wire \sw_330_module_data_in[1] ;
 wire \sw_330_module_data_in[2] ;
 wire \sw_330_module_data_in[3] ;
 wire \sw_330_module_data_in[4] ;
 wire \sw_330_module_data_in[5] ;
 wire \sw_330_module_data_in[6] ;
 wire \sw_330_module_data_in[7] ;
 wire \sw_330_module_data_out[0] ;
 wire \sw_330_module_data_out[1] ;
 wire \sw_330_module_data_out[2] ;
 wire \sw_330_module_data_out[3] ;
 wire \sw_330_module_data_out[4] ;
 wire \sw_330_module_data_out[5] ;
 wire \sw_330_module_data_out[6] ;
 wire \sw_330_module_data_out[7] ;
 wire sw_330_scan_out;
 wire sw_331_clk_out;
 wire sw_331_data_out;
 wire sw_331_latch_out;
 wire \sw_331_module_data_in[0] ;
 wire \sw_331_module_data_in[1] ;
 wire \sw_331_module_data_in[2] ;
 wire \sw_331_module_data_in[3] ;
 wire \sw_331_module_data_in[4] ;
 wire \sw_331_module_data_in[5] ;
 wire \sw_331_module_data_in[6] ;
 wire \sw_331_module_data_in[7] ;
 wire \sw_331_module_data_out[0] ;
 wire \sw_331_module_data_out[1] ;
 wire \sw_331_module_data_out[2] ;
 wire \sw_331_module_data_out[3] ;
 wire \sw_331_module_data_out[4] ;
 wire \sw_331_module_data_out[5] ;
 wire \sw_331_module_data_out[6] ;
 wire \sw_331_module_data_out[7] ;
 wire sw_331_scan_out;
 wire sw_332_clk_out;
 wire sw_332_data_out;
 wire sw_332_latch_out;
 wire \sw_332_module_data_in[0] ;
 wire \sw_332_module_data_in[1] ;
 wire \sw_332_module_data_in[2] ;
 wire \sw_332_module_data_in[3] ;
 wire \sw_332_module_data_in[4] ;
 wire \sw_332_module_data_in[5] ;
 wire \sw_332_module_data_in[6] ;
 wire \sw_332_module_data_in[7] ;
 wire \sw_332_module_data_out[0] ;
 wire \sw_332_module_data_out[1] ;
 wire \sw_332_module_data_out[2] ;
 wire \sw_332_module_data_out[3] ;
 wire \sw_332_module_data_out[4] ;
 wire \sw_332_module_data_out[5] ;
 wire \sw_332_module_data_out[6] ;
 wire \sw_332_module_data_out[7] ;
 wire sw_332_scan_out;
 wire sw_333_clk_out;
 wire sw_333_data_out;
 wire sw_333_latch_out;
 wire \sw_333_module_data_in[0] ;
 wire \sw_333_module_data_in[1] ;
 wire \sw_333_module_data_in[2] ;
 wire \sw_333_module_data_in[3] ;
 wire \sw_333_module_data_in[4] ;
 wire \sw_333_module_data_in[5] ;
 wire \sw_333_module_data_in[6] ;
 wire \sw_333_module_data_in[7] ;
 wire \sw_333_module_data_out[0] ;
 wire \sw_333_module_data_out[1] ;
 wire \sw_333_module_data_out[2] ;
 wire \sw_333_module_data_out[3] ;
 wire \sw_333_module_data_out[4] ;
 wire \sw_333_module_data_out[5] ;
 wire \sw_333_module_data_out[6] ;
 wire \sw_333_module_data_out[7] ;
 wire sw_333_scan_out;
 wire sw_334_clk_out;
 wire sw_334_data_out;
 wire sw_334_latch_out;
 wire \sw_334_module_data_in[0] ;
 wire \sw_334_module_data_in[1] ;
 wire \sw_334_module_data_in[2] ;
 wire \sw_334_module_data_in[3] ;
 wire \sw_334_module_data_in[4] ;
 wire \sw_334_module_data_in[5] ;
 wire \sw_334_module_data_in[6] ;
 wire \sw_334_module_data_in[7] ;
 wire \sw_334_module_data_out[0] ;
 wire \sw_334_module_data_out[1] ;
 wire \sw_334_module_data_out[2] ;
 wire \sw_334_module_data_out[3] ;
 wire \sw_334_module_data_out[4] ;
 wire \sw_334_module_data_out[5] ;
 wire \sw_334_module_data_out[6] ;
 wire \sw_334_module_data_out[7] ;
 wire sw_334_scan_out;
 wire sw_335_clk_out;
 wire sw_335_data_out;
 wire sw_335_latch_out;
 wire \sw_335_module_data_in[0] ;
 wire \sw_335_module_data_in[1] ;
 wire \sw_335_module_data_in[2] ;
 wire \sw_335_module_data_in[3] ;
 wire \sw_335_module_data_in[4] ;
 wire \sw_335_module_data_in[5] ;
 wire \sw_335_module_data_in[6] ;
 wire \sw_335_module_data_in[7] ;
 wire \sw_335_module_data_out[0] ;
 wire \sw_335_module_data_out[1] ;
 wire \sw_335_module_data_out[2] ;
 wire \sw_335_module_data_out[3] ;
 wire \sw_335_module_data_out[4] ;
 wire \sw_335_module_data_out[5] ;
 wire \sw_335_module_data_out[6] ;
 wire \sw_335_module_data_out[7] ;
 wire sw_335_scan_out;
 wire sw_336_clk_out;
 wire sw_336_data_out;
 wire sw_336_latch_out;
 wire \sw_336_module_data_in[0] ;
 wire \sw_336_module_data_in[1] ;
 wire \sw_336_module_data_in[2] ;
 wire \sw_336_module_data_in[3] ;
 wire \sw_336_module_data_in[4] ;
 wire \sw_336_module_data_in[5] ;
 wire \sw_336_module_data_in[6] ;
 wire \sw_336_module_data_in[7] ;
 wire \sw_336_module_data_out[0] ;
 wire \sw_336_module_data_out[1] ;
 wire \sw_336_module_data_out[2] ;
 wire \sw_336_module_data_out[3] ;
 wire \sw_336_module_data_out[4] ;
 wire \sw_336_module_data_out[5] ;
 wire \sw_336_module_data_out[6] ;
 wire \sw_336_module_data_out[7] ;
 wire sw_336_scan_out;
 wire sw_337_clk_out;
 wire sw_337_data_out;
 wire sw_337_latch_out;
 wire \sw_337_module_data_in[0] ;
 wire \sw_337_module_data_in[1] ;
 wire \sw_337_module_data_in[2] ;
 wire \sw_337_module_data_in[3] ;
 wire \sw_337_module_data_in[4] ;
 wire \sw_337_module_data_in[5] ;
 wire \sw_337_module_data_in[6] ;
 wire \sw_337_module_data_in[7] ;
 wire \sw_337_module_data_out[0] ;
 wire \sw_337_module_data_out[1] ;
 wire \sw_337_module_data_out[2] ;
 wire \sw_337_module_data_out[3] ;
 wire \sw_337_module_data_out[4] ;
 wire \sw_337_module_data_out[5] ;
 wire \sw_337_module_data_out[6] ;
 wire \sw_337_module_data_out[7] ;
 wire sw_337_scan_out;
 wire sw_338_clk_out;
 wire sw_338_data_out;
 wire sw_338_latch_out;
 wire \sw_338_module_data_in[0] ;
 wire \sw_338_module_data_in[1] ;
 wire \sw_338_module_data_in[2] ;
 wire \sw_338_module_data_in[3] ;
 wire \sw_338_module_data_in[4] ;
 wire \sw_338_module_data_in[5] ;
 wire \sw_338_module_data_in[6] ;
 wire \sw_338_module_data_in[7] ;
 wire \sw_338_module_data_out[0] ;
 wire \sw_338_module_data_out[1] ;
 wire \sw_338_module_data_out[2] ;
 wire \sw_338_module_data_out[3] ;
 wire \sw_338_module_data_out[4] ;
 wire \sw_338_module_data_out[5] ;
 wire \sw_338_module_data_out[6] ;
 wire \sw_338_module_data_out[7] ;
 wire sw_338_scan_out;
 wire sw_339_clk_out;
 wire sw_339_data_out;
 wire sw_339_latch_out;
 wire \sw_339_module_data_in[0] ;
 wire \sw_339_module_data_in[1] ;
 wire \sw_339_module_data_in[2] ;
 wire \sw_339_module_data_in[3] ;
 wire \sw_339_module_data_in[4] ;
 wire \sw_339_module_data_in[5] ;
 wire \sw_339_module_data_in[6] ;
 wire \sw_339_module_data_in[7] ;
 wire \sw_339_module_data_out[0] ;
 wire \sw_339_module_data_out[1] ;
 wire \sw_339_module_data_out[2] ;
 wire \sw_339_module_data_out[3] ;
 wire \sw_339_module_data_out[4] ;
 wire \sw_339_module_data_out[5] ;
 wire \sw_339_module_data_out[6] ;
 wire \sw_339_module_data_out[7] ;
 wire sw_339_scan_out;
 wire sw_340_clk_out;
 wire sw_340_data_out;
 wire sw_340_latch_out;
 wire \sw_340_module_data_in[0] ;
 wire \sw_340_module_data_in[1] ;
 wire \sw_340_module_data_in[2] ;
 wire \sw_340_module_data_in[3] ;
 wire \sw_340_module_data_in[4] ;
 wire \sw_340_module_data_in[5] ;
 wire \sw_340_module_data_in[6] ;
 wire \sw_340_module_data_in[7] ;
 wire \sw_340_module_data_out[0] ;
 wire \sw_340_module_data_out[1] ;
 wire \sw_340_module_data_out[2] ;
 wire \sw_340_module_data_out[3] ;
 wire \sw_340_module_data_out[4] ;
 wire \sw_340_module_data_out[5] ;
 wire \sw_340_module_data_out[6] ;
 wire \sw_340_module_data_out[7] ;
 wire sw_340_scan_out;
 wire sw_341_clk_out;
 wire sw_341_data_out;
 wire sw_341_latch_out;
 wire \sw_341_module_data_in[0] ;
 wire \sw_341_module_data_in[1] ;
 wire \sw_341_module_data_in[2] ;
 wire \sw_341_module_data_in[3] ;
 wire \sw_341_module_data_in[4] ;
 wire \sw_341_module_data_in[5] ;
 wire \sw_341_module_data_in[6] ;
 wire \sw_341_module_data_in[7] ;
 wire \sw_341_module_data_out[0] ;
 wire \sw_341_module_data_out[1] ;
 wire \sw_341_module_data_out[2] ;
 wire \sw_341_module_data_out[3] ;
 wire \sw_341_module_data_out[4] ;
 wire \sw_341_module_data_out[5] ;
 wire \sw_341_module_data_out[6] ;
 wire \sw_341_module_data_out[7] ;
 wire sw_341_scan_out;
 wire sw_342_clk_out;
 wire sw_342_data_out;
 wire sw_342_latch_out;
 wire \sw_342_module_data_in[0] ;
 wire \sw_342_module_data_in[1] ;
 wire \sw_342_module_data_in[2] ;
 wire \sw_342_module_data_in[3] ;
 wire \sw_342_module_data_in[4] ;
 wire \sw_342_module_data_in[5] ;
 wire \sw_342_module_data_in[6] ;
 wire \sw_342_module_data_in[7] ;
 wire \sw_342_module_data_out[0] ;
 wire \sw_342_module_data_out[1] ;
 wire \sw_342_module_data_out[2] ;
 wire \sw_342_module_data_out[3] ;
 wire \sw_342_module_data_out[4] ;
 wire \sw_342_module_data_out[5] ;
 wire \sw_342_module_data_out[6] ;
 wire \sw_342_module_data_out[7] ;
 wire sw_342_scan_out;
 wire sw_343_clk_out;
 wire sw_343_data_out;
 wire sw_343_latch_out;
 wire \sw_343_module_data_in[0] ;
 wire \sw_343_module_data_in[1] ;
 wire \sw_343_module_data_in[2] ;
 wire \sw_343_module_data_in[3] ;
 wire \sw_343_module_data_in[4] ;
 wire \sw_343_module_data_in[5] ;
 wire \sw_343_module_data_in[6] ;
 wire \sw_343_module_data_in[7] ;
 wire \sw_343_module_data_out[0] ;
 wire \sw_343_module_data_out[1] ;
 wire \sw_343_module_data_out[2] ;
 wire \sw_343_module_data_out[3] ;
 wire \sw_343_module_data_out[4] ;
 wire \sw_343_module_data_out[5] ;
 wire \sw_343_module_data_out[6] ;
 wire \sw_343_module_data_out[7] ;
 wire sw_343_scan_out;
 wire sw_344_clk_out;
 wire sw_344_data_out;
 wire sw_344_latch_out;
 wire \sw_344_module_data_in[0] ;
 wire \sw_344_module_data_in[1] ;
 wire \sw_344_module_data_in[2] ;
 wire \sw_344_module_data_in[3] ;
 wire \sw_344_module_data_in[4] ;
 wire \sw_344_module_data_in[5] ;
 wire \sw_344_module_data_in[6] ;
 wire \sw_344_module_data_in[7] ;
 wire \sw_344_module_data_out[0] ;
 wire \sw_344_module_data_out[1] ;
 wire \sw_344_module_data_out[2] ;
 wire \sw_344_module_data_out[3] ;
 wire \sw_344_module_data_out[4] ;
 wire \sw_344_module_data_out[5] ;
 wire \sw_344_module_data_out[6] ;
 wire \sw_344_module_data_out[7] ;
 wire sw_344_scan_out;
 wire sw_345_clk_out;
 wire sw_345_data_out;
 wire sw_345_latch_out;
 wire \sw_345_module_data_in[0] ;
 wire \sw_345_module_data_in[1] ;
 wire \sw_345_module_data_in[2] ;
 wire \sw_345_module_data_in[3] ;
 wire \sw_345_module_data_in[4] ;
 wire \sw_345_module_data_in[5] ;
 wire \sw_345_module_data_in[6] ;
 wire \sw_345_module_data_in[7] ;
 wire \sw_345_module_data_out[0] ;
 wire \sw_345_module_data_out[1] ;
 wire \sw_345_module_data_out[2] ;
 wire \sw_345_module_data_out[3] ;
 wire \sw_345_module_data_out[4] ;
 wire \sw_345_module_data_out[5] ;
 wire \sw_345_module_data_out[6] ;
 wire \sw_345_module_data_out[7] ;
 wire sw_345_scan_out;
 wire sw_346_clk_out;
 wire sw_346_data_out;
 wire sw_346_latch_out;
 wire \sw_346_module_data_in[0] ;
 wire \sw_346_module_data_in[1] ;
 wire \sw_346_module_data_in[2] ;
 wire \sw_346_module_data_in[3] ;
 wire \sw_346_module_data_in[4] ;
 wire \sw_346_module_data_in[5] ;
 wire \sw_346_module_data_in[6] ;
 wire \sw_346_module_data_in[7] ;
 wire \sw_346_module_data_out[0] ;
 wire \sw_346_module_data_out[1] ;
 wire \sw_346_module_data_out[2] ;
 wire \sw_346_module_data_out[3] ;
 wire \sw_346_module_data_out[4] ;
 wire \sw_346_module_data_out[5] ;
 wire \sw_346_module_data_out[6] ;
 wire \sw_346_module_data_out[7] ;
 wire sw_346_scan_out;
 wire sw_347_clk_out;
 wire sw_347_data_out;
 wire sw_347_latch_out;
 wire \sw_347_module_data_in[0] ;
 wire \sw_347_module_data_in[1] ;
 wire \sw_347_module_data_in[2] ;
 wire \sw_347_module_data_in[3] ;
 wire \sw_347_module_data_in[4] ;
 wire \sw_347_module_data_in[5] ;
 wire \sw_347_module_data_in[6] ;
 wire \sw_347_module_data_in[7] ;
 wire \sw_347_module_data_out[0] ;
 wire \sw_347_module_data_out[1] ;
 wire \sw_347_module_data_out[2] ;
 wire \sw_347_module_data_out[3] ;
 wire \sw_347_module_data_out[4] ;
 wire \sw_347_module_data_out[5] ;
 wire \sw_347_module_data_out[6] ;
 wire \sw_347_module_data_out[7] ;
 wire sw_347_scan_out;
 wire sw_348_clk_out;
 wire sw_348_data_out;
 wire sw_348_latch_out;
 wire \sw_348_module_data_in[0] ;
 wire \sw_348_module_data_in[1] ;
 wire \sw_348_module_data_in[2] ;
 wire \sw_348_module_data_in[3] ;
 wire \sw_348_module_data_in[4] ;
 wire \sw_348_module_data_in[5] ;
 wire \sw_348_module_data_in[6] ;
 wire \sw_348_module_data_in[7] ;
 wire \sw_348_module_data_out[0] ;
 wire \sw_348_module_data_out[1] ;
 wire \sw_348_module_data_out[2] ;
 wire \sw_348_module_data_out[3] ;
 wire \sw_348_module_data_out[4] ;
 wire \sw_348_module_data_out[5] ;
 wire \sw_348_module_data_out[6] ;
 wire \sw_348_module_data_out[7] ;
 wire sw_348_scan_out;
 wire sw_349_clk_out;
 wire sw_349_data_out;
 wire sw_349_latch_out;
 wire \sw_349_module_data_in[0] ;
 wire \sw_349_module_data_in[1] ;
 wire \sw_349_module_data_in[2] ;
 wire \sw_349_module_data_in[3] ;
 wire \sw_349_module_data_in[4] ;
 wire \sw_349_module_data_in[5] ;
 wire \sw_349_module_data_in[6] ;
 wire \sw_349_module_data_in[7] ;
 wire \sw_349_module_data_out[0] ;
 wire \sw_349_module_data_out[1] ;
 wire \sw_349_module_data_out[2] ;
 wire \sw_349_module_data_out[3] ;
 wire \sw_349_module_data_out[4] ;
 wire \sw_349_module_data_out[5] ;
 wire \sw_349_module_data_out[6] ;
 wire \sw_349_module_data_out[7] ;
 wire sw_349_scan_out;
 wire sw_350_clk_out;
 wire sw_350_data_out;
 wire sw_350_latch_out;
 wire \sw_350_module_data_in[0] ;
 wire \sw_350_module_data_in[1] ;
 wire \sw_350_module_data_in[2] ;
 wire \sw_350_module_data_in[3] ;
 wire \sw_350_module_data_in[4] ;
 wire \sw_350_module_data_in[5] ;
 wire \sw_350_module_data_in[6] ;
 wire \sw_350_module_data_in[7] ;
 wire \sw_350_module_data_out[0] ;
 wire \sw_350_module_data_out[1] ;
 wire \sw_350_module_data_out[2] ;
 wire \sw_350_module_data_out[3] ;
 wire \sw_350_module_data_out[4] ;
 wire \sw_350_module_data_out[5] ;
 wire \sw_350_module_data_out[6] ;
 wire \sw_350_module_data_out[7] ;
 wire sw_350_scan_out;
 wire sw_351_clk_out;
 wire sw_351_data_out;
 wire sw_351_latch_out;
 wire \sw_351_module_data_in[0] ;
 wire \sw_351_module_data_in[1] ;
 wire \sw_351_module_data_in[2] ;
 wire \sw_351_module_data_in[3] ;
 wire \sw_351_module_data_in[4] ;
 wire \sw_351_module_data_in[5] ;
 wire \sw_351_module_data_in[6] ;
 wire \sw_351_module_data_in[7] ;
 wire \sw_351_module_data_out[0] ;
 wire \sw_351_module_data_out[1] ;
 wire \sw_351_module_data_out[2] ;
 wire \sw_351_module_data_out[3] ;
 wire \sw_351_module_data_out[4] ;
 wire \sw_351_module_data_out[5] ;
 wire \sw_351_module_data_out[6] ;
 wire \sw_351_module_data_out[7] ;
 wire sw_351_scan_out;
 wire sw_352_clk_out;
 wire sw_352_data_out;
 wire sw_352_latch_out;
 wire \sw_352_module_data_in[0] ;
 wire \sw_352_module_data_in[1] ;
 wire \sw_352_module_data_in[2] ;
 wire \sw_352_module_data_in[3] ;
 wire \sw_352_module_data_in[4] ;
 wire \sw_352_module_data_in[5] ;
 wire \sw_352_module_data_in[6] ;
 wire \sw_352_module_data_in[7] ;
 wire \sw_352_module_data_out[0] ;
 wire \sw_352_module_data_out[1] ;
 wire \sw_352_module_data_out[2] ;
 wire \sw_352_module_data_out[3] ;
 wire \sw_352_module_data_out[4] ;
 wire \sw_352_module_data_out[5] ;
 wire \sw_352_module_data_out[6] ;
 wire \sw_352_module_data_out[7] ;
 wire sw_352_scan_out;
 wire sw_353_clk_out;
 wire sw_353_data_out;
 wire sw_353_latch_out;
 wire \sw_353_module_data_in[0] ;
 wire \sw_353_module_data_in[1] ;
 wire \sw_353_module_data_in[2] ;
 wire \sw_353_module_data_in[3] ;
 wire \sw_353_module_data_in[4] ;
 wire \sw_353_module_data_in[5] ;
 wire \sw_353_module_data_in[6] ;
 wire \sw_353_module_data_in[7] ;
 wire \sw_353_module_data_out[0] ;
 wire \sw_353_module_data_out[1] ;
 wire \sw_353_module_data_out[2] ;
 wire \sw_353_module_data_out[3] ;
 wire \sw_353_module_data_out[4] ;
 wire \sw_353_module_data_out[5] ;
 wire \sw_353_module_data_out[6] ;
 wire \sw_353_module_data_out[7] ;
 wire sw_353_scan_out;
 wire sw_354_clk_out;
 wire sw_354_data_out;
 wire sw_354_latch_out;
 wire \sw_354_module_data_in[0] ;
 wire \sw_354_module_data_in[1] ;
 wire \sw_354_module_data_in[2] ;
 wire \sw_354_module_data_in[3] ;
 wire \sw_354_module_data_in[4] ;
 wire \sw_354_module_data_in[5] ;
 wire \sw_354_module_data_in[6] ;
 wire \sw_354_module_data_in[7] ;
 wire \sw_354_module_data_out[0] ;
 wire \sw_354_module_data_out[1] ;
 wire \sw_354_module_data_out[2] ;
 wire \sw_354_module_data_out[3] ;
 wire \sw_354_module_data_out[4] ;
 wire \sw_354_module_data_out[5] ;
 wire \sw_354_module_data_out[6] ;
 wire \sw_354_module_data_out[7] ;
 wire sw_354_scan_out;
 wire sw_355_clk_out;
 wire sw_355_data_out;
 wire sw_355_latch_out;
 wire \sw_355_module_data_in[0] ;
 wire \sw_355_module_data_in[1] ;
 wire \sw_355_module_data_in[2] ;
 wire \sw_355_module_data_in[3] ;
 wire \sw_355_module_data_in[4] ;
 wire \sw_355_module_data_in[5] ;
 wire \sw_355_module_data_in[6] ;
 wire \sw_355_module_data_in[7] ;
 wire \sw_355_module_data_out[0] ;
 wire \sw_355_module_data_out[1] ;
 wire \sw_355_module_data_out[2] ;
 wire \sw_355_module_data_out[3] ;
 wire \sw_355_module_data_out[4] ;
 wire \sw_355_module_data_out[5] ;
 wire \sw_355_module_data_out[6] ;
 wire \sw_355_module_data_out[7] ;
 wire sw_355_scan_out;
 wire sw_356_clk_out;
 wire sw_356_data_out;
 wire sw_356_latch_out;
 wire \sw_356_module_data_in[0] ;
 wire \sw_356_module_data_in[1] ;
 wire \sw_356_module_data_in[2] ;
 wire \sw_356_module_data_in[3] ;
 wire \sw_356_module_data_in[4] ;
 wire \sw_356_module_data_in[5] ;
 wire \sw_356_module_data_in[6] ;
 wire \sw_356_module_data_in[7] ;
 wire \sw_356_module_data_out[0] ;
 wire \sw_356_module_data_out[1] ;
 wire \sw_356_module_data_out[2] ;
 wire \sw_356_module_data_out[3] ;
 wire \sw_356_module_data_out[4] ;
 wire \sw_356_module_data_out[5] ;
 wire \sw_356_module_data_out[6] ;
 wire \sw_356_module_data_out[7] ;
 wire sw_356_scan_out;
 wire sw_357_clk_out;
 wire sw_357_data_out;
 wire sw_357_latch_out;
 wire \sw_357_module_data_in[0] ;
 wire \sw_357_module_data_in[1] ;
 wire \sw_357_module_data_in[2] ;
 wire \sw_357_module_data_in[3] ;
 wire \sw_357_module_data_in[4] ;
 wire \sw_357_module_data_in[5] ;
 wire \sw_357_module_data_in[6] ;
 wire \sw_357_module_data_in[7] ;
 wire \sw_357_module_data_out[0] ;
 wire \sw_357_module_data_out[1] ;
 wire \sw_357_module_data_out[2] ;
 wire \sw_357_module_data_out[3] ;
 wire \sw_357_module_data_out[4] ;
 wire \sw_357_module_data_out[5] ;
 wire \sw_357_module_data_out[6] ;
 wire \sw_357_module_data_out[7] ;
 wire sw_357_scan_out;
 wire sw_358_clk_out;
 wire sw_358_data_out;
 wire sw_358_latch_out;
 wire \sw_358_module_data_in[0] ;
 wire \sw_358_module_data_in[1] ;
 wire \sw_358_module_data_in[2] ;
 wire \sw_358_module_data_in[3] ;
 wire \sw_358_module_data_in[4] ;
 wire \sw_358_module_data_in[5] ;
 wire \sw_358_module_data_in[6] ;
 wire \sw_358_module_data_in[7] ;
 wire \sw_358_module_data_out[0] ;
 wire \sw_358_module_data_out[1] ;
 wire \sw_358_module_data_out[2] ;
 wire \sw_358_module_data_out[3] ;
 wire \sw_358_module_data_out[4] ;
 wire \sw_358_module_data_out[5] ;
 wire \sw_358_module_data_out[6] ;
 wire \sw_358_module_data_out[7] ;
 wire sw_358_scan_out;
 wire sw_359_clk_out;
 wire sw_359_data_out;
 wire sw_359_latch_out;
 wire \sw_359_module_data_in[0] ;
 wire \sw_359_module_data_in[1] ;
 wire \sw_359_module_data_in[2] ;
 wire \sw_359_module_data_in[3] ;
 wire \sw_359_module_data_in[4] ;
 wire \sw_359_module_data_in[5] ;
 wire \sw_359_module_data_in[6] ;
 wire \sw_359_module_data_in[7] ;
 wire \sw_359_module_data_out[0] ;
 wire \sw_359_module_data_out[1] ;
 wire \sw_359_module_data_out[2] ;
 wire \sw_359_module_data_out[3] ;
 wire \sw_359_module_data_out[4] ;
 wire \sw_359_module_data_out[5] ;
 wire \sw_359_module_data_out[6] ;
 wire \sw_359_module_data_out[7] ;
 wire sw_359_scan_out;
 wire sw_360_clk_out;
 wire sw_360_data_out;
 wire sw_360_latch_out;
 wire \sw_360_module_data_in[0] ;
 wire \sw_360_module_data_in[1] ;
 wire \sw_360_module_data_in[2] ;
 wire \sw_360_module_data_in[3] ;
 wire \sw_360_module_data_in[4] ;
 wire \sw_360_module_data_in[5] ;
 wire \sw_360_module_data_in[6] ;
 wire \sw_360_module_data_in[7] ;
 wire \sw_360_module_data_out[0] ;
 wire \sw_360_module_data_out[1] ;
 wire \sw_360_module_data_out[2] ;
 wire \sw_360_module_data_out[3] ;
 wire \sw_360_module_data_out[4] ;
 wire \sw_360_module_data_out[5] ;
 wire \sw_360_module_data_out[6] ;
 wire \sw_360_module_data_out[7] ;
 wire sw_360_scan_out;
 wire sw_361_clk_out;
 wire sw_361_data_out;
 wire sw_361_latch_out;
 wire \sw_361_module_data_in[0] ;
 wire \sw_361_module_data_in[1] ;
 wire \sw_361_module_data_in[2] ;
 wire \sw_361_module_data_in[3] ;
 wire \sw_361_module_data_in[4] ;
 wire \sw_361_module_data_in[5] ;
 wire \sw_361_module_data_in[6] ;
 wire \sw_361_module_data_in[7] ;
 wire \sw_361_module_data_out[0] ;
 wire \sw_361_module_data_out[1] ;
 wire \sw_361_module_data_out[2] ;
 wire \sw_361_module_data_out[3] ;
 wire \sw_361_module_data_out[4] ;
 wire \sw_361_module_data_out[5] ;
 wire \sw_361_module_data_out[6] ;
 wire \sw_361_module_data_out[7] ;
 wire sw_361_scan_out;
 wire sw_362_clk_out;
 wire sw_362_data_out;
 wire sw_362_latch_out;
 wire \sw_362_module_data_in[0] ;
 wire \sw_362_module_data_in[1] ;
 wire \sw_362_module_data_in[2] ;
 wire \sw_362_module_data_in[3] ;
 wire \sw_362_module_data_in[4] ;
 wire \sw_362_module_data_in[5] ;
 wire \sw_362_module_data_in[6] ;
 wire \sw_362_module_data_in[7] ;
 wire \sw_362_module_data_out[0] ;
 wire \sw_362_module_data_out[1] ;
 wire \sw_362_module_data_out[2] ;
 wire \sw_362_module_data_out[3] ;
 wire \sw_362_module_data_out[4] ;
 wire \sw_362_module_data_out[5] ;
 wire \sw_362_module_data_out[6] ;
 wire \sw_362_module_data_out[7] ;
 wire sw_362_scan_out;
 wire sw_363_clk_out;
 wire sw_363_data_out;
 wire sw_363_latch_out;
 wire \sw_363_module_data_in[0] ;
 wire \sw_363_module_data_in[1] ;
 wire \sw_363_module_data_in[2] ;
 wire \sw_363_module_data_in[3] ;
 wire \sw_363_module_data_in[4] ;
 wire \sw_363_module_data_in[5] ;
 wire \sw_363_module_data_in[6] ;
 wire \sw_363_module_data_in[7] ;
 wire \sw_363_module_data_out[0] ;
 wire \sw_363_module_data_out[1] ;
 wire \sw_363_module_data_out[2] ;
 wire \sw_363_module_data_out[3] ;
 wire \sw_363_module_data_out[4] ;
 wire \sw_363_module_data_out[5] ;
 wire \sw_363_module_data_out[6] ;
 wire \sw_363_module_data_out[7] ;
 wire sw_363_scan_out;
 wire sw_364_clk_out;
 wire sw_364_data_out;
 wire sw_364_latch_out;
 wire \sw_364_module_data_in[0] ;
 wire \sw_364_module_data_in[1] ;
 wire \sw_364_module_data_in[2] ;
 wire \sw_364_module_data_in[3] ;
 wire \sw_364_module_data_in[4] ;
 wire \sw_364_module_data_in[5] ;
 wire \sw_364_module_data_in[6] ;
 wire \sw_364_module_data_in[7] ;
 wire \sw_364_module_data_out[0] ;
 wire \sw_364_module_data_out[1] ;
 wire \sw_364_module_data_out[2] ;
 wire \sw_364_module_data_out[3] ;
 wire \sw_364_module_data_out[4] ;
 wire \sw_364_module_data_out[5] ;
 wire \sw_364_module_data_out[6] ;
 wire \sw_364_module_data_out[7] ;
 wire sw_364_scan_out;
 wire sw_365_clk_out;
 wire sw_365_data_out;
 wire sw_365_latch_out;
 wire \sw_365_module_data_in[0] ;
 wire \sw_365_module_data_in[1] ;
 wire \sw_365_module_data_in[2] ;
 wire \sw_365_module_data_in[3] ;
 wire \sw_365_module_data_in[4] ;
 wire \sw_365_module_data_in[5] ;
 wire \sw_365_module_data_in[6] ;
 wire \sw_365_module_data_in[7] ;
 wire \sw_365_module_data_out[0] ;
 wire \sw_365_module_data_out[1] ;
 wire \sw_365_module_data_out[2] ;
 wire \sw_365_module_data_out[3] ;
 wire \sw_365_module_data_out[4] ;
 wire \sw_365_module_data_out[5] ;
 wire \sw_365_module_data_out[6] ;
 wire \sw_365_module_data_out[7] ;
 wire sw_365_scan_out;
 wire sw_366_clk_out;
 wire sw_366_data_out;
 wire sw_366_latch_out;
 wire \sw_366_module_data_in[0] ;
 wire \sw_366_module_data_in[1] ;
 wire \sw_366_module_data_in[2] ;
 wire \sw_366_module_data_in[3] ;
 wire \sw_366_module_data_in[4] ;
 wire \sw_366_module_data_in[5] ;
 wire \sw_366_module_data_in[6] ;
 wire \sw_366_module_data_in[7] ;
 wire \sw_366_module_data_out[0] ;
 wire \sw_366_module_data_out[1] ;
 wire \sw_366_module_data_out[2] ;
 wire \sw_366_module_data_out[3] ;
 wire \sw_366_module_data_out[4] ;
 wire \sw_366_module_data_out[5] ;
 wire \sw_366_module_data_out[6] ;
 wire \sw_366_module_data_out[7] ;
 wire sw_366_scan_out;
 wire sw_367_clk_out;
 wire sw_367_data_out;
 wire sw_367_latch_out;
 wire \sw_367_module_data_in[0] ;
 wire \sw_367_module_data_in[1] ;
 wire \sw_367_module_data_in[2] ;
 wire \sw_367_module_data_in[3] ;
 wire \sw_367_module_data_in[4] ;
 wire \sw_367_module_data_in[5] ;
 wire \sw_367_module_data_in[6] ;
 wire \sw_367_module_data_in[7] ;
 wire \sw_367_module_data_out[0] ;
 wire \sw_367_module_data_out[1] ;
 wire \sw_367_module_data_out[2] ;
 wire \sw_367_module_data_out[3] ;
 wire \sw_367_module_data_out[4] ;
 wire \sw_367_module_data_out[5] ;
 wire \sw_367_module_data_out[6] ;
 wire \sw_367_module_data_out[7] ;
 wire sw_367_scan_out;
 wire sw_368_clk_out;
 wire sw_368_data_out;
 wire sw_368_latch_out;
 wire \sw_368_module_data_in[0] ;
 wire \sw_368_module_data_in[1] ;
 wire \sw_368_module_data_in[2] ;
 wire \sw_368_module_data_in[3] ;
 wire \sw_368_module_data_in[4] ;
 wire \sw_368_module_data_in[5] ;
 wire \sw_368_module_data_in[6] ;
 wire \sw_368_module_data_in[7] ;
 wire \sw_368_module_data_out[0] ;
 wire \sw_368_module_data_out[1] ;
 wire \sw_368_module_data_out[2] ;
 wire \sw_368_module_data_out[3] ;
 wire \sw_368_module_data_out[4] ;
 wire \sw_368_module_data_out[5] ;
 wire \sw_368_module_data_out[6] ;
 wire \sw_368_module_data_out[7] ;
 wire sw_368_scan_out;
 wire sw_369_clk_out;
 wire sw_369_data_out;
 wire sw_369_latch_out;
 wire \sw_369_module_data_in[0] ;
 wire \sw_369_module_data_in[1] ;
 wire \sw_369_module_data_in[2] ;
 wire \sw_369_module_data_in[3] ;
 wire \sw_369_module_data_in[4] ;
 wire \sw_369_module_data_in[5] ;
 wire \sw_369_module_data_in[6] ;
 wire \sw_369_module_data_in[7] ;
 wire \sw_369_module_data_out[0] ;
 wire \sw_369_module_data_out[1] ;
 wire \sw_369_module_data_out[2] ;
 wire \sw_369_module_data_out[3] ;
 wire \sw_369_module_data_out[4] ;
 wire \sw_369_module_data_out[5] ;
 wire \sw_369_module_data_out[6] ;
 wire \sw_369_module_data_out[7] ;
 wire sw_369_scan_out;
 wire sw_370_clk_out;
 wire sw_370_data_out;
 wire sw_370_latch_out;
 wire \sw_370_module_data_in[0] ;
 wire \sw_370_module_data_in[1] ;
 wire \sw_370_module_data_in[2] ;
 wire \sw_370_module_data_in[3] ;
 wire \sw_370_module_data_in[4] ;
 wire \sw_370_module_data_in[5] ;
 wire \sw_370_module_data_in[6] ;
 wire \sw_370_module_data_in[7] ;
 wire \sw_370_module_data_out[0] ;
 wire \sw_370_module_data_out[1] ;
 wire \sw_370_module_data_out[2] ;
 wire \sw_370_module_data_out[3] ;
 wire \sw_370_module_data_out[4] ;
 wire \sw_370_module_data_out[5] ;
 wire \sw_370_module_data_out[6] ;
 wire \sw_370_module_data_out[7] ;
 wire sw_370_scan_out;
 wire sw_371_clk_out;
 wire sw_371_data_out;
 wire sw_371_latch_out;
 wire \sw_371_module_data_in[0] ;
 wire \sw_371_module_data_in[1] ;
 wire \sw_371_module_data_in[2] ;
 wire \sw_371_module_data_in[3] ;
 wire \sw_371_module_data_in[4] ;
 wire \sw_371_module_data_in[5] ;
 wire \sw_371_module_data_in[6] ;
 wire \sw_371_module_data_in[7] ;
 wire \sw_371_module_data_out[0] ;
 wire \sw_371_module_data_out[1] ;
 wire \sw_371_module_data_out[2] ;
 wire \sw_371_module_data_out[3] ;
 wire \sw_371_module_data_out[4] ;
 wire \sw_371_module_data_out[5] ;
 wire \sw_371_module_data_out[6] ;
 wire \sw_371_module_data_out[7] ;
 wire sw_371_scan_out;
 wire sw_372_clk_out;
 wire sw_372_data_out;
 wire sw_372_latch_out;
 wire \sw_372_module_data_in[0] ;
 wire \sw_372_module_data_in[1] ;
 wire \sw_372_module_data_in[2] ;
 wire \sw_372_module_data_in[3] ;
 wire \sw_372_module_data_in[4] ;
 wire \sw_372_module_data_in[5] ;
 wire \sw_372_module_data_in[6] ;
 wire \sw_372_module_data_in[7] ;
 wire \sw_372_module_data_out[0] ;
 wire \sw_372_module_data_out[1] ;
 wire \sw_372_module_data_out[2] ;
 wire \sw_372_module_data_out[3] ;
 wire \sw_372_module_data_out[4] ;
 wire \sw_372_module_data_out[5] ;
 wire \sw_372_module_data_out[6] ;
 wire \sw_372_module_data_out[7] ;
 wire sw_372_scan_out;
 wire sw_373_clk_out;
 wire sw_373_data_out;
 wire sw_373_latch_out;
 wire \sw_373_module_data_in[0] ;
 wire \sw_373_module_data_in[1] ;
 wire \sw_373_module_data_in[2] ;
 wire \sw_373_module_data_in[3] ;
 wire \sw_373_module_data_in[4] ;
 wire \sw_373_module_data_in[5] ;
 wire \sw_373_module_data_in[6] ;
 wire \sw_373_module_data_in[7] ;
 wire \sw_373_module_data_out[0] ;
 wire \sw_373_module_data_out[1] ;
 wire \sw_373_module_data_out[2] ;
 wire \sw_373_module_data_out[3] ;
 wire \sw_373_module_data_out[4] ;
 wire \sw_373_module_data_out[5] ;
 wire \sw_373_module_data_out[6] ;
 wire \sw_373_module_data_out[7] ;
 wire sw_373_scan_out;
 wire sw_374_clk_out;
 wire sw_374_data_out;
 wire sw_374_latch_out;
 wire \sw_374_module_data_in[0] ;
 wire \sw_374_module_data_in[1] ;
 wire \sw_374_module_data_in[2] ;
 wire \sw_374_module_data_in[3] ;
 wire \sw_374_module_data_in[4] ;
 wire \sw_374_module_data_in[5] ;
 wire \sw_374_module_data_in[6] ;
 wire \sw_374_module_data_in[7] ;
 wire \sw_374_module_data_out[0] ;
 wire \sw_374_module_data_out[1] ;
 wire \sw_374_module_data_out[2] ;
 wire \sw_374_module_data_out[3] ;
 wire \sw_374_module_data_out[4] ;
 wire \sw_374_module_data_out[5] ;
 wire \sw_374_module_data_out[6] ;
 wire \sw_374_module_data_out[7] ;
 wire sw_374_scan_out;
 wire sw_375_clk_out;
 wire sw_375_data_out;
 wire sw_375_latch_out;
 wire \sw_375_module_data_in[0] ;
 wire \sw_375_module_data_in[1] ;
 wire \sw_375_module_data_in[2] ;
 wire \sw_375_module_data_in[3] ;
 wire \sw_375_module_data_in[4] ;
 wire \sw_375_module_data_in[5] ;
 wire \sw_375_module_data_in[6] ;
 wire \sw_375_module_data_in[7] ;
 wire \sw_375_module_data_out[0] ;
 wire \sw_375_module_data_out[1] ;
 wire \sw_375_module_data_out[2] ;
 wire \sw_375_module_data_out[3] ;
 wire \sw_375_module_data_out[4] ;
 wire \sw_375_module_data_out[5] ;
 wire \sw_375_module_data_out[6] ;
 wire \sw_375_module_data_out[7] ;
 wire sw_375_scan_out;
 wire sw_376_clk_out;
 wire sw_376_data_out;
 wire sw_376_latch_out;
 wire \sw_376_module_data_in[0] ;
 wire \sw_376_module_data_in[1] ;
 wire \sw_376_module_data_in[2] ;
 wire \sw_376_module_data_in[3] ;
 wire \sw_376_module_data_in[4] ;
 wire \sw_376_module_data_in[5] ;
 wire \sw_376_module_data_in[6] ;
 wire \sw_376_module_data_in[7] ;
 wire \sw_376_module_data_out[0] ;
 wire \sw_376_module_data_out[1] ;
 wire \sw_376_module_data_out[2] ;
 wire \sw_376_module_data_out[3] ;
 wire \sw_376_module_data_out[4] ;
 wire \sw_376_module_data_out[5] ;
 wire \sw_376_module_data_out[6] ;
 wire \sw_376_module_data_out[7] ;
 wire sw_376_scan_out;
 wire sw_377_clk_out;
 wire sw_377_data_out;
 wire sw_377_latch_out;
 wire \sw_377_module_data_in[0] ;
 wire \sw_377_module_data_in[1] ;
 wire \sw_377_module_data_in[2] ;
 wire \sw_377_module_data_in[3] ;
 wire \sw_377_module_data_in[4] ;
 wire \sw_377_module_data_in[5] ;
 wire \sw_377_module_data_in[6] ;
 wire \sw_377_module_data_in[7] ;
 wire \sw_377_module_data_out[0] ;
 wire \sw_377_module_data_out[1] ;
 wire \sw_377_module_data_out[2] ;
 wire \sw_377_module_data_out[3] ;
 wire \sw_377_module_data_out[4] ;
 wire \sw_377_module_data_out[5] ;
 wire \sw_377_module_data_out[6] ;
 wire \sw_377_module_data_out[7] ;
 wire sw_377_scan_out;
 wire sw_378_clk_out;
 wire sw_378_data_out;
 wire sw_378_latch_out;
 wire \sw_378_module_data_in[0] ;
 wire \sw_378_module_data_in[1] ;
 wire \sw_378_module_data_in[2] ;
 wire \sw_378_module_data_in[3] ;
 wire \sw_378_module_data_in[4] ;
 wire \sw_378_module_data_in[5] ;
 wire \sw_378_module_data_in[6] ;
 wire \sw_378_module_data_in[7] ;
 wire \sw_378_module_data_out[0] ;
 wire \sw_378_module_data_out[1] ;
 wire \sw_378_module_data_out[2] ;
 wire \sw_378_module_data_out[3] ;
 wire \sw_378_module_data_out[4] ;
 wire \sw_378_module_data_out[5] ;
 wire \sw_378_module_data_out[6] ;
 wire \sw_378_module_data_out[7] ;
 wire sw_378_scan_out;
 wire sw_379_clk_out;
 wire sw_379_data_out;
 wire sw_379_latch_out;
 wire \sw_379_module_data_in[0] ;
 wire \sw_379_module_data_in[1] ;
 wire \sw_379_module_data_in[2] ;
 wire \sw_379_module_data_in[3] ;
 wire \sw_379_module_data_in[4] ;
 wire \sw_379_module_data_in[5] ;
 wire \sw_379_module_data_in[6] ;
 wire \sw_379_module_data_in[7] ;
 wire \sw_379_module_data_out[0] ;
 wire \sw_379_module_data_out[1] ;
 wire \sw_379_module_data_out[2] ;
 wire \sw_379_module_data_out[3] ;
 wire \sw_379_module_data_out[4] ;
 wire \sw_379_module_data_out[5] ;
 wire \sw_379_module_data_out[6] ;
 wire \sw_379_module_data_out[7] ;
 wire sw_379_scan_out;
 wire sw_380_clk_out;
 wire sw_380_data_out;
 wire sw_380_latch_out;
 wire \sw_380_module_data_in[0] ;
 wire \sw_380_module_data_in[1] ;
 wire \sw_380_module_data_in[2] ;
 wire \sw_380_module_data_in[3] ;
 wire \sw_380_module_data_in[4] ;
 wire \sw_380_module_data_in[5] ;
 wire \sw_380_module_data_in[6] ;
 wire \sw_380_module_data_in[7] ;
 wire \sw_380_module_data_out[0] ;
 wire \sw_380_module_data_out[1] ;
 wire \sw_380_module_data_out[2] ;
 wire \sw_380_module_data_out[3] ;
 wire \sw_380_module_data_out[4] ;
 wire \sw_380_module_data_out[5] ;
 wire \sw_380_module_data_out[6] ;
 wire \sw_380_module_data_out[7] ;
 wire sw_380_scan_out;
 wire sw_381_clk_out;
 wire sw_381_data_out;
 wire sw_381_latch_out;
 wire \sw_381_module_data_in[0] ;
 wire \sw_381_module_data_in[1] ;
 wire \sw_381_module_data_in[2] ;
 wire \sw_381_module_data_in[3] ;
 wire \sw_381_module_data_in[4] ;
 wire \sw_381_module_data_in[5] ;
 wire \sw_381_module_data_in[6] ;
 wire \sw_381_module_data_in[7] ;
 wire \sw_381_module_data_out[0] ;
 wire \sw_381_module_data_out[1] ;
 wire \sw_381_module_data_out[2] ;
 wire \sw_381_module_data_out[3] ;
 wire \sw_381_module_data_out[4] ;
 wire \sw_381_module_data_out[5] ;
 wire \sw_381_module_data_out[6] ;
 wire \sw_381_module_data_out[7] ;
 wire sw_381_scan_out;
 wire sw_382_clk_out;
 wire sw_382_data_out;
 wire sw_382_latch_out;
 wire \sw_382_module_data_in[0] ;
 wire \sw_382_module_data_in[1] ;
 wire \sw_382_module_data_in[2] ;
 wire \sw_382_module_data_in[3] ;
 wire \sw_382_module_data_in[4] ;
 wire \sw_382_module_data_in[5] ;
 wire \sw_382_module_data_in[6] ;
 wire \sw_382_module_data_in[7] ;
 wire \sw_382_module_data_out[0] ;
 wire \sw_382_module_data_out[1] ;
 wire \sw_382_module_data_out[2] ;
 wire \sw_382_module_data_out[3] ;
 wire \sw_382_module_data_out[4] ;
 wire \sw_382_module_data_out[5] ;
 wire \sw_382_module_data_out[6] ;
 wire \sw_382_module_data_out[7] ;
 wire sw_382_scan_out;
 wire sw_383_clk_out;
 wire sw_383_data_out;
 wire sw_383_latch_out;
 wire \sw_383_module_data_in[0] ;
 wire \sw_383_module_data_in[1] ;
 wire \sw_383_module_data_in[2] ;
 wire \sw_383_module_data_in[3] ;
 wire \sw_383_module_data_in[4] ;
 wire \sw_383_module_data_in[5] ;
 wire \sw_383_module_data_in[6] ;
 wire \sw_383_module_data_in[7] ;
 wire \sw_383_module_data_out[0] ;
 wire \sw_383_module_data_out[1] ;
 wire \sw_383_module_data_out[2] ;
 wire \sw_383_module_data_out[3] ;
 wire \sw_383_module_data_out[4] ;
 wire \sw_383_module_data_out[5] ;
 wire \sw_383_module_data_out[6] ;
 wire \sw_383_module_data_out[7] ;
 wire sw_383_scan_out;
 wire sw_384_clk_out;
 wire sw_384_data_out;
 wire sw_384_latch_out;
 wire \sw_384_module_data_in[0] ;
 wire \sw_384_module_data_in[1] ;
 wire \sw_384_module_data_in[2] ;
 wire \sw_384_module_data_in[3] ;
 wire \sw_384_module_data_in[4] ;
 wire \sw_384_module_data_in[5] ;
 wire \sw_384_module_data_in[6] ;
 wire \sw_384_module_data_in[7] ;
 wire \sw_384_module_data_out[0] ;
 wire \sw_384_module_data_out[1] ;
 wire \sw_384_module_data_out[2] ;
 wire \sw_384_module_data_out[3] ;
 wire \sw_384_module_data_out[4] ;
 wire \sw_384_module_data_out[5] ;
 wire \sw_384_module_data_out[6] ;
 wire \sw_384_module_data_out[7] ;
 wire sw_384_scan_out;
 wire sw_385_clk_out;
 wire sw_385_data_out;
 wire sw_385_latch_out;
 wire \sw_385_module_data_in[0] ;
 wire \sw_385_module_data_in[1] ;
 wire \sw_385_module_data_in[2] ;
 wire \sw_385_module_data_in[3] ;
 wire \sw_385_module_data_in[4] ;
 wire \sw_385_module_data_in[5] ;
 wire \sw_385_module_data_in[6] ;
 wire \sw_385_module_data_in[7] ;
 wire \sw_385_module_data_out[0] ;
 wire \sw_385_module_data_out[1] ;
 wire \sw_385_module_data_out[2] ;
 wire \sw_385_module_data_out[3] ;
 wire \sw_385_module_data_out[4] ;
 wire \sw_385_module_data_out[5] ;
 wire \sw_385_module_data_out[6] ;
 wire \sw_385_module_data_out[7] ;
 wire sw_385_scan_out;
 wire sw_386_clk_out;
 wire sw_386_data_out;
 wire sw_386_latch_out;
 wire \sw_386_module_data_in[0] ;
 wire \sw_386_module_data_in[1] ;
 wire \sw_386_module_data_in[2] ;
 wire \sw_386_module_data_in[3] ;
 wire \sw_386_module_data_in[4] ;
 wire \sw_386_module_data_in[5] ;
 wire \sw_386_module_data_in[6] ;
 wire \sw_386_module_data_in[7] ;
 wire \sw_386_module_data_out[0] ;
 wire \sw_386_module_data_out[1] ;
 wire \sw_386_module_data_out[2] ;
 wire \sw_386_module_data_out[3] ;
 wire \sw_386_module_data_out[4] ;
 wire \sw_386_module_data_out[5] ;
 wire \sw_386_module_data_out[6] ;
 wire \sw_386_module_data_out[7] ;
 wire sw_386_scan_out;
 wire sw_387_clk_out;
 wire sw_387_data_out;
 wire sw_387_latch_out;
 wire \sw_387_module_data_in[0] ;
 wire \sw_387_module_data_in[1] ;
 wire \sw_387_module_data_in[2] ;
 wire \sw_387_module_data_in[3] ;
 wire \sw_387_module_data_in[4] ;
 wire \sw_387_module_data_in[5] ;
 wire \sw_387_module_data_in[6] ;
 wire \sw_387_module_data_in[7] ;
 wire \sw_387_module_data_out[0] ;
 wire \sw_387_module_data_out[1] ;
 wire \sw_387_module_data_out[2] ;
 wire \sw_387_module_data_out[3] ;
 wire \sw_387_module_data_out[4] ;
 wire \sw_387_module_data_out[5] ;
 wire \sw_387_module_data_out[6] ;
 wire \sw_387_module_data_out[7] ;
 wire sw_387_scan_out;
 wire sw_388_clk_out;
 wire sw_388_data_out;
 wire sw_388_latch_out;
 wire \sw_388_module_data_in[0] ;
 wire \sw_388_module_data_in[1] ;
 wire \sw_388_module_data_in[2] ;
 wire \sw_388_module_data_in[3] ;
 wire \sw_388_module_data_in[4] ;
 wire \sw_388_module_data_in[5] ;
 wire \sw_388_module_data_in[6] ;
 wire \sw_388_module_data_in[7] ;
 wire \sw_388_module_data_out[0] ;
 wire \sw_388_module_data_out[1] ;
 wire \sw_388_module_data_out[2] ;
 wire \sw_388_module_data_out[3] ;
 wire \sw_388_module_data_out[4] ;
 wire \sw_388_module_data_out[5] ;
 wire \sw_388_module_data_out[6] ;
 wire \sw_388_module_data_out[7] ;
 wire sw_388_scan_out;
 wire sw_389_clk_out;
 wire sw_389_data_out;
 wire sw_389_latch_out;
 wire \sw_389_module_data_in[0] ;
 wire \sw_389_module_data_in[1] ;
 wire \sw_389_module_data_in[2] ;
 wire \sw_389_module_data_in[3] ;
 wire \sw_389_module_data_in[4] ;
 wire \sw_389_module_data_in[5] ;
 wire \sw_389_module_data_in[6] ;
 wire \sw_389_module_data_in[7] ;
 wire \sw_389_module_data_out[0] ;
 wire \sw_389_module_data_out[1] ;
 wire \sw_389_module_data_out[2] ;
 wire \sw_389_module_data_out[3] ;
 wire \sw_389_module_data_out[4] ;
 wire \sw_389_module_data_out[5] ;
 wire \sw_389_module_data_out[6] ;
 wire \sw_389_module_data_out[7] ;
 wire sw_389_scan_out;
 wire sw_390_clk_out;
 wire sw_390_data_out;
 wire sw_390_latch_out;
 wire \sw_390_module_data_in[0] ;
 wire \sw_390_module_data_in[1] ;
 wire \sw_390_module_data_in[2] ;
 wire \sw_390_module_data_in[3] ;
 wire \sw_390_module_data_in[4] ;
 wire \sw_390_module_data_in[5] ;
 wire \sw_390_module_data_in[6] ;
 wire \sw_390_module_data_in[7] ;
 wire \sw_390_module_data_out[0] ;
 wire \sw_390_module_data_out[1] ;
 wire \sw_390_module_data_out[2] ;
 wire \sw_390_module_data_out[3] ;
 wire \sw_390_module_data_out[4] ;
 wire \sw_390_module_data_out[5] ;
 wire \sw_390_module_data_out[6] ;
 wire \sw_390_module_data_out[7] ;
 wire sw_390_scan_out;
 wire sw_391_clk_out;
 wire sw_391_data_out;
 wire sw_391_latch_out;
 wire \sw_391_module_data_in[0] ;
 wire \sw_391_module_data_in[1] ;
 wire \sw_391_module_data_in[2] ;
 wire \sw_391_module_data_in[3] ;
 wire \sw_391_module_data_in[4] ;
 wire \sw_391_module_data_in[5] ;
 wire \sw_391_module_data_in[6] ;
 wire \sw_391_module_data_in[7] ;
 wire \sw_391_module_data_out[0] ;
 wire \sw_391_module_data_out[1] ;
 wire \sw_391_module_data_out[2] ;
 wire \sw_391_module_data_out[3] ;
 wire \sw_391_module_data_out[4] ;
 wire \sw_391_module_data_out[5] ;
 wire \sw_391_module_data_out[6] ;
 wire \sw_391_module_data_out[7] ;
 wire sw_391_scan_out;
 wire sw_392_clk_out;
 wire sw_392_data_out;
 wire sw_392_latch_out;
 wire \sw_392_module_data_in[0] ;
 wire \sw_392_module_data_in[1] ;
 wire \sw_392_module_data_in[2] ;
 wire \sw_392_module_data_in[3] ;
 wire \sw_392_module_data_in[4] ;
 wire \sw_392_module_data_in[5] ;
 wire \sw_392_module_data_in[6] ;
 wire \sw_392_module_data_in[7] ;
 wire \sw_392_module_data_out[0] ;
 wire \sw_392_module_data_out[1] ;
 wire \sw_392_module_data_out[2] ;
 wire \sw_392_module_data_out[3] ;
 wire \sw_392_module_data_out[4] ;
 wire \sw_392_module_data_out[5] ;
 wire \sw_392_module_data_out[6] ;
 wire \sw_392_module_data_out[7] ;
 wire sw_392_scan_out;
 wire sw_393_clk_out;
 wire sw_393_data_out;
 wire sw_393_latch_out;
 wire \sw_393_module_data_in[0] ;
 wire \sw_393_module_data_in[1] ;
 wire \sw_393_module_data_in[2] ;
 wire \sw_393_module_data_in[3] ;
 wire \sw_393_module_data_in[4] ;
 wire \sw_393_module_data_in[5] ;
 wire \sw_393_module_data_in[6] ;
 wire \sw_393_module_data_in[7] ;
 wire \sw_393_module_data_out[0] ;
 wire \sw_393_module_data_out[1] ;
 wire \sw_393_module_data_out[2] ;
 wire \sw_393_module_data_out[3] ;
 wire \sw_393_module_data_out[4] ;
 wire \sw_393_module_data_out[5] ;
 wire \sw_393_module_data_out[6] ;
 wire \sw_393_module_data_out[7] ;
 wire sw_393_scan_out;
 wire sw_394_clk_out;
 wire sw_394_data_out;
 wire sw_394_latch_out;
 wire \sw_394_module_data_in[0] ;
 wire \sw_394_module_data_in[1] ;
 wire \sw_394_module_data_in[2] ;
 wire \sw_394_module_data_in[3] ;
 wire \sw_394_module_data_in[4] ;
 wire \sw_394_module_data_in[5] ;
 wire \sw_394_module_data_in[6] ;
 wire \sw_394_module_data_in[7] ;
 wire \sw_394_module_data_out[0] ;
 wire \sw_394_module_data_out[1] ;
 wire \sw_394_module_data_out[2] ;
 wire \sw_394_module_data_out[3] ;
 wire \sw_394_module_data_out[4] ;
 wire \sw_394_module_data_out[5] ;
 wire \sw_394_module_data_out[6] ;
 wire \sw_394_module_data_out[7] ;
 wire sw_394_scan_out;
 wire sw_395_clk_out;
 wire sw_395_data_out;
 wire sw_395_latch_out;
 wire \sw_395_module_data_in[0] ;
 wire \sw_395_module_data_in[1] ;
 wire \sw_395_module_data_in[2] ;
 wire \sw_395_module_data_in[3] ;
 wire \sw_395_module_data_in[4] ;
 wire \sw_395_module_data_in[5] ;
 wire \sw_395_module_data_in[6] ;
 wire \sw_395_module_data_in[7] ;
 wire \sw_395_module_data_out[0] ;
 wire \sw_395_module_data_out[1] ;
 wire \sw_395_module_data_out[2] ;
 wire \sw_395_module_data_out[3] ;
 wire \sw_395_module_data_out[4] ;
 wire \sw_395_module_data_out[5] ;
 wire \sw_395_module_data_out[6] ;
 wire \sw_395_module_data_out[7] ;
 wire sw_395_scan_out;
 wire sw_396_clk_out;
 wire sw_396_data_out;
 wire sw_396_latch_out;
 wire \sw_396_module_data_in[0] ;
 wire \sw_396_module_data_in[1] ;
 wire \sw_396_module_data_in[2] ;
 wire \sw_396_module_data_in[3] ;
 wire \sw_396_module_data_in[4] ;
 wire \sw_396_module_data_in[5] ;
 wire \sw_396_module_data_in[6] ;
 wire \sw_396_module_data_in[7] ;
 wire \sw_396_module_data_out[0] ;
 wire \sw_396_module_data_out[1] ;
 wire \sw_396_module_data_out[2] ;
 wire \sw_396_module_data_out[3] ;
 wire \sw_396_module_data_out[4] ;
 wire \sw_396_module_data_out[5] ;
 wire \sw_396_module_data_out[6] ;
 wire \sw_396_module_data_out[7] ;
 wire sw_396_scan_out;
 wire sw_397_clk_out;
 wire sw_397_data_out;
 wire sw_397_latch_out;
 wire \sw_397_module_data_in[0] ;
 wire \sw_397_module_data_in[1] ;
 wire \sw_397_module_data_in[2] ;
 wire \sw_397_module_data_in[3] ;
 wire \sw_397_module_data_in[4] ;
 wire \sw_397_module_data_in[5] ;
 wire \sw_397_module_data_in[6] ;
 wire \sw_397_module_data_in[7] ;
 wire \sw_397_module_data_out[0] ;
 wire \sw_397_module_data_out[1] ;
 wire \sw_397_module_data_out[2] ;
 wire \sw_397_module_data_out[3] ;
 wire \sw_397_module_data_out[4] ;
 wire \sw_397_module_data_out[5] ;
 wire \sw_397_module_data_out[6] ;
 wire \sw_397_module_data_out[7] ;
 wire sw_397_scan_out;
 wire sw_398_clk_out;
 wire sw_398_data_out;
 wire sw_398_latch_out;
 wire \sw_398_module_data_in[0] ;
 wire \sw_398_module_data_in[1] ;
 wire \sw_398_module_data_in[2] ;
 wire \sw_398_module_data_in[3] ;
 wire \sw_398_module_data_in[4] ;
 wire \sw_398_module_data_in[5] ;
 wire \sw_398_module_data_in[6] ;
 wire \sw_398_module_data_in[7] ;
 wire \sw_398_module_data_out[0] ;
 wire \sw_398_module_data_out[1] ;
 wire \sw_398_module_data_out[2] ;
 wire \sw_398_module_data_out[3] ;
 wire \sw_398_module_data_out[4] ;
 wire \sw_398_module_data_out[5] ;
 wire \sw_398_module_data_out[6] ;
 wire \sw_398_module_data_out[7] ;
 wire sw_398_scan_out;
 wire sw_399_clk_out;
 wire sw_399_data_out;
 wire sw_399_latch_out;
 wire \sw_399_module_data_in[0] ;
 wire \sw_399_module_data_in[1] ;
 wire \sw_399_module_data_in[2] ;
 wire \sw_399_module_data_in[3] ;
 wire \sw_399_module_data_in[4] ;
 wire \sw_399_module_data_in[5] ;
 wire \sw_399_module_data_in[6] ;
 wire \sw_399_module_data_in[7] ;
 wire \sw_399_module_data_out[0] ;
 wire \sw_399_module_data_out[1] ;
 wire \sw_399_module_data_out[2] ;
 wire \sw_399_module_data_out[3] ;
 wire \sw_399_module_data_out[4] ;
 wire \sw_399_module_data_out[5] ;
 wire \sw_399_module_data_out[6] ;
 wire \sw_399_module_data_out[7] ;
 wire sw_399_scan_out;
 wire sw_400_clk_out;
 wire sw_400_data_out;
 wire sw_400_latch_out;
 wire \sw_400_module_data_in[0] ;
 wire \sw_400_module_data_in[1] ;
 wire \sw_400_module_data_in[2] ;
 wire \sw_400_module_data_in[3] ;
 wire \sw_400_module_data_in[4] ;
 wire \sw_400_module_data_in[5] ;
 wire \sw_400_module_data_in[6] ;
 wire \sw_400_module_data_in[7] ;
 wire \sw_400_module_data_out[0] ;
 wire \sw_400_module_data_out[1] ;
 wire \sw_400_module_data_out[2] ;
 wire \sw_400_module_data_out[3] ;
 wire \sw_400_module_data_out[4] ;
 wire \sw_400_module_data_out[5] ;
 wire \sw_400_module_data_out[6] ;
 wire \sw_400_module_data_out[7] ;
 wire sw_400_scan_out;
 wire sw_401_clk_out;
 wire sw_401_data_out;
 wire sw_401_latch_out;
 wire \sw_401_module_data_in[0] ;
 wire \sw_401_module_data_in[1] ;
 wire \sw_401_module_data_in[2] ;
 wire \sw_401_module_data_in[3] ;
 wire \sw_401_module_data_in[4] ;
 wire \sw_401_module_data_in[5] ;
 wire \sw_401_module_data_in[6] ;
 wire \sw_401_module_data_in[7] ;
 wire \sw_401_module_data_out[0] ;
 wire \sw_401_module_data_out[1] ;
 wire \sw_401_module_data_out[2] ;
 wire \sw_401_module_data_out[3] ;
 wire \sw_401_module_data_out[4] ;
 wire \sw_401_module_data_out[5] ;
 wire \sw_401_module_data_out[6] ;
 wire \sw_401_module_data_out[7] ;
 wire sw_401_scan_out;
 wire sw_402_clk_out;
 wire sw_402_data_out;
 wire sw_402_latch_out;
 wire \sw_402_module_data_in[0] ;
 wire \sw_402_module_data_in[1] ;
 wire \sw_402_module_data_in[2] ;
 wire \sw_402_module_data_in[3] ;
 wire \sw_402_module_data_in[4] ;
 wire \sw_402_module_data_in[5] ;
 wire \sw_402_module_data_in[6] ;
 wire \sw_402_module_data_in[7] ;
 wire \sw_402_module_data_out[0] ;
 wire \sw_402_module_data_out[1] ;
 wire \sw_402_module_data_out[2] ;
 wire \sw_402_module_data_out[3] ;
 wire \sw_402_module_data_out[4] ;
 wire \sw_402_module_data_out[5] ;
 wire \sw_402_module_data_out[6] ;
 wire \sw_402_module_data_out[7] ;
 wire sw_402_scan_out;
 wire sw_403_clk_out;
 wire sw_403_data_out;
 wire sw_403_latch_out;
 wire \sw_403_module_data_in[0] ;
 wire \sw_403_module_data_in[1] ;
 wire \sw_403_module_data_in[2] ;
 wire \sw_403_module_data_in[3] ;
 wire \sw_403_module_data_in[4] ;
 wire \sw_403_module_data_in[5] ;
 wire \sw_403_module_data_in[6] ;
 wire \sw_403_module_data_in[7] ;
 wire \sw_403_module_data_out[0] ;
 wire \sw_403_module_data_out[1] ;
 wire \sw_403_module_data_out[2] ;
 wire \sw_403_module_data_out[3] ;
 wire \sw_403_module_data_out[4] ;
 wire \sw_403_module_data_out[5] ;
 wire \sw_403_module_data_out[6] ;
 wire \sw_403_module_data_out[7] ;
 wire sw_403_scan_out;
 wire sw_404_clk_out;
 wire sw_404_data_out;
 wire sw_404_latch_out;
 wire \sw_404_module_data_in[0] ;
 wire \sw_404_module_data_in[1] ;
 wire \sw_404_module_data_in[2] ;
 wire \sw_404_module_data_in[3] ;
 wire \sw_404_module_data_in[4] ;
 wire \sw_404_module_data_in[5] ;
 wire \sw_404_module_data_in[6] ;
 wire \sw_404_module_data_in[7] ;
 wire \sw_404_module_data_out[0] ;
 wire \sw_404_module_data_out[1] ;
 wire \sw_404_module_data_out[2] ;
 wire \sw_404_module_data_out[3] ;
 wire \sw_404_module_data_out[4] ;
 wire \sw_404_module_data_out[5] ;
 wire \sw_404_module_data_out[6] ;
 wire \sw_404_module_data_out[7] ;
 wire sw_404_scan_out;
 wire sw_405_clk_out;
 wire sw_405_data_out;
 wire sw_405_latch_out;
 wire \sw_405_module_data_in[0] ;
 wire \sw_405_module_data_in[1] ;
 wire \sw_405_module_data_in[2] ;
 wire \sw_405_module_data_in[3] ;
 wire \sw_405_module_data_in[4] ;
 wire \sw_405_module_data_in[5] ;
 wire \sw_405_module_data_in[6] ;
 wire \sw_405_module_data_in[7] ;
 wire \sw_405_module_data_out[0] ;
 wire \sw_405_module_data_out[1] ;
 wire \sw_405_module_data_out[2] ;
 wire \sw_405_module_data_out[3] ;
 wire \sw_405_module_data_out[4] ;
 wire \sw_405_module_data_out[5] ;
 wire \sw_405_module_data_out[6] ;
 wire \sw_405_module_data_out[7] ;
 wire sw_405_scan_out;
 wire sw_406_clk_out;
 wire sw_406_data_out;
 wire sw_406_latch_out;
 wire \sw_406_module_data_in[0] ;
 wire \sw_406_module_data_in[1] ;
 wire \sw_406_module_data_in[2] ;
 wire \sw_406_module_data_in[3] ;
 wire \sw_406_module_data_in[4] ;
 wire \sw_406_module_data_in[5] ;
 wire \sw_406_module_data_in[6] ;
 wire \sw_406_module_data_in[7] ;
 wire \sw_406_module_data_out[0] ;
 wire \sw_406_module_data_out[1] ;
 wire \sw_406_module_data_out[2] ;
 wire \sw_406_module_data_out[3] ;
 wire \sw_406_module_data_out[4] ;
 wire \sw_406_module_data_out[5] ;
 wire \sw_406_module_data_out[6] ;
 wire \sw_406_module_data_out[7] ;
 wire sw_406_scan_out;
 wire sw_407_clk_out;
 wire sw_407_data_out;
 wire sw_407_latch_out;
 wire \sw_407_module_data_in[0] ;
 wire \sw_407_module_data_in[1] ;
 wire \sw_407_module_data_in[2] ;
 wire \sw_407_module_data_in[3] ;
 wire \sw_407_module_data_in[4] ;
 wire \sw_407_module_data_in[5] ;
 wire \sw_407_module_data_in[6] ;
 wire \sw_407_module_data_in[7] ;
 wire \sw_407_module_data_out[0] ;
 wire \sw_407_module_data_out[1] ;
 wire \sw_407_module_data_out[2] ;
 wire \sw_407_module_data_out[3] ;
 wire \sw_407_module_data_out[4] ;
 wire \sw_407_module_data_out[5] ;
 wire \sw_407_module_data_out[6] ;
 wire \sw_407_module_data_out[7] ;
 wire sw_407_scan_out;
 wire sw_408_clk_out;
 wire sw_408_data_out;
 wire sw_408_latch_out;
 wire \sw_408_module_data_in[0] ;
 wire \sw_408_module_data_in[1] ;
 wire \sw_408_module_data_in[2] ;
 wire \sw_408_module_data_in[3] ;
 wire \sw_408_module_data_in[4] ;
 wire \sw_408_module_data_in[5] ;
 wire \sw_408_module_data_in[6] ;
 wire \sw_408_module_data_in[7] ;
 wire \sw_408_module_data_out[0] ;
 wire \sw_408_module_data_out[1] ;
 wire \sw_408_module_data_out[2] ;
 wire \sw_408_module_data_out[3] ;
 wire \sw_408_module_data_out[4] ;
 wire \sw_408_module_data_out[5] ;
 wire \sw_408_module_data_out[6] ;
 wire \sw_408_module_data_out[7] ;
 wire sw_408_scan_out;
 wire sw_409_clk_out;
 wire sw_409_data_out;
 wire sw_409_latch_out;
 wire \sw_409_module_data_in[0] ;
 wire \sw_409_module_data_in[1] ;
 wire \sw_409_module_data_in[2] ;
 wire \sw_409_module_data_in[3] ;
 wire \sw_409_module_data_in[4] ;
 wire \sw_409_module_data_in[5] ;
 wire \sw_409_module_data_in[6] ;
 wire \sw_409_module_data_in[7] ;
 wire \sw_409_module_data_out[0] ;
 wire \sw_409_module_data_out[1] ;
 wire \sw_409_module_data_out[2] ;
 wire \sw_409_module_data_out[3] ;
 wire \sw_409_module_data_out[4] ;
 wire \sw_409_module_data_out[5] ;
 wire \sw_409_module_data_out[6] ;
 wire \sw_409_module_data_out[7] ;
 wire sw_409_scan_out;
 wire sw_410_clk_out;
 wire sw_410_data_out;
 wire sw_410_latch_out;
 wire \sw_410_module_data_in[0] ;
 wire \sw_410_module_data_in[1] ;
 wire \sw_410_module_data_in[2] ;
 wire \sw_410_module_data_in[3] ;
 wire \sw_410_module_data_in[4] ;
 wire \sw_410_module_data_in[5] ;
 wire \sw_410_module_data_in[6] ;
 wire \sw_410_module_data_in[7] ;
 wire \sw_410_module_data_out[0] ;
 wire \sw_410_module_data_out[1] ;
 wire \sw_410_module_data_out[2] ;
 wire \sw_410_module_data_out[3] ;
 wire \sw_410_module_data_out[4] ;
 wire \sw_410_module_data_out[5] ;
 wire \sw_410_module_data_out[6] ;
 wire \sw_410_module_data_out[7] ;
 wire sw_410_scan_out;
 wire sw_411_clk_out;
 wire sw_411_data_out;
 wire sw_411_latch_out;
 wire \sw_411_module_data_in[0] ;
 wire \sw_411_module_data_in[1] ;
 wire \sw_411_module_data_in[2] ;
 wire \sw_411_module_data_in[3] ;
 wire \sw_411_module_data_in[4] ;
 wire \sw_411_module_data_in[5] ;
 wire \sw_411_module_data_in[6] ;
 wire \sw_411_module_data_in[7] ;
 wire \sw_411_module_data_out[0] ;
 wire \sw_411_module_data_out[1] ;
 wire \sw_411_module_data_out[2] ;
 wire \sw_411_module_data_out[3] ;
 wire \sw_411_module_data_out[4] ;
 wire \sw_411_module_data_out[5] ;
 wire \sw_411_module_data_out[6] ;
 wire \sw_411_module_data_out[7] ;
 wire sw_411_scan_out;
 wire sw_412_clk_out;
 wire sw_412_data_out;
 wire sw_412_latch_out;
 wire \sw_412_module_data_in[0] ;
 wire \sw_412_module_data_in[1] ;
 wire \sw_412_module_data_in[2] ;
 wire \sw_412_module_data_in[3] ;
 wire \sw_412_module_data_in[4] ;
 wire \sw_412_module_data_in[5] ;
 wire \sw_412_module_data_in[6] ;
 wire \sw_412_module_data_in[7] ;
 wire \sw_412_module_data_out[0] ;
 wire \sw_412_module_data_out[1] ;
 wire \sw_412_module_data_out[2] ;
 wire \sw_412_module_data_out[3] ;
 wire \sw_412_module_data_out[4] ;
 wire \sw_412_module_data_out[5] ;
 wire \sw_412_module_data_out[6] ;
 wire \sw_412_module_data_out[7] ;
 wire sw_412_scan_out;
 wire sw_413_clk_out;
 wire sw_413_data_out;
 wire sw_413_latch_out;
 wire \sw_413_module_data_in[0] ;
 wire \sw_413_module_data_in[1] ;
 wire \sw_413_module_data_in[2] ;
 wire \sw_413_module_data_in[3] ;
 wire \sw_413_module_data_in[4] ;
 wire \sw_413_module_data_in[5] ;
 wire \sw_413_module_data_in[6] ;
 wire \sw_413_module_data_in[7] ;
 wire \sw_413_module_data_out[0] ;
 wire \sw_413_module_data_out[1] ;
 wire \sw_413_module_data_out[2] ;
 wire \sw_413_module_data_out[3] ;
 wire \sw_413_module_data_out[4] ;
 wire \sw_413_module_data_out[5] ;
 wire \sw_413_module_data_out[6] ;
 wire \sw_413_module_data_out[7] ;
 wire sw_413_scan_out;
 wire sw_414_clk_out;
 wire sw_414_data_out;
 wire sw_414_latch_out;
 wire \sw_414_module_data_in[0] ;
 wire \sw_414_module_data_in[1] ;
 wire \sw_414_module_data_in[2] ;
 wire \sw_414_module_data_in[3] ;
 wire \sw_414_module_data_in[4] ;
 wire \sw_414_module_data_in[5] ;
 wire \sw_414_module_data_in[6] ;
 wire \sw_414_module_data_in[7] ;
 wire \sw_414_module_data_out[0] ;
 wire \sw_414_module_data_out[1] ;
 wire \sw_414_module_data_out[2] ;
 wire \sw_414_module_data_out[3] ;
 wire \sw_414_module_data_out[4] ;
 wire \sw_414_module_data_out[5] ;
 wire \sw_414_module_data_out[6] ;
 wire \sw_414_module_data_out[7] ;
 wire sw_414_scan_out;
 wire sw_415_clk_out;
 wire sw_415_data_out;
 wire sw_415_latch_out;
 wire \sw_415_module_data_in[0] ;
 wire \sw_415_module_data_in[1] ;
 wire \sw_415_module_data_in[2] ;
 wire \sw_415_module_data_in[3] ;
 wire \sw_415_module_data_in[4] ;
 wire \sw_415_module_data_in[5] ;
 wire \sw_415_module_data_in[6] ;
 wire \sw_415_module_data_in[7] ;
 wire \sw_415_module_data_out[0] ;
 wire \sw_415_module_data_out[1] ;
 wire \sw_415_module_data_out[2] ;
 wire \sw_415_module_data_out[3] ;
 wire \sw_415_module_data_out[4] ;
 wire \sw_415_module_data_out[5] ;
 wire \sw_415_module_data_out[6] ;
 wire \sw_415_module_data_out[7] ;
 wire sw_415_scan_out;
 wire sw_416_clk_out;
 wire sw_416_data_out;
 wire sw_416_latch_out;
 wire \sw_416_module_data_in[0] ;
 wire \sw_416_module_data_in[1] ;
 wire \sw_416_module_data_in[2] ;
 wire \sw_416_module_data_in[3] ;
 wire \sw_416_module_data_in[4] ;
 wire \sw_416_module_data_in[5] ;
 wire \sw_416_module_data_in[6] ;
 wire \sw_416_module_data_in[7] ;
 wire \sw_416_module_data_out[0] ;
 wire \sw_416_module_data_out[1] ;
 wire \sw_416_module_data_out[2] ;
 wire \sw_416_module_data_out[3] ;
 wire \sw_416_module_data_out[4] ;
 wire \sw_416_module_data_out[5] ;
 wire \sw_416_module_data_out[6] ;
 wire \sw_416_module_data_out[7] ;
 wire sw_416_scan_out;
 wire sw_417_clk_out;
 wire sw_417_data_out;
 wire sw_417_latch_out;
 wire \sw_417_module_data_in[0] ;
 wire \sw_417_module_data_in[1] ;
 wire \sw_417_module_data_in[2] ;
 wire \sw_417_module_data_in[3] ;
 wire \sw_417_module_data_in[4] ;
 wire \sw_417_module_data_in[5] ;
 wire \sw_417_module_data_in[6] ;
 wire \sw_417_module_data_in[7] ;
 wire \sw_417_module_data_out[0] ;
 wire \sw_417_module_data_out[1] ;
 wire \sw_417_module_data_out[2] ;
 wire \sw_417_module_data_out[3] ;
 wire \sw_417_module_data_out[4] ;
 wire \sw_417_module_data_out[5] ;
 wire \sw_417_module_data_out[6] ;
 wire \sw_417_module_data_out[7] ;
 wire sw_417_scan_out;
 wire sw_418_clk_out;
 wire sw_418_data_out;
 wire sw_418_latch_out;
 wire \sw_418_module_data_in[0] ;
 wire \sw_418_module_data_in[1] ;
 wire \sw_418_module_data_in[2] ;
 wire \sw_418_module_data_in[3] ;
 wire \sw_418_module_data_in[4] ;
 wire \sw_418_module_data_in[5] ;
 wire \sw_418_module_data_in[6] ;
 wire \sw_418_module_data_in[7] ;
 wire \sw_418_module_data_out[0] ;
 wire \sw_418_module_data_out[1] ;
 wire \sw_418_module_data_out[2] ;
 wire \sw_418_module_data_out[3] ;
 wire \sw_418_module_data_out[4] ;
 wire \sw_418_module_data_out[5] ;
 wire \sw_418_module_data_out[6] ;
 wire \sw_418_module_data_out[7] ;
 wire sw_418_scan_out;
 wire sw_419_clk_out;
 wire sw_419_data_out;
 wire sw_419_latch_out;
 wire \sw_419_module_data_in[0] ;
 wire \sw_419_module_data_in[1] ;
 wire \sw_419_module_data_in[2] ;
 wire \sw_419_module_data_in[3] ;
 wire \sw_419_module_data_in[4] ;
 wire \sw_419_module_data_in[5] ;
 wire \sw_419_module_data_in[6] ;
 wire \sw_419_module_data_in[7] ;
 wire \sw_419_module_data_out[0] ;
 wire \sw_419_module_data_out[1] ;
 wire \sw_419_module_data_out[2] ;
 wire \sw_419_module_data_out[3] ;
 wire \sw_419_module_data_out[4] ;
 wire \sw_419_module_data_out[5] ;
 wire \sw_419_module_data_out[6] ;
 wire \sw_419_module_data_out[7] ;
 wire sw_419_scan_out;
 wire sw_420_clk_out;
 wire sw_420_data_out;
 wire sw_420_latch_out;
 wire \sw_420_module_data_in[0] ;
 wire \sw_420_module_data_in[1] ;
 wire \sw_420_module_data_in[2] ;
 wire \sw_420_module_data_in[3] ;
 wire \sw_420_module_data_in[4] ;
 wire \sw_420_module_data_in[5] ;
 wire \sw_420_module_data_in[6] ;
 wire \sw_420_module_data_in[7] ;
 wire \sw_420_module_data_out[0] ;
 wire \sw_420_module_data_out[1] ;
 wire \sw_420_module_data_out[2] ;
 wire \sw_420_module_data_out[3] ;
 wire \sw_420_module_data_out[4] ;
 wire \sw_420_module_data_out[5] ;
 wire \sw_420_module_data_out[6] ;
 wire \sw_420_module_data_out[7] ;
 wire sw_420_scan_out;
 wire sw_421_clk_out;
 wire sw_421_data_out;
 wire sw_421_latch_out;
 wire \sw_421_module_data_in[0] ;
 wire \sw_421_module_data_in[1] ;
 wire \sw_421_module_data_in[2] ;
 wire \sw_421_module_data_in[3] ;
 wire \sw_421_module_data_in[4] ;
 wire \sw_421_module_data_in[5] ;
 wire \sw_421_module_data_in[6] ;
 wire \sw_421_module_data_in[7] ;
 wire \sw_421_module_data_out[0] ;
 wire \sw_421_module_data_out[1] ;
 wire \sw_421_module_data_out[2] ;
 wire \sw_421_module_data_out[3] ;
 wire \sw_421_module_data_out[4] ;
 wire \sw_421_module_data_out[5] ;
 wire \sw_421_module_data_out[6] ;
 wire \sw_421_module_data_out[7] ;
 wire sw_421_scan_out;
 wire sw_422_clk_out;
 wire sw_422_data_out;
 wire sw_422_latch_out;
 wire \sw_422_module_data_in[0] ;
 wire \sw_422_module_data_in[1] ;
 wire \sw_422_module_data_in[2] ;
 wire \sw_422_module_data_in[3] ;
 wire \sw_422_module_data_in[4] ;
 wire \sw_422_module_data_in[5] ;
 wire \sw_422_module_data_in[6] ;
 wire \sw_422_module_data_in[7] ;
 wire \sw_422_module_data_out[0] ;
 wire \sw_422_module_data_out[1] ;
 wire \sw_422_module_data_out[2] ;
 wire \sw_422_module_data_out[3] ;
 wire \sw_422_module_data_out[4] ;
 wire \sw_422_module_data_out[5] ;
 wire \sw_422_module_data_out[6] ;
 wire \sw_422_module_data_out[7] ;
 wire sw_422_scan_out;
 wire sw_423_clk_out;
 wire sw_423_data_out;
 wire sw_423_latch_out;
 wire \sw_423_module_data_in[0] ;
 wire \sw_423_module_data_in[1] ;
 wire \sw_423_module_data_in[2] ;
 wire \sw_423_module_data_in[3] ;
 wire \sw_423_module_data_in[4] ;
 wire \sw_423_module_data_in[5] ;
 wire \sw_423_module_data_in[6] ;
 wire \sw_423_module_data_in[7] ;
 wire \sw_423_module_data_out[0] ;
 wire \sw_423_module_data_out[1] ;
 wire \sw_423_module_data_out[2] ;
 wire \sw_423_module_data_out[3] ;
 wire \sw_423_module_data_out[4] ;
 wire \sw_423_module_data_out[5] ;
 wire \sw_423_module_data_out[6] ;
 wire \sw_423_module_data_out[7] ;
 wire sw_423_scan_out;
 wire sw_424_clk_out;
 wire sw_424_data_out;
 wire sw_424_latch_out;
 wire \sw_424_module_data_in[0] ;
 wire \sw_424_module_data_in[1] ;
 wire \sw_424_module_data_in[2] ;
 wire \sw_424_module_data_in[3] ;
 wire \sw_424_module_data_in[4] ;
 wire \sw_424_module_data_in[5] ;
 wire \sw_424_module_data_in[6] ;
 wire \sw_424_module_data_in[7] ;
 wire \sw_424_module_data_out[0] ;
 wire \sw_424_module_data_out[1] ;
 wire \sw_424_module_data_out[2] ;
 wire \sw_424_module_data_out[3] ;
 wire \sw_424_module_data_out[4] ;
 wire \sw_424_module_data_out[5] ;
 wire \sw_424_module_data_out[6] ;
 wire \sw_424_module_data_out[7] ;
 wire sw_424_scan_out;
 wire sw_425_clk_out;
 wire sw_425_data_out;
 wire sw_425_latch_out;
 wire \sw_425_module_data_in[0] ;
 wire \sw_425_module_data_in[1] ;
 wire \sw_425_module_data_in[2] ;
 wire \sw_425_module_data_in[3] ;
 wire \sw_425_module_data_in[4] ;
 wire \sw_425_module_data_in[5] ;
 wire \sw_425_module_data_in[6] ;
 wire \sw_425_module_data_in[7] ;
 wire \sw_425_module_data_out[0] ;
 wire \sw_425_module_data_out[1] ;
 wire \sw_425_module_data_out[2] ;
 wire \sw_425_module_data_out[3] ;
 wire \sw_425_module_data_out[4] ;
 wire \sw_425_module_data_out[5] ;
 wire \sw_425_module_data_out[6] ;
 wire \sw_425_module_data_out[7] ;
 wire sw_425_scan_out;
 wire sw_426_clk_out;
 wire sw_426_data_out;
 wire sw_426_latch_out;
 wire \sw_426_module_data_in[0] ;
 wire \sw_426_module_data_in[1] ;
 wire \sw_426_module_data_in[2] ;
 wire \sw_426_module_data_in[3] ;
 wire \sw_426_module_data_in[4] ;
 wire \sw_426_module_data_in[5] ;
 wire \sw_426_module_data_in[6] ;
 wire \sw_426_module_data_in[7] ;
 wire \sw_426_module_data_out[0] ;
 wire \sw_426_module_data_out[1] ;
 wire \sw_426_module_data_out[2] ;
 wire \sw_426_module_data_out[3] ;
 wire \sw_426_module_data_out[4] ;
 wire \sw_426_module_data_out[5] ;
 wire \sw_426_module_data_out[6] ;
 wire \sw_426_module_data_out[7] ;
 wire sw_426_scan_out;
 wire sw_427_clk_out;
 wire sw_427_data_out;
 wire sw_427_latch_out;
 wire \sw_427_module_data_in[0] ;
 wire \sw_427_module_data_in[1] ;
 wire \sw_427_module_data_in[2] ;
 wire \sw_427_module_data_in[3] ;
 wire \sw_427_module_data_in[4] ;
 wire \sw_427_module_data_in[5] ;
 wire \sw_427_module_data_in[6] ;
 wire \sw_427_module_data_in[7] ;
 wire \sw_427_module_data_out[0] ;
 wire \sw_427_module_data_out[1] ;
 wire \sw_427_module_data_out[2] ;
 wire \sw_427_module_data_out[3] ;
 wire \sw_427_module_data_out[4] ;
 wire \sw_427_module_data_out[5] ;
 wire \sw_427_module_data_out[6] ;
 wire \sw_427_module_data_out[7] ;
 wire sw_427_scan_out;
 wire sw_428_clk_out;
 wire sw_428_data_out;
 wire sw_428_latch_out;
 wire \sw_428_module_data_in[0] ;
 wire \sw_428_module_data_in[1] ;
 wire \sw_428_module_data_in[2] ;
 wire \sw_428_module_data_in[3] ;
 wire \sw_428_module_data_in[4] ;
 wire \sw_428_module_data_in[5] ;
 wire \sw_428_module_data_in[6] ;
 wire \sw_428_module_data_in[7] ;
 wire \sw_428_module_data_out[0] ;
 wire \sw_428_module_data_out[1] ;
 wire \sw_428_module_data_out[2] ;
 wire \sw_428_module_data_out[3] ;
 wire \sw_428_module_data_out[4] ;
 wire \sw_428_module_data_out[5] ;
 wire \sw_428_module_data_out[6] ;
 wire \sw_428_module_data_out[7] ;
 wire sw_428_scan_out;
 wire sw_429_clk_out;
 wire sw_429_data_out;
 wire sw_429_latch_out;
 wire \sw_429_module_data_in[0] ;
 wire \sw_429_module_data_in[1] ;
 wire \sw_429_module_data_in[2] ;
 wire \sw_429_module_data_in[3] ;
 wire \sw_429_module_data_in[4] ;
 wire \sw_429_module_data_in[5] ;
 wire \sw_429_module_data_in[6] ;
 wire \sw_429_module_data_in[7] ;
 wire \sw_429_module_data_out[0] ;
 wire \sw_429_module_data_out[1] ;
 wire \sw_429_module_data_out[2] ;
 wire \sw_429_module_data_out[3] ;
 wire \sw_429_module_data_out[4] ;
 wire \sw_429_module_data_out[5] ;
 wire \sw_429_module_data_out[6] ;
 wire \sw_429_module_data_out[7] ;
 wire sw_429_scan_out;
 wire sw_430_clk_out;
 wire sw_430_data_out;
 wire sw_430_latch_out;
 wire \sw_430_module_data_in[0] ;
 wire \sw_430_module_data_in[1] ;
 wire \sw_430_module_data_in[2] ;
 wire \sw_430_module_data_in[3] ;
 wire \sw_430_module_data_in[4] ;
 wire \sw_430_module_data_in[5] ;
 wire \sw_430_module_data_in[6] ;
 wire \sw_430_module_data_in[7] ;
 wire \sw_430_module_data_out[0] ;
 wire \sw_430_module_data_out[1] ;
 wire \sw_430_module_data_out[2] ;
 wire \sw_430_module_data_out[3] ;
 wire \sw_430_module_data_out[4] ;
 wire \sw_430_module_data_out[5] ;
 wire \sw_430_module_data_out[6] ;
 wire \sw_430_module_data_out[7] ;
 wire sw_430_scan_out;
 wire sw_431_clk_out;
 wire sw_431_data_out;
 wire sw_431_latch_out;
 wire \sw_431_module_data_in[0] ;
 wire \sw_431_module_data_in[1] ;
 wire \sw_431_module_data_in[2] ;
 wire \sw_431_module_data_in[3] ;
 wire \sw_431_module_data_in[4] ;
 wire \sw_431_module_data_in[5] ;
 wire \sw_431_module_data_in[6] ;
 wire \sw_431_module_data_in[7] ;
 wire \sw_431_module_data_out[0] ;
 wire \sw_431_module_data_out[1] ;
 wire \sw_431_module_data_out[2] ;
 wire \sw_431_module_data_out[3] ;
 wire \sw_431_module_data_out[4] ;
 wire \sw_431_module_data_out[5] ;
 wire \sw_431_module_data_out[6] ;
 wire \sw_431_module_data_out[7] ;
 wire sw_431_scan_out;
 wire sw_432_clk_out;
 wire sw_432_data_out;
 wire sw_432_latch_out;
 wire \sw_432_module_data_in[0] ;
 wire \sw_432_module_data_in[1] ;
 wire \sw_432_module_data_in[2] ;
 wire \sw_432_module_data_in[3] ;
 wire \sw_432_module_data_in[4] ;
 wire \sw_432_module_data_in[5] ;
 wire \sw_432_module_data_in[6] ;
 wire \sw_432_module_data_in[7] ;
 wire \sw_432_module_data_out[0] ;
 wire \sw_432_module_data_out[1] ;
 wire \sw_432_module_data_out[2] ;
 wire \sw_432_module_data_out[3] ;
 wire \sw_432_module_data_out[4] ;
 wire \sw_432_module_data_out[5] ;
 wire \sw_432_module_data_out[6] ;
 wire \sw_432_module_data_out[7] ;
 wire sw_432_scan_out;
 wire sw_433_clk_out;
 wire sw_433_data_out;
 wire sw_433_latch_out;
 wire \sw_433_module_data_in[0] ;
 wire \sw_433_module_data_in[1] ;
 wire \sw_433_module_data_in[2] ;
 wire \sw_433_module_data_in[3] ;
 wire \sw_433_module_data_in[4] ;
 wire \sw_433_module_data_in[5] ;
 wire \sw_433_module_data_in[6] ;
 wire \sw_433_module_data_in[7] ;
 wire \sw_433_module_data_out[0] ;
 wire \sw_433_module_data_out[1] ;
 wire \sw_433_module_data_out[2] ;
 wire \sw_433_module_data_out[3] ;
 wire \sw_433_module_data_out[4] ;
 wire \sw_433_module_data_out[5] ;
 wire \sw_433_module_data_out[6] ;
 wire \sw_433_module_data_out[7] ;
 wire sw_433_scan_out;
 wire sw_434_clk_out;
 wire sw_434_data_out;
 wire sw_434_latch_out;
 wire \sw_434_module_data_in[0] ;
 wire \sw_434_module_data_in[1] ;
 wire \sw_434_module_data_in[2] ;
 wire \sw_434_module_data_in[3] ;
 wire \sw_434_module_data_in[4] ;
 wire \sw_434_module_data_in[5] ;
 wire \sw_434_module_data_in[6] ;
 wire \sw_434_module_data_in[7] ;
 wire \sw_434_module_data_out[0] ;
 wire \sw_434_module_data_out[1] ;
 wire \sw_434_module_data_out[2] ;
 wire \sw_434_module_data_out[3] ;
 wire \sw_434_module_data_out[4] ;
 wire \sw_434_module_data_out[5] ;
 wire \sw_434_module_data_out[6] ;
 wire \sw_434_module_data_out[7] ;
 wire sw_434_scan_out;
 wire sw_435_clk_out;
 wire sw_435_data_out;
 wire sw_435_latch_out;
 wire \sw_435_module_data_in[0] ;
 wire \sw_435_module_data_in[1] ;
 wire \sw_435_module_data_in[2] ;
 wire \sw_435_module_data_in[3] ;
 wire \sw_435_module_data_in[4] ;
 wire \sw_435_module_data_in[5] ;
 wire \sw_435_module_data_in[6] ;
 wire \sw_435_module_data_in[7] ;
 wire \sw_435_module_data_out[0] ;
 wire \sw_435_module_data_out[1] ;
 wire \sw_435_module_data_out[2] ;
 wire \sw_435_module_data_out[3] ;
 wire \sw_435_module_data_out[4] ;
 wire \sw_435_module_data_out[5] ;
 wire \sw_435_module_data_out[6] ;
 wire \sw_435_module_data_out[7] ;
 wire sw_435_scan_out;
 wire sw_436_clk_out;
 wire sw_436_data_out;
 wire sw_436_latch_out;
 wire \sw_436_module_data_in[0] ;
 wire \sw_436_module_data_in[1] ;
 wire \sw_436_module_data_in[2] ;
 wire \sw_436_module_data_in[3] ;
 wire \sw_436_module_data_in[4] ;
 wire \sw_436_module_data_in[5] ;
 wire \sw_436_module_data_in[6] ;
 wire \sw_436_module_data_in[7] ;
 wire \sw_436_module_data_out[0] ;
 wire \sw_436_module_data_out[1] ;
 wire \sw_436_module_data_out[2] ;
 wire \sw_436_module_data_out[3] ;
 wire \sw_436_module_data_out[4] ;
 wire \sw_436_module_data_out[5] ;
 wire \sw_436_module_data_out[6] ;
 wire \sw_436_module_data_out[7] ;
 wire sw_436_scan_out;
 wire sw_437_clk_out;
 wire sw_437_data_out;
 wire sw_437_latch_out;
 wire \sw_437_module_data_in[0] ;
 wire \sw_437_module_data_in[1] ;
 wire \sw_437_module_data_in[2] ;
 wire \sw_437_module_data_in[3] ;
 wire \sw_437_module_data_in[4] ;
 wire \sw_437_module_data_in[5] ;
 wire \sw_437_module_data_in[6] ;
 wire \sw_437_module_data_in[7] ;
 wire \sw_437_module_data_out[0] ;
 wire \sw_437_module_data_out[1] ;
 wire \sw_437_module_data_out[2] ;
 wire \sw_437_module_data_out[3] ;
 wire \sw_437_module_data_out[4] ;
 wire \sw_437_module_data_out[5] ;
 wire \sw_437_module_data_out[6] ;
 wire \sw_437_module_data_out[7] ;
 wire sw_437_scan_out;
 wire sw_438_clk_out;
 wire sw_438_data_out;
 wire sw_438_latch_out;
 wire \sw_438_module_data_in[0] ;
 wire \sw_438_module_data_in[1] ;
 wire \sw_438_module_data_in[2] ;
 wire \sw_438_module_data_in[3] ;
 wire \sw_438_module_data_in[4] ;
 wire \sw_438_module_data_in[5] ;
 wire \sw_438_module_data_in[6] ;
 wire \sw_438_module_data_in[7] ;
 wire \sw_438_module_data_out[0] ;
 wire \sw_438_module_data_out[1] ;
 wire \sw_438_module_data_out[2] ;
 wire \sw_438_module_data_out[3] ;
 wire \sw_438_module_data_out[4] ;
 wire \sw_438_module_data_out[5] ;
 wire \sw_438_module_data_out[6] ;
 wire \sw_438_module_data_out[7] ;
 wire sw_438_scan_out;
 wire sw_439_clk_out;
 wire sw_439_data_out;
 wire sw_439_latch_out;
 wire \sw_439_module_data_in[0] ;
 wire \sw_439_module_data_in[1] ;
 wire \sw_439_module_data_in[2] ;
 wire \sw_439_module_data_in[3] ;
 wire \sw_439_module_data_in[4] ;
 wire \sw_439_module_data_in[5] ;
 wire \sw_439_module_data_in[6] ;
 wire \sw_439_module_data_in[7] ;
 wire \sw_439_module_data_out[0] ;
 wire \sw_439_module_data_out[1] ;
 wire \sw_439_module_data_out[2] ;
 wire \sw_439_module_data_out[3] ;
 wire \sw_439_module_data_out[4] ;
 wire \sw_439_module_data_out[5] ;
 wire \sw_439_module_data_out[6] ;
 wire \sw_439_module_data_out[7] ;
 wire sw_439_scan_out;
 wire sw_440_clk_out;
 wire sw_440_data_out;
 wire sw_440_latch_out;
 wire \sw_440_module_data_in[0] ;
 wire \sw_440_module_data_in[1] ;
 wire \sw_440_module_data_in[2] ;
 wire \sw_440_module_data_in[3] ;
 wire \sw_440_module_data_in[4] ;
 wire \sw_440_module_data_in[5] ;
 wire \sw_440_module_data_in[6] ;
 wire \sw_440_module_data_in[7] ;
 wire \sw_440_module_data_out[0] ;
 wire \sw_440_module_data_out[1] ;
 wire \sw_440_module_data_out[2] ;
 wire \sw_440_module_data_out[3] ;
 wire \sw_440_module_data_out[4] ;
 wire \sw_440_module_data_out[5] ;
 wire \sw_440_module_data_out[6] ;
 wire \sw_440_module_data_out[7] ;
 wire sw_440_scan_out;
 wire sw_441_clk_out;
 wire sw_441_data_out;
 wire sw_441_latch_out;
 wire \sw_441_module_data_in[0] ;
 wire \sw_441_module_data_in[1] ;
 wire \sw_441_module_data_in[2] ;
 wire \sw_441_module_data_in[3] ;
 wire \sw_441_module_data_in[4] ;
 wire \sw_441_module_data_in[5] ;
 wire \sw_441_module_data_in[6] ;
 wire \sw_441_module_data_in[7] ;
 wire \sw_441_module_data_out[0] ;
 wire \sw_441_module_data_out[1] ;
 wire \sw_441_module_data_out[2] ;
 wire \sw_441_module_data_out[3] ;
 wire \sw_441_module_data_out[4] ;
 wire \sw_441_module_data_out[5] ;
 wire \sw_441_module_data_out[6] ;
 wire \sw_441_module_data_out[7] ;
 wire sw_441_scan_out;
 wire sw_442_clk_out;
 wire sw_442_data_out;
 wire sw_442_latch_out;
 wire \sw_442_module_data_in[0] ;
 wire \sw_442_module_data_in[1] ;
 wire \sw_442_module_data_in[2] ;
 wire \sw_442_module_data_in[3] ;
 wire \sw_442_module_data_in[4] ;
 wire \sw_442_module_data_in[5] ;
 wire \sw_442_module_data_in[6] ;
 wire \sw_442_module_data_in[7] ;
 wire \sw_442_module_data_out[0] ;
 wire \sw_442_module_data_out[1] ;
 wire \sw_442_module_data_out[2] ;
 wire \sw_442_module_data_out[3] ;
 wire \sw_442_module_data_out[4] ;
 wire \sw_442_module_data_out[5] ;
 wire \sw_442_module_data_out[6] ;
 wire \sw_442_module_data_out[7] ;
 wire sw_442_scan_out;
 wire sw_443_clk_out;
 wire sw_443_data_out;
 wire sw_443_latch_out;
 wire \sw_443_module_data_in[0] ;
 wire \sw_443_module_data_in[1] ;
 wire \sw_443_module_data_in[2] ;
 wire \sw_443_module_data_in[3] ;
 wire \sw_443_module_data_in[4] ;
 wire \sw_443_module_data_in[5] ;
 wire \sw_443_module_data_in[6] ;
 wire \sw_443_module_data_in[7] ;
 wire \sw_443_module_data_out[0] ;
 wire \sw_443_module_data_out[1] ;
 wire \sw_443_module_data_out[2] ;
 wire \sw_443_module_data_out[3] ;
 wire \sw_443_module_data_out[4] ;
 wire \sw_443_module_data_out[5] ;
 wire \sw_443_module_data_out[6] ;
 wire \sw_443_module_data_out[7] ;
 wire sw_443_scan_out;
 wire sw_444_clk_out;
 wire sw_444_data_out;
 wire sw_444_latch_out;
 wire \sw_444_module_data_in[0] ;
 wire \sw_444_module_data_in[1] ;
 wire \sw_444_module_data_in[2] ;
 wire \sw_444_module_data_in[3] ;
 wire \sw_444_module_data_in[4] ;
 wire \sw_444_module_data_in[5] ;
 wire \sw_444_module_data_in[6] ;
 wire \sw_444_module_data_in[7] ;
 wire \sw_444_module_data_out[0] ;
 wire \sw_444_module_data_out[1] ;
 wire \sw_444_module_data_out[2] ;
 wire \sw_444_module_data_out[3] ;
 wire \sw_444_module_data_out[4] ;
 wire \sw_444_module_data_out[5] ;
 wire \sw_444_module_data_out[6] ;
 wire \sw_444_module_data_out[7] ;
 wire sw_444_scan_out;
 wire sw_445_clk_out;
 wire sw_445_data_out;
 wire sw_445_latch_out;
 wire \sw_445_module_data_in[0] ;
 wire \sw_445_module_data_in[1] ;
 wire \sw_445_module_data_in[2] ;
 wire \sw_445_module_data_in[3] ;
 wire \sw_445_module_data_in[4] ;
 wire \sw_445_module_data_in[5] ;
 wire \sw_445_module_data_in[6] ;
 wire \sw_445_module_data_in[7] ;
 wire \sw_445_module_data_out[0] ;
 wire \sw_445_module_data_out[1] ;
 wire \sw_445_module_data_out[2] ;
 wire \sw_445_module_data_out[3] ;
 wire \sw_445_module_data_out[4] ;
 wire \sw_445_module_data_out[5] ;
 wire \sw_445_module_data_out[6] ;
 wire \sw_445_module_data_out[7] ;
 wire sw_445_scan_out;
 wire sw_446_clk_out;
 wire sw_446_data_out;
 wire sw_446_latch_out;
 wire \sw_446_module_data_in[0] ;
 wire \sw_446_module_data_in[1] ;
 wire \sw_446_module_data_in[2] ;
 wire \sw_446_module_data_in[3] ;
 wire \sw_446_module_data_in[4] ;
 wire \sw_446_module_data_in[5] ;
 wire \sw_446_module_data_in[6] ;
 wire \sw_446_module_data_in[7] ;
 wire \sw_446_module_data_out[0] ;
 wire \sw_446_module_data_out[1] ;
 wire \sw_446_module_data_out[2] ;
 wire \sw_446_module_data_out[3] ;
 wire \sw_446_module_data_out[4] ;
 wire \sw_446_module_data_out[5] ;
 wire \sw_446_module_data_out[6] ;
 wire \sw_446_module_data_out[7] ;
 wire sw_446_scan_out;
 wire sw_447_clk_out;
 wire sw_447_data_out;
 wire sw_447_latch_out;
 wire \sw_447_module_data_in[0] ;
 wire \sw_447_module_data_in[1] ;
 wire \sw_447_module_data_in[2] ;
 wire \sw_447_module_data_in[3] ;
 wire \sw_447_module_data_in[4] ;
 wire \sw_447_module_data_in[5] ;
 wire \sw_447_module_data_in[6] ;
 wire \sw_447_module_data_in[7] ;
 wire \sw_447_module_data_out[0] ;
 wire \sw_447_module_data_out[1] ;
 wire \sw_447_module_data_out[2] ;
 wire \sw_447_module_data_out[3] ;
 wire \sw_447_module_data_out[4] ;
 wire \sw_447_module_data_out[5] ;
 wire \sw_447_module_data_out[6] ;
 wire \sw_447_module_data_out[7] ;
 wire sw_447_scan_out;
 wire sw_448_clk_out;
 wire sw_448_data_out;
 wire sw_448_latch_out;
 wire \sw_448_module_data_in[0] ;
 wire \sw_448_module_data_in[1] ;
 wire \sw_448_module_data_in[2] ;
 wire \sw_448_module_data_in[3] ;
 wire \sw_448_module_data_in[4] ;
 wire \sw_448_module_data_in[5] ;
 wire \sw_448_module_data_in[6] ;
 wire \sw_448_module_data_in[7] ;
 wire \sw_448_module_data_out[0] ;
 wire \sw_448_module_data_out[1] ;
 wire \sw_448_module_data_out[2] ;
 wire \sw_448_module_data_out[3] ;
 wire \sw_448_module_data_out[4] ;
 wire \sw_448_module_data_out[5] ;
 wire \sw_448_module_data_out[6] ;
 wire \sw_448_module_data_out[7] ;
 wire sw_448_scan_out;
 wire sw_449_clk_out;
 wire sw_449_data_out;
 wire sw_449_latch_out;
 wire \sw_449_module_data_in[0] ;
 wire \sw_449_module_data_in[1] ;
 wire \sw_449_module_data_in[2] ;
 wire \sw_449_module_data_in[3] ;
 wire \sw_449_module_data_in[4] ;
 wire \sw_449_module_data_in[5] ;
 wire \sw_449_module_data_in[6] ;
 wire \sw_449_module_data_in[7] ;
 wire \sw_449_module_data_out[0] ;
 wire \sw_449_module_data_out[1] ;
 wire \sw_449_module_data_out[2] ;
 wire \sw_449_module_data_out[3] ;
 wire \sw_449_module_data_out[4] ;
 wire \sw_449_module_data_out[5] ;
 wire \sw_449_module_data_out[6] ;
 wire \sw_449_module_data_out[7] ;
 wire sw_449_scan_out;
 wire sw_450_clk_out;
 wire sw_450_data_out;
 wire sw_450_latch_out;
 wire \sw_450_module_data_in[0] ;
 wire \sw_450_module_data_in[1] ;
 wire \sw_450_module_data_in[2] ;
 wire \sw_450_module_data_in[3] ;
 wire \sw_450_module_data_in[4] ;
 wire \sw_450_module_data_in[5] ;
 wire \sw_450_module_data_in[6] ;
 wire \sw_450_module_data_in[7] ;
 wire \sw_450_module_data_out[0] ;
 wire \sw_450_module_data_out[1] ;
 wire \sw_450_module_data_out[2] ;
 wire \sw_450_module_data_out[3] ;
 wire \sw_450_module_data_out[4] ;
 wire \sw_450_module_data_out[5] ;
 wire \sw_450_module_data_out[6] ;
 wire \sw_450_module_data_out[7] ;
 wire sw_450_scan_out;
 wire sw_451_clk_out;
 wire sw_451_data_out;
 wire sw_451_latch_out;
 wire \sw_451_module_data_in[0] ;
 wire \sw_451_module_data_in[1] ;
 wire \sw_451_module_data_in[2] ;
 wire \sw_451_module_data_in[3] ;
 wire \sw_451_module_data_in[4] ;
 wire \sw_451_module_data_in[5] ;
 wire \sw_451_module_data_in[6] ;
 wire \sw_451_module_data_in[7] ;
 wire \sw_451_module_data_out[0] ;
 wire \sw_451_module_data_out[1] ;
 wire \sw_451_module_data_out[2] ;
 wire \sw_451_module_data_out[3] ;
 wire \sw_451_module_data_out[4] ;
 wire \sw_451_module_data_out[5] ;
 wire \sw_451_module_data_out[6] ;
 wire \sw_451_module_data_out[7] ;
 wire sw_451_scan_out;
 wire sw_452_clk_out;
 wire sw_452_data_out;
 wire sw_452_latch_out;
 wire \sw_452_module_data_in[0] ;
 wire \sw_452_module_data_in[1] ;
 wire \sw_452_module_data_in[2] ;
 wire \sw_452_module_data_in[3] ;
 wire \sw_452_module_data_in[4] ;
 wire \sw_452_module_data_in[5] ;
 wire \sw_452_module_data_in[6] ;
 wire \sw_452_module_data_in[7] ;
 wire \sw_452_module_data_out[0] ;
 wire \sw_452_module_data_out[1] ;
 wire \sw_452_module_data_out[2] ;
 wire \sw_452_module_data_out[3] ;
 wire \sw_452_module_data_out[4] ;
 wire \sw_452_module_data_out[5] ;
 wire \sw_452_module_data_out[6] ;
 wire \sw_452_module_data_out[7] ;
 wire sw_452_scan_out;
 wire sw_453_clk_out;
 wire sw_453_data_out;
 wire sw_453_latch_out;
 wire \sw_453_module_data_in[0] ;
 wire \sw_453_module_data_in[1] ;
 wire \sw_453_module_data_in[2] ;
 wire \sw_453_module_data_in[3] ;
 wire \sw_453_module_data_in[4] ;
 wire \sw_453_module_data_in[5] ;
 wire \sw_453_module_data_in[6] ;
 wire \sw_453_module_data_in[7] ;
 wire \sw_453_module_data_out[0] ;
 wire \sw_453_module_data_out[1] ;
 wire \sw_453_module_data_out[2] ;
 wire \sw_453_module_data_out[3] ;
 wire \sw_453_module_data_out[4] ;
 wire \sw_453_module_data_out[5] ;
 wire \sw_453_module_data_out[6] ;
 wire \sw_453_module_data_out[7] ;
 wire sw_453_scan_out;
 wire sw_454_clk_out;
 wire sw_454_data_out;
 wire sw_454_latch_out;
 wire \sw_454_module_data_in[0] ;
 wire \sw_454_module_data_in[1] ;
 wire \sw_454_module_data_in[2] ;
 wire \sw_454_module_data_in[3] ;
 wire \sw_454_module_data_in[4] ;
 wire \sw_454_module_data_in[5] ;
 wire \sw_454_module_data_in[6] ;
 wire \sw_454_module_data_in[7] ;
 wire \sw_454_module_data_out[0] ;
 wire \sw_454_module_data_out[1] ;
 wire \sw_454_module_data_out[2] ;
 wire \sw_454_module_data_out[3] ;
 wire \sw_454_module_data_out[4] ;
 wire \sw_454_module_data_out[5] ;
 wire \sw_454_module_data_out[6] ;
 wire \sw_454_module_data_out[7] ;
 wire sw_454_scan_out;
 wire sw_455_clk_out;
 wire sw_455_data_out;
 wire sw_455_latch_out;
 wire \sw_455_module_data_in[0] ;
 wire \sw_455_module_data_in[1] ;
 wire \sw_455_module_data_in[2] ;
 wire \sw_455_module_data_in[3] ;
 wire \sw_455_module_data_in[4] ;
 wire \sw_455_module_data_in[5] ;
 wire \sw_455_module_data_in[6] ;
 wire \sw_455_module_data_in[7] ;
 wire \sw_455_module_data_out[0] ;
 wire \sw_455_module_data_out[1] ;
 wire \sw_455_module_data_out[2] ;
 wire \sw_455_module_data_out[3] ;
 wire \sw_455_module_data_out[4] ;
 wire \sw_455_module_data_out[5] ;
 wire \sw_455_module_data_out[6] ;
 wire \sw_455_module_data_out[7] ;
 wire sw_455_scan_out;
 wire sw_456_clk_out;
 wire sw_456_data_out;
 wire sw_456_latch_out;
 wire \sw_456_module_data_in[0] ;
 wire \sw_456_module_data_in[1] ;
 wire \sw_456_module_data_in[2] ;
 wire \sw_456_module_data_in[3] ;
 wire \sw_456_module_data_in[4] ;
 wire \sw_456_module_data_in[5] ;
 wire \sw_456_module_data_in[6] ;
 wire \sw_456_module_data_in[7] ;
 wire \sw_456_module_data_out[0] ;
 wire \sw_456_module_data_out[1] ;
 wire \sw_456_module_data_out[2] ;
 wire \sw_456_module_data_out[3] ;
 wire \sw_456_module_data_out[4] ;
 wire \sw_456_module_data_out[5] ;
 wire \sw_456_module_data_out[6] ;
 wire \sw_456_module_data_out[7] ;
 wire sw_456_scan_out;
 wire sw_457_clk_out;
 wire sw_457_data_out;
 wire sw_457_latch_out;
 wire \sw_457_module_data_in[0] ;
 wire \sw_457_module_data_in[1] ;
 wire \sw_457_module_data_in[2] ;
 wire \sw_457_module_data_in[3] ;
 wire \sw_457_module_data_in[4] ;
 wire \sw_457_module_data_in[5] ;
 wire \sw_457_module_data_in[6] ;
 wire \sw_457_module_data_in[7] ;
 wire \sw_457_module_data_out[0] ;
 wire \sw_457_module_data_out[1] ;
 wire \sw_457_module_data_out[2] ;
 wire \sw_457_module_data_out[3] ;
 wire \sw_457_module_data_out[4] ;
 wire \sw_457_module_data_out[5] ;
 wire \sw_457_module_data_out[6] ;
 wire \sw_457_module_data_out[7] ;
 wire sw_457_scan_out;
 wire sw_458_clk_out;
 wire sw_458_data_out;
 wire sw_458_latch_out;
 wire \sw_458_module_data_in[0] ;
 wire \sw_458_module_data_in[1] ;
 wire \sw_458_module_data_in[2] ;
 wire \sw_458_module_data_in[3] ;
 wire \sw_458_module_data_in[4] ;
 wire \sw_458_module_data_in[5] ;
 wire \sw_458_module_data_in[6] ;
 wire \sw_458_module_data_in[7] ;
 wire \sw_458_module_data_out[0] ;
 wire \sw_458_module_data_out[1] ;
 wire \sw_458_module_data_out[2] ;
 wire \sw_458_module_data_out[3] ;
 wire \sw_458_module_data_out[4] ;
 wire \sw_458_module_data_out[5] ;
 wire \sw_458_module_data_out[6] ;
 wire \sw_458_module_data_out[7] ;
 wire sw_458_scan_out;
 wire sw_459_clk_out;
 wire sw_459_data_out;
 wire sw_459_latch_out;
 wire \sw_459_module_data_in[0] ;
 wire \sw_459_module_data_in[1] ;
 wire \sw_459_module_data_in[2] ;
 wire \sw_459_module_data_in[3] ;
 wire \sw_459_module_data_in[4] ;
 wire \sw_459_module_data_in[5] ;
 wire \sw_459_module_data_in[6] ;
 wire \sw_459_module_data_in[7] ;
 wire \sw_459_module_data_out[0] ;
 wire \sw_459_module_data_out[1] ;
 wire \sw_459_module_data_out[2] ;
 wire \sw_459_module_data_out[3] ;
 wire \sw_459_module_data_out[4] ;
 wire \sw_459_module_data_out[5] ;
 wire \sw_459_module_data_out[6] ;
 wire \sw_459_module_data_out[7] ;
 wire sw_459_scan_out;
 wire sw_460_clk_out;
 wire sw_460_data_out;
 wire sw_460_latch_out;
 wire \sw_460_module_data_in[0] ;
 wire \sw_460_module_data_in[1] ;
 wire \sw_460_module_data_in[2] ;
 wire \sw_460_module_data_in[3] ;
 wire \sw_460_module_data_in[4] ;
 wire \sw_460_module_data_in[5] ;
 wire \sw_460_module_data_in[6] ;
 wire \sw_460_module_data_in[7] ;
 wire \sw_460_module_data_out[0] ;
 wire \sw_460_module_data_out[1] ;
 wire \sw_460_module_data_out[2] ;
 wire \sw_460_module_data_out[3] ;
 wire \sw_460_module_data_out[4] ;
 wire \sw_460_module_data_out[5] ;
 wire \sw_460_module_data_out[6] ;
 wire \sw_460_module_data_out[7] ;
 wire sw_460_scan_out;
 wire sw_461_clk_out;
 wire sw_461_data_out;
 wire sw_461_latch_out;
 wire \sw_461_module_data_in[0] ;
 wire \sw_461_module_data_in[1] ;
 wire \sw_461_module_data_in[2] ;
 wire \sw_461_module_data_in[3] ;
 wire \sw_461_module_data_in[4] ;
 wire \sw_461_module_data_in[5] ;
 wire \sw_461_module_data_in[6] ;
 wire \sw_461_module_data_in[7] ;
 wire \sw_461_module_data_out[0] ;
 wire \sw_461_module_data_out[1] ;
 wire \sw_461_module_data_out[2] ;
 wire \sw_461_module_data_out[3] ;
 wire \sw_461_module_data_out[4] ;
 wire \sw_461_module_data_out[5] ;
 wire \sw_461_module_data_out[6] ;
 wire \sw_461_module_data_out[7] ;
 wire sw_461_scan_out;
 wire sw_462_clk_out;
 wire sw_462_data_out;
 wire sw_462_latch_out;
 wire \sw_462_module_data_in[0] ;
 wire \sw_462_module_data_in[1] ;
 wire \sw_462_module_data_in[2] ;
 wire \sw_462_module_data_in[3] ;
 wire \sw_462_module_data_in[4] ;
 wire \sw_462_module_data_in[5] ;
 wire \sw_462_module_data_in[6] ;
 wire \sw_462_module_data_in[7] ;
 wire \sw_462_module_data_out[0] ;
 wire \sw_462_module_data_out[1] ;
 wire \sw_462_module_data_out[2] ;
 wire \sw_462_module_data_out[3] ;
 wire \sw_462_module_data_out[4] ;
 wire \sw_462_module_data_out[5] ;
 wire \sw_462_module_data_out[6] ;
 wire \sw_462_module_data_out[7] ;
 wire sw_462_scan_out;
 wire sw_463_clk_out;
 wire sw_463_data_out;
 wire sw_463_latch_out;
 wire \sw_463_module_data_in[0] ;
 wire \sw_463_module_data_in[1] ;
 wire \sw_463_module_data_in[2] ;
 wire \sw_463_module_data_in[3] ;
 wire \sw_463_module_data_in[4] ;
 wire \sw_463_module_data_in[5] ;
 wire \sw_463_module_data_in[6] ;
 wire \sw_463_module_data_in[7] ;
 wire \sw_463_module_data_out[0] ;
 wire \sw_463_module_data_out[1] ;
 wire \sw_463_module_data_out[2] ;
 wire \sw_463_module_data_out[3] ;
 wire \sw_463_module_data_out[4] ;
 wire \sw_463_module_data_out[5] ;
 wire \sw_463_module_data_out[6] ;
 wire \sw_463_module_data_out[7] ;
 wire sw_463_scan_out;
 wire sw_464_clk_out;
 wire sw_464_data_out;
 wire sw_464_latch_out;
 wire \sw_464_module_data_in[0] ;
 wire \sw_464_module_data_in[1] ;
 wire \sw_464_module_data_in[2] ;
 wire \sw_464_module_data_in[3] ;
 wire \sw_464_module_data_in[4] ;
 wire \sw_464_module_data_in[5] ;
 wire \sw_464_module_data_in[6] ;
 wire \sw_464_module_data_in[7] ;
 wire \sw_464_module_data_out[0] ;
 wire \sw_464_module_data_out[1] ;
 wire \sw_464_module_data_out[2] ;
 wire \sw_464_module_data_out[3] ;
 wire \sw_464_module_data_out[4] ;
 wire \sw_464_module_data_out[5] ;
 wire \sw_464_module_data_out[6] ;
 wire \sw_464_module_data_out[7] ;
 wire sw_464_scan_out;
 wire sw_465_clk_out;
 wire sw_465_data_out;
 wire sw_465_latch_out;
 wire \sw_465_module_data_in[0] ;
 wire \sw_465_module_data_in[1] ;
 wire \sw_465_module_data_in[2] ;
 wire \sw_465_module_data_in[3] ;
 wire \sw_465_module_data_in[4] ;
 wire \sw_465_module_data_in[5] ;
 wire \sw_465_module_data_in[6] ;
 wire \sw_465_module_data_in[7] ;
 wire \sw_465_module_data_out[0] ;
 wire \sw_465_module_data_out[1] ;
 wire \sw_465_module_data_out[2] ;
 wire \sw_465_module_data_out[3] ;
 wire \sw_465_module_data_out[4] ;
 wire \sw_465_module_data_out[5] ;
 wire \sw_465_module_data_out[6] ;
 wire \sw_465_module_data_out[7] ;
 wire sw_465_scan_out;
 wire sw_466_clk_out;
 wire sw_466_data_out;
 wire sw_466_latch_out;
 wire \sw_466_module_data_in[0] ;
 wire \sw_466_module_data_in[1] ;
 wire \sw_466_module_data_in[2] ;
 wire \sw_466_module_data_in[3] ;
 wire \sw_466_module_data_in[4] ;
 wire \sw_466_module_data_in[5] ;
 wire \sw_466_module_data_in[6] ;
 wire \sw_466_module_data_in[7] ;
 wire \sw_466_module_data_out[0] ;
 wire \sw_466_module_data_out[1] ;
 wire \sw_466_module_data_out[2] ;
 wire \sw_466_module_data_out[3] ;
 wire \sw_466_module_data_out[4] ;
 wire \sw_466_module_data_out[5] ;
 wire \sw_466_module_data_out[6] ;
 wire \sw_466_module_data_out[7] ;
 wire sw_466_scan_out;
 wire sw_467_clk_out;
 wire sw_467_data_out;
 wire sw_467_latch_out;
 wire \sw_467_module_data_in[0] ;
 wire \sw_467_module_data_in[1] ;
 wire \sw_467_module_data_in[2] ;
 wire \sw_467_module_data_in[3] ;
 wire \sw_467_module_data_in[4] ;
 wire \sw_467_module_data_in[5] ;
 wire \sw_467_module_data_in[6] ;
 wire \sw_467_module_data_in[7] ;
 wire \sw_467_module_data_out[0] ;
 wire \sw_467_module_data_out[1] ;
 wire \sw_467_module_data_out[2] ;
 wire \sw_467_module_data_out[3] ;
 wire \sw_467_module_data_out[4] ;
 wire \sw_467_module_data_out[5] ;
 wire \sw_467_module_data_out[6] ;
 wire \sw_467_module_data_out[7] ;
 wire sw_467_scan_out;
 wire sw_468_clk_out;
 wire sw_468_data_out;
 wire sw_468_latch_out;
 wire \sw_468_module_data_in[0] ;
 wire \sw_468_module_data_in[1] ;
 wire \sw_468_module_data_in[2] ;
 wire \sw_468_module_data_in[3] ;
 wire \sw_468_module_data_in[4] ;
 wire \sw_468_module_data_in[5] ;
 wire \sw_468_module_data_in[6] ;
 wire \sw_468_module_data_in[7] ;
 wire \sw_468_module_data_out[0] ;
 wire \sw_468_module_data_out[1] ;
 wire \sw_468_module_data_out[2] ;
 wire \sw_468_module_data_out[3] ;
 wire \sw_468_module_data_out[4] ;
 wire \sw_468_module_data_out[5] ;
 wire \sw_468_module_data_out[6] ;
 wire \sw_468_module_data_out[7] ;
 wire sw_468_scan_out;
 wire sw_469_clk_out;
 wire sw_469_data_out;
 wire sw_469_latch_out;
 wire \sw_469_module_data_in[0] ;
 wire \sw_469_module_data_in[1] ;
 wire \sw_469_module_data_in[2] ;
 wire \sw_469_module_data_in[3] ;
 wire \sw_469_module_data_in[4] ;
 wire \sw_469_module_data_in[5] ;
 wire \sw_469_module_data_in[6] ;
 wire \sw_469_module_data_in[7] ;
 wire \sw_469_module_data_out[0] ;
 wire \sw_469_module_data_out[1] ;
 wire \sw_469_module_data_out[2] ;
 wire \sw_469_module_data_out[3] ;
 wire \sw_469_module_data_out[4] ;
 wire \sw_469_module_data_out[5] ;
 wire \sw_469_module_data_out[6] ;
 wire \sw_469_module_data_out[7] ;
 wire sw_469_scan_out;
 wire sw_470_clk_out;
 wire sw_470_data_out;
 wire sw_470_latch_out;
 wire \sw_470_module_data_in[0] ;
 wire \sw_470_module_data_in[1] ;
 wire \sw_470_module_data_in[2] ;
 wire \sw_470_module_data_in[3] ;
 wire \sw_470_module_data_in[4] ;
 wire \sw_470_module_data_in[5] ;
 wire \sw_470_module_data_in[6] ;
 wire \sw_470_module_data_in[7] ;
 wire \sw_470_module_data_out[0] ;
 wire \sw_470_module_data_out[1] ;
 wire \sw_470_module_data_out[2] ;
 wire \sw_470_module_data_out[3] ;
 wire \sw_470_module_data_out[4] ;
 wire \sw_470_module_data_out[5] ;
 wire \sw_470_module_data_out[6] ;
 wire \sw_470_module_data_out[7] ;
 wire sw_470_scan_out;
 wire sw_471_clk_out;
 wire sw_471_data_out;
 wire sw_471_latch_out;
 wire \sw_471_module_data_in[0] ;
 wire \sw_471_module_data_in[1] ;
 wire \sw_471_module_data_in[2] ;
 wire \sw_471_module_data_in[3] ;
 wire \sw_471_module_data_in[4] ;
 wire \sw_471_module_data_in[5] ;
 wire \sw_471_module_data_in[6] ;
 wire \sw_471_module_data_in[7] ;
 wire \sw_471_module_data_out[0] ;
 wire \sw_471_module_data_out[1] ;
 wire \sw_471_module_data_out[2] ;
 wire \sw_471_module_data_out[3] ;
 wire \sw_471_module_data_out[4] ;
 wire \sw_471_module_data_out[5] ;
 wire \sw_471_module_data_out[6] ;
 wire \sw_471_module_data_out[7] ;
 wire sw_471_scan_out;
 wire sw_472_latch_out;
 wire \sw_472_module_data_in[0] ;
 wire \sw_472_module_data_in[1] ;
 wire \sw_472_module_data_in[2] ;
 wire \sw_472_module_data_in[3] ;
 wire \sw_472_module_data_in[4] ;
 wire \sw_472_module_data_in[5] ;
 wire \sw_472_module_data_in[6] ;
 wire \sw_472_module_data_in[7] ;
 wire \sw_472_module_data_out[0] ;
 wire \sw_472_module_data_out[1] ;
 wire \sw_472_module_data_out[2] ;
 wire \sw_472_module_data_out[3] ;
 wire \sw_472_module_data_out[4] ;
 wire \sw_472_module_data_out[5] ;
 wire \sw_472_module_data_out[6] ;
 wire \sw_472_module_data_out[7] ;
 wire sw_472_scan_out;

 aidan_McCoy aidan_McCoy_8 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_008_module_data_in[7] ,
    \sw_008_module_data_in[6] ,
    \sw_008_module_data_in[5] ,
    \sw_008_module_data_in[4] ,
    \sw_008_module_data_in[3] ,
    \sw_008_module_data_in[2] ,
    \sw_008_module_data_in[1] ,
    \sw_008_module_data_in[0] }),
    .io_out({\sw_008_module_data_out[7] ,
    \sw_008_module_data_out[6] ,
    \sw_008_module_data_out[5] ,
    \sw_008_module_data_out[4] ,
    \sw_008_module_data_out[3] ,
    \sw_008_module_data_out[2] ,
    \sw_008_module_data_out[1] ,
    \sw_008_module_data_out[0] }));
 alu_top alu_top_7 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_007_module_data_in[7] ,
    \sw_007_module_data_in[6] ,
    \sw_007_module_data_in[5] ,
    \sw_007_module_data_in[4] ,
    \sw_007_module_data_in[3] ,
    \sw_007_module_data_in[2] ,
    \sw_007_module_data_in[1] ,
    \sw_007_module_data_in[0] }),
    .io_out({\sw_007_module_data_out[7] ,
    \sw_007_module_data_out[6] ,
    \sw_007_module_data_out[5] ,
    \sw_007_module_data_out[4] ,
    \sw_007_module_data_out[3] ,
    \sw_007_module_data_out[2] ,
    \sw_007_module_data_out[1] ,
    \sw_007_module_data_out[0] }));
 asic_multiplier_wrapper asic_multiplier_wrapper_23 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_023_module_data_in[7] ,
    \sw_023_module_data_in[6] ,
    \sw_023_module_data_in[5] ,
    \sw_023_module_data_in[4] ,
    \sw_023_module_data_in[3] ,
    \sw_023_module_data_in[2] ,
    \sw_023_module_data_in[1] ,
    \sw_023_module_data_in[0] }),
    .io_out({\sw_023_module_data_out[7] ,
    \sw_023_module_data_out[6] ,
    \sw_023_module_data_out[5] ,
    \sw_023_module_data_out[4] ,
    \sw_023_module_data_out[3] ,
    \sw_023_module_data_out[2] ,
    \sw_023_module_data_out[1] ,
    \sw_023_module_data_out[0] }));
 azdle_binary_clock azdle_binary_clock_9 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_009_module_data_in[7] ,
    \sw_009_module_data_in[6] ,
    \sw_009_module_data_in[5] ,
    \sw_009_module_data_in[4] ,
    \sw_009_module_data_in[3] ,
    \sw_009_module_data_in[2] ,
    \sw_009_module_data_in[1] ,
    \sw_009_module_data_in[0] }),
    .io_out({\sw_009_module_data_out[7] ,
    \sw_009_module_data_out[6] ,
    \sw_009_module_data_out[5] ,
    \sw_009_module_data_out[4] ,
    \sw_009_module_data_out[3] ,
    \sw_009_module_data_out[2] ,
    \sw_009_module_data_out[1] ,
    \sw_009_module_data_out[0] }));
 chase_the_beat chase_the_beat_20 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_020_module_data_in[7] ,
    \sw_020_module_data_in[6] ,
    \sw_020_module_data_in[5] ,
    \sw_020_module_data_in[4] ,
    \sw_020_module_data_in[3] ,
    \sw_020_module_data_in[2] ,
    \sw_020_module_data_in[1] ,
    \sw_020_module_data_in[0] }),
    .io_out({\sw_020_module_data_out[7] ,
    \sw_020_module_data_out[6] ,
    \sw_020_module_data_out[5] ,
    \sw_020_module_data_out[4] ,
    \sw_020_module_data_out[3] ,
    \sw_020_module_data_out[2] ,
    \sw_020_module_data_out[1] ,
    \sw_020_module_data_out[0] }));
 chrisruk_matrix chrisruk_matrix_3 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_003_module_data_in[7] ,
    \sw_003_module_data_in[6] ,
    \sw_003_module_data_in[5] ,
    \sw_003_module_data_in[4] ,
    \sw_003_module_data_in[3] ,
    \sw_003_module_data_in[2] ,
    \sw_003_module_data_in[1] ,
    \sw_003_module_data_in[0] }),
    .io_out({\sw_003_module_data_out[7] ,
    \sw_003_module_data_out[6] ,
    \sw_003_module_data_out[5] ,
    \sw_003_module_data_out[4] ,
    \sw_003_module_data_out[3] ,
    \sw_003_module_data_out[2] ,
    \sw_003_module_data_out[1] ,
    \sw_003_module_data_out[0] }));
 fraserbc_simon fraserbc_simon_1 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_001_module_data_in[7] ,
    \sw_001_module_data_in[6] ,
    \sw_001_module_data_in[5] ,
    \sw_001_module_data_in[4] ,
    \sw_001_module_data_in[3] ,
    \sw_001_module_data_in[2] ,
    \sw_001_module_data_in[1] ,
    \sw_001_module_data_in[0] }),
    .io_out({\sw_001_module_data_out[7] ,
    \sw_001_module_data_out[6] ,
    \sw_001_module_data_out[5] ,
    \sw_001_module_data_out[4] ,
    \sw_001_module_data_out[3] ,
    \sw_001_module_data_out[2] ,
    \sw_001_module_data_out[1] ,
    \sw_001_module_data_out[0] }));
 jar_sram_top jar_sram_top_11 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_011_module_data_in[7] ,
    \sw_011_module_data_in[6] ,
    \sw_011_module_data_in[5] ,
    \sw_011_module_data_in[4] ,
    \sw_011_module_data_in[3] ,
    \sw_011_module_data_in[2] ,
    \sw_011_module_data_in[1] ,
    \sw_011_module_data_in[0] }),
    .io_out({\sw_011_module_data_out[7] ,
    \sw_011_module_data_out[6] ,
    \sw_011_module_data_out[5] ,
    \sw_011_module_data_out[4] ,
    \sw_011_module_data_out[3] ,
    \sw_011_module_data_out[2] ,
    \sw_011_module_data_out[1] ,
    \sw_011_module_data_out[0] }));
 loxodes_sequencer loxodes_sequencer_4 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_004_module_data_in[7] ,
    \sw_004_module_data_in[6] ,
    \sw_004_module_data_in[5] ,
    \sw_004_module_data_in[4] ,
    \sw_004_module_data_in[3] ,
    \sw_004_module_data_in[2] ,
    \sw_004_module_data_in[1] ,
    \sw_004_module_data_in[0] }),
    .io_out({\sw_004_module_data_out[7] ,
    \sw_004_module_data_out[6] ,
    \sw_004_module_data_out[5] ,
    \sw_004_module_data_out[4] ,
    \sw_004_module_data_out[3] ,
    \sw_004_module_data_out[2] ,
    \sw_004_module_data_out[1] ,
    \sw_004_module_data_out[0] }));
 migcorre_pwm migcorre_pwm_5 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_005_module_data_in[7] ,
    \sw_005_module_data_in[6] ,
    \sw_005_module_data_in[5] ,
    \sw_005_module_data_in[4] ,
    \sw_005_module_data_in[3] ,
    \sw_005_module_data_in[2] ,
    \sw_005_module_data_in[1] ,
    \sw_005_module_data_in[0] }),
    .io_out({\sw_005_module_data_out[7] ,
    \sw_005_module_data_out[6] ,
    \sw_005_module_data_out[5] ,
    \sw_005_module_data_out[4] ,
    \sw_005_module_data_out[3] ,
    \sw_005_module_data_out[2] ,
    \sw_005_module_data_out[1] ,
    \sw_005_module_data_out[0] }));
 mm21_LEDMatrixTop mm21_LEDMatrixTop_26 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_026_module_data_in[7] ,
    \sw_026_module_data_in[6] ,
    \sw_026_module_data_in[5] ,
    \sw_026_module_data_in[4] ,
    \sw_026_module_data_in[3] ,
    \sw_026_module_data_in[2] ,
    \sw_026_module_data_in[1] ,
    \sw_026_module_data_in[0] }),
    .io_out({\sw_026_module_data_out[7] ,
    \sw_026_module_data_out[6] ,
    \sw_026_module_data_out[5] ,
    \sw_026_module_data_out[4] ,
    \sw_026_module_data_out[3] ,
    \sw_026_module_data_out[2] ,
    \sw_026_module_data_out[1] ,
    \sw_026_module_data_out[0] }));
 s4ga s4ga_6 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_006_module_data_in[7] ,
    \sw_006_module_data_in[6] ,
    \sw_006_module_data_in[5] ,
    \sw_006_module_data_in[4] ,
    \sw_006_module_data_in[3] ,
    \sw_006_module_data_in[2] ,
    \sw_006_module_data_in[1] ,
    \sw_006_module_data_in[0] }),
    .io_out({\sw_006_module_data_out[7] ,
    \sw_006_module_data_out[6] ,
    \sw_006_module_data_out[5] ,
    \sw_006_module_data_out[4] ,
    \sw_006_module_data_out[3] ,
    \sw_006_module_data_out[2] ,
    \sw_006_module_data_out[1] ,
    \sw_006_module_data_out[0] }));
 scan_controller scan_controller (.clk(wb_clk_i),
    .la_scan_clk_in(la_data_in[0]),
    .la_scan_data_in(la_data_in[1]),
    .la_scan_data_out(la_data_out[0]),
    .la_scan_latch_en(la_data_in[3]),
    .la_scan_select(la_data_in[2]),
    .ready(io_out[37]),
    .reset(wb_rst_i),
    .scan_clk_in(sc_clk_in),
    .scan_clk_out(sc_clk_out),
    .scan_data_in(sc_data_in),
    .scan_data_out(sc_data_out),
    .scan_latch_en(sc_latch_out),
    .scan_select(sc_scan_out),
    .set_clk_div(io_in[11]),
    .slow_clk(io_out[10]),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .active_select({io_in[20],
    io_in[19],
    io_in[18],
    io_in[17],
    io_in[16],
    io_in[15],
    io_in[14],
    io_in[13],
    io_in[12]}),
    .driver_sel({io_in[9],
    io_in[8]}),
    .inputs({io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24],
    io_in[23],
    io_in[22],
    io_in[21]}),
    .oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .outputs({io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29]}));
 scanchain scanchain_0 (.clk_in(sc_clk_out),
    .clk_out(sw_000_clk_out),
    .data_in(sc_data_out),
    .data_out(sw_000_data_out),
    .latch_enable_in(sc_latch_out),
    .latch_enable_out(sw_000_latch_out),
    .scan_select_in(sc_scan_out),
    .scan_select_out(sw_000_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_000_module_data_in[7] ,
    \sw_000_module_data_in[6] ,
    \sw_000_module_data_in[5] ,
    \sw_000_module_data_in[4] ,
    \sw_000_module_data_in[3] ,
    \sw_000_module_data_in[2] ,
    \sw_000_module_data_in[1] ,
    \sw_000_module_data_in[0] }),
    .module_data_out({\sw_000_module_data_out[7] ,
    \sw_000_module_data_out[6] ,
    \sw_000_module_data_out[5] ,
    \sw_000_module_data_out[4] ,
    \sw_000_module_data_out[3] ,
    \sw_000_module_data_out[2] ,
    \sw_000_module_data_out[1] ,
    \sw_000_module_data_out[0] }));
 scanchain scanchain_1 (.clk_in(sw_000_clk_out),
    .clk_out(sw_001_clk_out),
    .data_in(sw_000_data_out),
    .data_out(sw_001_data_out),
    .latch_enable_in(sw_000_latch_out),
    .latch_enable_out(sw_001_latch_out),
    .scan_select_in(sw_000_scan_out),
    .scan_select_out(sw_001_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_001_module_data_in[7] ,
    \sw_001_module_data_in[6] ,
    \sw_001_module_data_in[5] ,
    \sw_001_module_data_in[4] ,
    \sw_001_module_data_in[3] ,
    \sw_001_module_data_in[2] ,
    \sw_001_module_data_in[1] ,
    \sw_001_module_data_in[0] }),
    .module_data_out({\sw_001_module_data_out[7] ,
    \sw_001_module_data_out[6] ,
    \sw_001_module_data_out[5] ,
    \sw_001_module_data_out[4] ,
    \sw_001_module_data_out[3] ,
    \sw_001_module_data_out[2] ,
    \sw_001_module_data_out[1] ,
    \sw_001_module_data_out[0] }));
 scanchain scanchain_10 (.clk_in(sw_009_clk_out),
    .clk_out(sw_010_clk_out),
    .data_in(sw_009_data_out),
    .data_out(sw_010_data_out),
    .latch_enable_in(sw_009_latch_out),
    .latch_enable_out(sw_010_latch_out),
    .scan_select_in(sw_009_scan_out),
    .scan_select_out(sw_010_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_010_module_data_in[7] ,
    \sw_010_module_data_in[6] ,
    \sw_010_module_data_in[5] ,
    \sw_010_module_data_in[4] ,
    \sw_010_module_data_in[3] ,
    \sw_010_module_data_in[2] ,
    \sw_010_module_data_in[1] ,
    \sw_010_module_data_in[0] }),
    .module_data_out({\sw_010_module_data_out[7] ,
    \sw_010_module_data_out[6] ,
    \sw_010_module_data_out[5] ,
    \sw_010_module_data_out[4] ,
    \sw_010_module_data_out[3] ,
    \sw_010_module_data_out[2] ,
    \sw_010_module_data_out[1] ,
    \sw_010_module_data_out[0] }));
 scanchain scanchain_100 (.clk_in(sw_099_clk_out),
    .clk_out(sw_100_clk_out),
    .data_in(sw_099_data_out),
    .data_out(sw_100_data_out),
    .latch_enable_in(sw_099_latch_out),
    .latch_enable_out(sw_100_latch_out),
    .scan_select_in(sw_099_scan_out),
    .scan_select_out(sw_100_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_100_module_data_in[7] ,
    \sw_100_module_data_in[6] ,
    \sw_100_module_data_in[5] ,
    \sw_100_module_data_in[4] ,
    \sw_100_module_data_in[3] ,
    \sw_100_module_data_in[2] ,
    \sw_100_module_data_in[1] ,
    \sw_100_module_data_in[0] }),
    .module_data_out({\sw_100_module_data_out[7] ,
    \sw_100_module_data_out[6] ,
    \sw_100_module_data_out[5] ,
    \sw_100_module_data_out[4] ,
    \sw_100_module_data_out[3] ,
    \sw_100_module_data_out[2] ,
    \sw_100_module_data_out[1] ,
    \sw_100_module_data_out[0] }));
 scanchain scanchain_101 (.clk_in(sw_100_clk_out),
    .clk_out(sw_101_clk_out),
    .data_in(sw_100_data_out),
    .data_out(sw_101_data_out),
    .latch_enable_in(sw_100_latch_out),
    .latch_enable_out(sw_101_latch_out),
    .scan_select_in(sw_100_scan_out),
    .scan_select_out(sw_101_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_101_module_data_in[7] ,
    \sw_101_module_data_in[6] ,
    \sw_101_module_data_in[5] ,
    \sw_101_module_data_in[4] ,
    \sw_101_module_data_in[3] ,
    \sw_101_module_data_in[2] ,
    \sw_101_module_data_in[1] ,
    \sw_101_module_data_in[0] }),
    .module_data_out({\sw_101_module_data_out[7] ,
    \sw_101_module_data_out[6] ,
    \sw_101_module_data_out[5] ,
    \sw_101_module_data_out[4] ,
    \sw_101_module_data_out[3] ,
    \sw_101_module_data_out[2] ,
    \sw_101_module_data_out[1] ,
    \sw_101_module_data_out[0] }));
 scanchain scanchain_102 (.clk_in(sw_101_clk_out),
    .clk_out(sw_102_clk_out),
    .data_in(sw_101_data_out),
    .data_out(sw_102_data_out),
    .latch_enable_in(sw_101_latch_out),
    .latch_enable_out(sw_102_latch_out),
    .scan_select_in(sw_101_scan_out),
    .scan_select_out(sw_102_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_102_module_data_in[7] ,
    \sw_102_module_data_in[6] ,
    \sw_102_module_data_in[5] ,
    \sw_102_module_data_in[4] ,
    \sw_102_module_data_in[3] ,
    \sw_102_module_data_in[2] ,
    \sw_102_module_data_in[1] ,
    \sw_102_module_data_in[0] }),
    .module_data_out({\sw_102_module_data_out[7] ,
    \sw_102_module_data_out[6] ,
    \sw_102_module_data_out[5] ,
    \sw_102_module_data_out[4] ,
    \sw_102_module_data_out[3] ,
    \sw_102_module_data_out[2] ,
    \sw_102_module_data_out[1] ,
    \sw_102_module_data_out[0] }));
 scanchain scanchain_103 (.clk_in(sw_102_clk_out),
    .clk_out(sw_103_clk_out),
    .data_in(sw_102_data_out),
    .data_out(sw_103_data_out),
    .latch_enable_in(sw_102_latch_out),
    .latch_enable_out(sw_103_latch_out),
    .scan_select_in(sw_102_scan_out),
    .scan_select_out(sw_103_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_103_module_data_in[7] ,
    \sw_103_module_data_in[6] ,
    \sw_103_module_data_in[5] ,
    \sw_103_module_data_in[4] ,
    \sw_103_module_data_in[3] ,
    \sw_103_module_data_in[2] ,
    \sw_103_module_data_in[1] ,
    \sw_103_module_data_in[0] }),
    .module_data_out({\sw_103_module_data_out[7] ,
    \sw_103_module_data_out[6] ,
    \sw_103_module_data_out[5] ,
    \sw_103_module_data_out[4] ,
    \sw_103_module_data_out[3] ,
    \sw_103_module_data_out[2] ,
    \sw_103_module_data_out[1] ,
    \sw_103_module_data_out[0] }));
 scanchain scanchain_104 (.clk_in(sw_103_clk_out),
    .clk_out(sw_104_clk_out),
    .data_in(sw_103_data_out),
    .data_out(sw_104_data_out),
    .latch_enable_in(sw_103_latch_out),
    .latch_enable_out(sw_104_latch_out),
    .scan_select_in(sw_103_scan_out),
    .scan_select_out(sw_104_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_104_module_data_in[7] ,
    \sw_104_module_data_in[6] ,
    \sw_104_module_data_in[5] ,
    \sw_104_module_data_in[4] ,
    \sw_104_module_data_in[3] ,
    \sw_104_module_data_in[2] ,
    \sw_104_module_data_in[1] ,
    \sw_104_module_data_in[0] }),
    .module_data_out({\sw_104_module_data_out[7] ,
    \sw_104_module_data_out[6] ,
    \sw_104_module_data_out[5] ,
    \sw_104_module_data_out[4] ,
    \sw_104_module_data_out[3] ,
    \sw_104_module_data_out[2] ,
    \sw_104_module_data_out[1] ,
    \sw_104_module_data_out[0] }));
 scanchain scanchain_105 (.clk_in(sw_104_clk_out),
    .clk_out(sw_105_clk_out),
    .data_in(sw_104_data_out),
    .data_out(sw_105_data_out),
    .latch_enable_in(sw_104_latch_out),
    .latch_enable_out(sw_105_latch_out),
    .scan_select_in(sw_104_scan_out),
    .scan_select_out(sw_105_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_105_module_data_in[7] ,
    \sw_105_module_data_in[6] ,
    \sw_105_module_data_in[5] ,
    \sw_105_module_data_in[4] ,
    \sw_105_module_data_in[3] ,
    \sw_105_module_data_in[2] ,
    \sw_105_module_data_in[1] ,
    \sw_105_module_data_in[0] }),
    .module_data_out({\sw_105_module_data_out[7] ,
    \sw_105_module_data_out[6] ,
    \sw_105_module_data_out[5] ,
    \sw_105_module_data_out[4] ,
    \sw_105_module_data_out[3] ,
    \sw_105_module_data_out[2] ,
    \sw_105_module_data_out[1] ,
    \sw_105_module_data_out[0] }));
 scanchain scanchain_106 (.clk_in(sw_105_clk_out),
    .clk_out(sw_106_clk_out),
    .data_in(sw_105_data_out),
    .data_out(sw_106_data_out),
    .latch_enable_in(sw_105_latch_out),
    .latch_enable_out(sw_106_latch_out),
    .scan_select_in(sw_105_scan_out),
    .scan_select_out(sw_106_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_106_module_data_in[7] ,
    \sw_106_module_data_in[6] ,
    \sw_106_module_data_in[5] ,
    \sw_106_module_data_in[4] ,
    \sw_106_module_data_in[3] ,
    \sw_106_module_data_in[2] ,
    \sw_106_module_data_in[1] ,
    \sw_106_module_data_in[0] }),
    .module_data_out({\sw_106_module_data_out[7] ,
    \sw_106_module_data_out[6] ,
    \sw_106_module_data_out[5] ,
    \sw_106_module_data_out[4] ,
    \sw_106_module_data_out[3] ,
    \sw_106_module_data_out[2] ,
    \sw_106_module_data_out[1] ,
    \sw_106_module_data_out[0] }));
 scanchain scanchain_107 (.clk_in(sw_106_clk_out),
    .clk_out(sw_107_clk_out),
    .data_in(sw_106_data_out),
    .data_out(sw_107_data_out),
    .latch_enable_in(sw_106_latch_out),
    .latch_enable_out(sw_107_latch_out),
    .scan_select_in(sw_106_scan_out),
    .scan_select_out(sw_107_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_107_module_data_in[7] ,
    \sw_107_module_data_in[6] ,
    \sw_107_module_data_in[5] ,
    \sw_107_module_data_in[4] ,
    \sw_107_module_data_in[3] ,
    \sw_107_module_data_in[2] ,
    \sw_107_module_data_in[1] ,
    \sw_107_module_data_in[0] }),
    .module_data_out({\sw_107_module_data_out[7] ,
    \sw_107_module_data_out[6] ,
    \sw_107_module_data_out[5] ,
    \sw_107_module_data_out[4] ,
    \sw_107_module_data_out[3] ,
    \sw_107_module_data_out[2] ,
    \sw_107_module_data_out[1] ,
    \sw_107_module_data_out[0] }));
 scanchain scanchain_108 (.clk_in(sw_107_clk_out),
    .clk_out(sw_108_clk_out),
    .data_in(sw_107_data_out),
    .data_out(sw_108_data_out),
    .latch_enable_in(sw_107_latch_out),
    .latch_enable_out(sw_108_latch_out),
    .scan_select_in(sw_107_scan_out),
    .scan_select_out(sw_108_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_108_module_data_in[7] ,
    \sw_108_module_data_in[6] ,
    \sw_108_module_data_in[5] ,
    \sw_108_module_data_in[4] ,
    \sw_108_module_data_in[3] ,
    \sw_108_module_data_in[2] ,
    \sw_108_module_data_in[1] ,
    \sw_108_module_data_in[0] }),
    .module_data_out({\sw_108_module_data_out[7] ,
    \sw_108_module_data_out[6] ,
    \sw_108_module_data_out[5] ,
    \sw_108_module_data_out[4] ,
    \sw_108_module_data_out[3] ,
    \sw_108_module_data_out[2] ,
    \sw_108_module_data_out[1] ,
    \sw_108_module_data_out[0] }));
 scanchain scanchain_109 (.clk_in(sw_108_clk_out),
    .clk_out(sw_109_clk_out),
    .data_in(sw_108_data_out),
    .data_out(sw_109_data_out),
    .latch_enable_in(sw_108_latch_out),
    .latch_enable_out(sw_109_latch_out),
    .scan_select_in(sw_108_scan_out),
    .scan_select_out(sw_109_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_109_module_data_in[7] ,
    \sw_109_module_data_in[6] ,
    \sw_109_module_data_in[5] ,
    \sw_109_module_data_in[4] ,
    \sw_109_module_data_in[3] ,
    \sw_109_module_data_in[2] ,
    \sw_109_module_data_in[1] ,
    \sw_109_module_data_in[0] }),
    .module_data_out({\sw_109_module_data_out[7] ,
    \sw_109_module_data_out[6] ,
    \sw_109_module_data_out[5] ,
    \sw_109_module_data_out[4] ,
    \sw_109_module_data_out[3] ,
    \sw_109_module_data_out[2] ,
    \sw_109_module_data_out[1] ,
    \sw_109_module_data_out[0] }));
 scanchain scanchain_11 (.clk_in(sw_010_clk_out),
    .clk_out(sw_011_clk_out),
    .data_in(sw_010_data_out),
    .data_out(sw_011_data_out),
    .latch_enable_in(sw_010_latch_out),
    .latch_enable_out(sw_011_latch_out),
    .scan_select_in(sw_010_scan_out),
    .scan_select_out(sw_011_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_011_module_data_in[7] ,
    \sw_011_module_data_in[6] ,
    \sw_011_module_data_in[5] ,
    \sw_011_module_data_in[4] ,
    \sw_011_module_data_in[3] ,
    \sw_011_module_data_in[2] ,
    \sw_011_module_data_in[1] ,
    \sw_011_module_data_in[0] }),
    .module_data_out({\sw_011_module_data_out[7] ,
    \sw_011_module_data_out[6] ,
    \sw_011_module_data_out[5] ,
    \sw_011_module_data_out[4] ,
    \sw_011_module_data_out[3] ,
    \sw_011_module_data_out[2] ,
    \sw_011_module_data_out[1] ,
    \sw_011_module_data_out[0] }));
 scanchain scanchain_110 (.clk_in(sw_109_clk_out),
    .clk_out(sw_110_clk_out),
    .data_in(sw_109_data_out),
    .data_out(sw_110_data_out),
    .latch_enable_in(sw_109_latch_out),
    .latch_enable_out(sw_110_latch_out),
    .scan_select_in(sw_109_scan_out),
    .scan_select_out(sw_110_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_110_module_data_in[7] ,
    \sw_110_module_data_in[6] ,
    \sw_110_module_data_in[5] ,
    \sw_110_module_data_in[4] ,
    \sw_110_module_data_in[3] ,
    \sw_110_module_data_in[2] ,
    \sw_110_module_data_in[1] ,
    \sw_110_module_data_in[0] }),
    .module_data_out({\sw_110_module_data_out[7] ,
    \sw_110_module_data_out[6] ,
    \sw_110_module_data_out[5] ,
    \sw_110_module_data_out[4] ,
    \sw_110_module_data_out[3] ,
    \sw_110_module_data_out[2] ,
    \sw_110_module_data_out[1] ,
    \sw_110_module_data_out[0] }));
 scanchain scanchain_111 (.clk_in(sw_110_clk_out),
    .clk_out(sw_111_clk_out),
    .data_in(sw_110_data_out),
    .data_out(sw_111_data_out),
    .latch_enable_in(sw_110_latch_out),
    .latch_enable_out(sw_111_latch_out),
    .scan_select_in(sw_110_scan_out),
    .scan_select_out(sw_111_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_111_module_data_in[7] ,
    \sw_111_module_data_in[6] ,
    \sw_111_module_data_in[5] ,
    \sw_111_module_data_in[4] ,
    \sw_111_module_data_in[3] ,
    \sw_111_module_data_in[2] ,
    \sw_111_module_data_in[1] ,
    \sw_111_module_data_in[0] }),
    .module_data_out({\sw_111_module_data_out[7] ,
    \sw_111_module_data_out[6] ,
    \sw_111_module_data_out[5] ,
    \sw_111_module_data_out[4] ,
    \sw_111_module_data_out[3] ,
    \sw_111_module_data_out[2] ,
    \sw_111_module_data_out[1] ,
    \sw_111_module_data_out[0] }));
 scanchain scanchain_112 (.clk_in(sw_111_clk_out),
    .clk_out(sw_112_clk_out),
    .data_in(sw_111_data_out),
    .data_out(sw_112_data_out),
    .latch_enable_in(sw_111_latch_out),
    .latch_enable_out(sw_112_latch_out),
    .scan_select_in(sw_111_scan_out),
    .scan_select_out(sw_112_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_112_module_data_in[7] ,
    \sw_112_module_data_in[6] ,
    \sw_112_module_data_in[5] ,
    \sw_112_module_data_in[4] ,
    \sw_112_module_data_in[3] ,
    \sw_112_module_data_in[2] ,
    \sw_112_module_data_in[1] ,
    \sw_112_module_data_in[0] }),
    .module_data_out({\sw_112_module_data_out[7] ,
    \sw_112_module_data_out[6] ,
    \sw_112_module_data_out[5] ,
    \sw_112_module_data_out[4] ,
    \sw_112_module_data_out[3] ,
    \sw_112_module_data_out[2] ,
    \sw_112_module_data_out[1] ,
    \sw_112_module_data_out[0] }));
 scanchain scanchain_113 (.clk_in(sw_112_clk_out),
    .clk_out(sw_113_clk_out),
    .data_in(sw_112_data_out),
    .data_out(sw_113_data_out),
    .latch_enable_in(sw_112_latch_out),
    .latch_enable_out(sw_113_latch_out),
    .scan_select_in(sw_112_scan_out),
    .scan_select_out(sw_113_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_113_module_data_in[7] ,
    \sw_113_module_data_in[6] ,
    \sw_113_module_data_in[5] ,
    \sw_113_module_data_in[4] ,
    \sw_113_module_data_in[3] ,
    \sw_113_module_data_in[2] ,
    \sw_113_module_data_in[1] ,
    \sw_113_module_data_in[0] }),
    .module_data_out({\sw_113_module_data_out[7] ,
    \sw_113_module_data_out[6] ,
    \sw_113_module_data_out[5] ,
    \sw_113_module_data_out[4] ,
    \sw_113_module_data_out[3] ,
    \sw_113_module_data_out[2] ,
    \sw_113_module_data_out[1] ,
    \sw_113_module_data_out[0] }));
 scanchain scanchain_114 (.clk_in(sw_113_clk_out),
    .clk_out(sw_114_clk_out),
    .data_in(sw_113_data_out),
    .data_out(sw_114_data_out),
    .latch_enable_in(sw_113_latch_out),
    .latch_enable_out(sw_114_latch_out),
    .scan_select_in(sw_113_scan_out),
    .scan_select_out(sw_114_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_114_module_data_in[7] ,
    \sw_114_module_data_in[6] ,
    \sw_114_module_data_in[5] ,
    \sw_114_module_data_in[4] ,
    \sw_114_module_data_in[3] ,
    \sw_114_module_data_in[2] ,
    \sw_114_module_data_in[1] ,
    \sw_114_module_data_in[0] }),
    .module_data_out({\sw_114_module_data_out[7] ,
    \sw_114_module_data_out[6] ,
    \sw_114_module_data_out[5] ,
    \sw_114_module_data_out[4] ,
    \sw_114_module_data_out[3] ,
    \sw_114_module_data_out[2] ,
    \sw_114_module_data_out[1] ,
    \sw_114_module_data_out[0] }));
 scanchain scanchain_115 (.clk_in(sw_114_clk_out),
    .clk_out(sw_115_clk_out),
    .data_in(sw_114_data_out),
    .data_out(sw_115_data_out),
    .latch_enable_in(sw_114_latch_out),
    .latch_enable_out(sw_115_latch_out),
    .scan_select_in(sw_114_scan_out),
    .scan_select_out(sw_115_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_115_module_data_in[7] ,
    \sw_115_module_data_in[6] ,
    \sw_115_module_data_in[5] ,
    \sw_115_module_data_in[4] ,
    \sw_115_module_data_in[3] ,
    \sw_115_module_data_in[2] ,
    \sw_115_module_data_in[1] ,
    \sw_115_module_data_in[0] }),
    .module_data_out({\sw_115_module_data_out[7] ,
    \sw_115_module_data_out[6] ,
    \sw_115_module_data_out[5] ,
    \sw_115_module_data_out[4] ,
    \sw_115_module_data_out[3] ,
    \sw_115_module_data_out[2] ,
    \sw_115_module_data_out[1] ,
    \sw_115_module_data_out[0] }));
 scanchain scanchain_116 (.clk_in(sw_115_clk_out),
    .clk_out(sw_116_clk_out),
    .data_in(sw_115_data_out),
    .data_out(sw_116_data_out),
    .latch_enable_in(sw_115_latch_out),
    .latch_enable_out(sw_116_latch_out),
    .scan_select_in(sw_115_scan_out),
    .scan_select_out(sw_116_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_116_module_data_in[7] ,
    \sw_116_module_data_in[6] ,
    \sw_116_module_data_in[5] ,
    \sw_116_module_data_in[4] ,
    \sw_116_module_data_in[3] ,
    \sw_116_module_data_in[2] ,
    \sw_116_module_data_in[1] ,
    \sw_116_module_data_in[0] }),
    .module_data_out({\sw_116_module_data_out[7] ,
    \sw_116_module_data_out[6] ,
    \sw_116_module_data_out[5] ,
    \sw_116_module_data_out[4] ,
    \sw_116_module_data_out[3] ,
    \sw_116_module_data_out[2] ,
    \sw_116_module_data_out[1] ,
    \sw_116_module_data_out[0] }));
 scanchain scanchain_117 (.clk_in(sw_116_clk_out),
    .clk_out(sw_117_clk_out),
    .data_in(sw_116_data_out),
    .data_out(sw_117_data_out),
    .latch_enable_in(sw_116_latch_out),
    .latch_enable_out(sw_117_latch_out),
    .scan_select_in(sw_116_scan_out),
    .scan_select_out(sw_117_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_117_module_data_in[7] ,
    \sw_117_module_data_in[6] ,
    \sw_117_module_data_in[5] ,
    \sw_117_module_data_in[4] ,
    \sw_117_module_data_in[3] ,
    \sw_117_module_data_in[2] ,
    \sw_117_module_data_in[1] ,
    \sw_117_module_data_in[0] }),
    .module_data_out({\sw_117_module_data_out[7] ,
    \sw_117_module_data_out[6] ,
    \sw_117_module_data_out[5] ,
    \sw_117_module_data_out[4] ,
    \sw_117_module_data_out[3] ,
    \sw_117_module_data_out[2] ,
    \sw_117_module_data_out[1] ,
    \sw_117_module_data_out[0] }));
 scanchain scanchain_118 (.clk_in(sw_117_clk_out),
    .clk_out(sw_118_clk_out),
    .data_in(sw_117_data_out),
    .data_out(sw_118_data_out),
    .latch_enable_in(sw_117_latch_out),
    .latch_enable_out(sw_118_latch_out),
    .scan_select_in(sw_117_scan_out),
    .scan_select_out(sw_118_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_118_module_data_in[7] ,
    \sw_118_module_data_in[6] ,
    \sw_118_module_data_in[5] ,
    \sw_118_module_data_in[4] ,
    \sw_118_module_data_in[3] ,
    \sw_118_module_data_in[2] ,
    \sw_118_module_data_in[1] ,
    \sw_118_module_data_in[0] }),
    .module_data_out({\sw_118_module_data_out[7] ,
    \sw_118_module_data_out[6] ,
    \sw_118_module_data_out[5] ,
    \sw_118_module_data_out[4] ,
    \sw_118_module_data_out[3] ,
    \sw_118_module_data_out[2] ,
    \sw_118_module_data_out[1] ,
    \sw_118_module_data_out[0] }));
 scanchain scanchain_119 (.clk_in(sw_118_clk_out),
    .clk_out(sw_119_clk_out),
    .data_in(sw_118_data_out),
    .data_out(sw_119_data_out),
    .latch_enable_in(sw_118_latch_out),
    .latch_enable_out(sw_119_latch_out),
    .scan_select_in(sw_118_scan_out),
    .scan_select_out(sw_119_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_119_module_data_in[7] ,
    \sw_119_module_data_in[6] ,
    \sw_119_module_data_in[5] ,
    \sw_119_module_data_in[4] ,
    \sw_119_module_data_in[3] ,
    \sw_119_module_data_in[2] ,
    \sw_119_module_data_in[1] ,
    \sw_119_module_data_in[0] }),
    .module_data_out({\sw_119_module_data_out[7] ,
    \sw_119_module_data_out[6] ,
    \sw_119_module_data_out[5] ,
    \sw_119_module_data_out[4] ,
    \sw_119_module_data_out[3] ,
    \sw_119_module_data_out[2] ,
    \sw_119_module_data_out[1] ,
    \sw_119_module_data_out[0] }));
 scanchain scanchain_12 (.clk_in(sw_011_clk_out),
    .clk_out(sw_012_clk_out),
    .data_in(sw_011_data_out),
    .data_out(sw_012_data_out),
    .latch_enable_in(sw_011_latch_out),
    .latch_enable_out(sw_012_latch_out),
    .scan_select_in(sw_011_scan_out),
    .scan_select_out(sw_012_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_012_module_data_in[7] ,
    \sw_012_module_data_in[6] ,
    \sw_012_module_data_in[5] ,
    \sw_012_module_data_in[4] ,
    \sw_012_module_data_in[3] ,
    \sw_012_module_data_in[2] ,
    \sw_012_module_data_in[1] ,
    \sw_012_module_data_in[0] }),
    .module_data_out({\sw_012_module_data_out[7] ,
    \sw_012_module_data_out[6] ,
    \sw_012_module_data_out[5] ,
    \sw_012_module_data_out[4] ,
    \sw_012_module_data_out[3] ,
    \sw_012_module_data_out[2] ,
    \sw_012_module_data_out[1] ,
    \sw_012_module_data_out[0] }));
 scanchain scanchain_120 (.clk_in(sw_119_clk_out),
    .clk_out(sw_120_clk_out),
    .data_in(sw_119_data_out),
    .data_out(sw_120_data_out),
    .latch_enable_in(sw_119_latch_out),
    .latch_enable_out(sw_120_latch_out),
    .scan_select_in(sw_119_scan_out),
    .scan_select_out(sw_120_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_120_module_data_in[7] ,
    \sw_120_module_data_in[6] ,
    \sw_120_module_data_in[5] ,
    \sw_120_module_data_in[4] ,
    \sw_120_module_data_in[3] ,
    \sw_120_module_data_in[2] ,
    \sw_120_module_data_in[1] ,
    \sw_120_module_data_in[0] }),
    .module_data_out({\sw_120_module_data_out[7] ,
    \sw_120_module_data_out[6] ,
    \sw_120_module_data_out[5] ,
    \sw_120_module_data_out[4] ,
    \sw_120_module_data_out[3] ,
    \sw_120_module_data_out[2] ,
    \sw_120_module_data_out[1] ,
    \sw_120_module_data_out[0] }));
 scanchain scanchain_121 (.clk_in(sw_120_clk_out),
    .clk_out(sw_121_clk_out),
    .data_in(sw_120_data_out),
    .data_out(sw_121_data_out),
    .latch_enable_in(sw_120_latch_out),
    .latch_enable_out(sw_121_latch_out),
    .scan_select_in(sw_120_scan_out),
    .scan_select_out(sw_121_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_121_module_data_in[7] ,
    \sw_121_module_data_in[6] ,
    \sw_121_module_data_in[5] ,
    \sw_121_module_data_in[4] ,
    \sw_121_module_data_in[3] ,
    \sw_121_module_data_in[2] ,
    \sw_121_module_data_in[1] ,
    \sw_121_module_data_in[0] }),
    .module_data_out({\sw_121_module_data_out[7] ,
    \sw_121_module_data_out[6] ,
    \sw_121_module_data_out[5] ,
    \sw_121_module_data_out[4] ,
    \sw_121_module_data_out[3] ,
    \sw_121_module_data_out[2] ,
    \sw_121_module_data_out[1] ,
    \sw_121_module_data_out[0] }));
 scanchain scanchain_122 (.clk_in(sw_121_clk_out),
    .clk_out(sw_122_clk_out),
    .data_in(sw_121_data_out),
    .data_out(sw_122_data_out),
    .latch_enable_in(sw_121_latch_out),
    .latch_enable_out(sw_122_latch_out),
    .scan_select_in(sw_121_scan_out),
    .scan_select_out(sw_122_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_122_module_data_in[7] ,
    \sw_122_module_data_in[6] ,
    \sw_122_module_data_in[5] ,
    \sw_122_module_data_in[4] ,
    \sw_122_module_data_in[3] ,
    \sw_122_module_data_in[2] ,
    \sw_122_module_data_in[1] ,
    \sw_122_module_data_in[0] }),
    .module_data_out({\sw_122_module_data_out[7] ,
    \sw_122_module_data_out[6] ,
    \sw_122_module_data_out[5] ,
    \sw_122_module_data_out[4] ,
    \sw_122_module_data_out[3] ,
    \sw_122_module_data_out[2] ,
    \sw_122_module_data_out[1] ,
    \sw_122_module_data_out[0] }));
 scanchain scanchain_123 (.clk_in(sw_122_clk_out),
    .clk_out(sw_123_clk_out),
    .data_in(sw_122_data_out),
    .data_out(sw_123_data_out),
    .latch_enable_in(sw_122_latch_out),
    .latch_enable_out(sw_123_latch_out),
    .scan_select_in(sw_122_scan_out),
    .scan_select_out(sw_123_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_123_module_data_in[7] ,
    \sw_123_module_data_in[6] ,
    \sw_123_module_data_in[5] ,
    \sw_123_module_data_in[4] ,
    \sw_123_module_data_in[3] ,
    \sw_123_module_data_in[2] ,
    \sw_123_module_data_in[1] ,
    \sw_123_module_data_in[0] }),
    .module_data_out({\sw_123_module_data_out[7] ,
    \sw_123_module_data_out[6] ,
    \sw_123_module_data_out[5] ,
    \sw_123_module_data_out[4] ,
    \sw_123_module_data_out[3] ,
    \sw_123_module_data_out[2] ,
    \sw_123_module_data_out[1] ,
    \sw_123_module_data_out[0] }));
 scanchain scanchain_124 (.clk_in(sw_123_clk_out),
    .clk_out(sw_124_clk_out),
    .data_in(sw_123_data_out),
    .data_out(sw_124_data_out),
    .latch_enable_in(sw_123_latch_out),
    .latch_enable_out(sw_124_latch_out),
    .scan_select_in(sw_123_scan_out),
    .scan_select_out(sw_124_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_124_module_data_in[7] ,
    \sw_124_module_data_in[6] ,
    \sw_124_module_data_in[5] ,
    \sw_124_module_data_in[4] ,
    \sw_124_module_data_in[3] ,
    \sw_124_module_data_in[2] ,
    \sw_124_module_data_in[1] ,
    \sw_124_module_data_in[0] }),
    .module_data_out({\sw_124_module_data_out[7] ,
    \sw_124_module_data_out[6] ,
    \sw_124_module_data_out[5] ,
    \sw_124_module_data_out[4] ,
    \sw_124_module_data_out[3] ,
    \sw_124_module_data_out[2] ,
    \sw_124_module_data_out[1] ,
    \sw_124_module_data_out[0] }));
 scanchain scanchain_125 (.clk_in(sw_124_clk_out),
    .clk_out(sw_125_clk_out),
    .data_in(sw_124_data_out),
    .data_out(sw_125_data_out),
    .latch_enable_in(sw_124_latch_out),
    .latch_enable_out(sw_125_latch_out),
    .scan_select_in(sw_124_scan_out),
    .scan_select_out(sw_125_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_125_module_data_in[7] ,
    \sw_125_module_data_in[6] ,
    \sw_125_module_data_in[5] ,
    \sw_125_module_data_in[4] ,
    \sw_125_module_data_in[3] ,
    \sw_125_module_data_in[2] ,
    \sw_125_module_data_in[1] ,
    \sw_125_module_data_in[0] }),
    .module_data_out({\sw_125_module_data_out[7] ,
    \sw_125_module_data_out[6] ,
    \sw_125_module_data_out[5] ,
    \sw_125_module_data_out[4] ,
    \sw_125_module_data_out[3] ,
    \sw_125_module_data_out[2] ,
    \sw_125_module_data_out[1] ,
    \sw_125_module_data_out[0] }));
 scanchain scanchain_126 (.clk_in(sw_125_clk_out),
    .clk_out(sw_126_clk_out),
    .data_in(sw_125_data_out),
    .data_out(sw_126_data_out),
    .latch_enable_in(sw_125_latch_out),
    .latch_enable_out(sw_126_latch_out),
    .scan_select_in(sw_125_scan_out),
    .scan_select_out(sw_126_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_126_module_data_in[7] ,
    \sw_126_module_data_in[6] ,
    \sw_126_module_data_in[5] ,
    \sw_126_module_data_in[4] ,
    \sw_126_module_data_in[3] ,
    \sw_126_module_data_in[2] ,
    \sw_126_module_data_in[1] ,
    \sw_126_module_data_in[0] }),
    .module_data_out({\sw_126_module_data_out[7] ,
    \sw_126_module_data_out[6] ,
    \sw_126_module_data_out[5] ,
    \sw_126_module_data_out[4] ,
    \sw_126_module_data_out[3] ,
    \sw_126_module_data_out[2] ,
    \sw_126_module_data_out[1] ,
    \sw_126_module_data_out[0] }));
 scanchain scanchain_127 (.clk_in(sw_126_clk_out),
    .clk_out(sw_127_clk_out),
    .data_in(sw_126_data_out),
    .data_out(sw_127_data_out),
    .latch_enable_in(sw_126_latch_out),
    .latch_enable_out(sw_127_latch_out),
    .scan_select_in(sw_126_scan_out),
    .scan_select_out(sw_127_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_127_module_data_in[7] ,
    \sw_127_module_data_in[6] ,
    \sw_127_module_data_in[5] ,
    \sw_127_module_data_in[4] ,
    \sw_127_module_data_in[3] ,
    \sw_127_module_data_in[2] ,
    \sw_127_module_data_in[1] ,
    \sw_127_module_data_in[0] }),
    .module_data_out({\sw_127_module_data_out[7] ,
    \sw_127_module_data_out[6] ,
    \sw_127_module_data_out[5] ,
    \sw_127_module_data_out[4] ,
    \sw_127_module_data_out[3] ,
    \sw_127_module_data_out[2] ,
    \sw_127_module_data_out[1] ,
    \sw_127_module_data_out[0] }));
 scanchain scanchain_128 (.clk_in(sw_127_clk_out),
    .clk_out(sw_128_clk_out),
    .data_in(sw_127_data_out),
    .data_out(sw_128_data_out),
    .latch_enable_in(sw_127_latch_out),
    .latch_enable_out(sw_128_latch_out),
    .scan_select_in(sw_127_scan_out),
    .scan_select_out(sw_128_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_128_module_data_in[7] ,
    \sw_128_module_data_in[6] ,
    \sw_128_module_data_in[5] ,
    \sw_128_module_data_in[4] ,
    \sw_128_module_data_in[3] ,
    \sw_128_module_data_in[2] ,
    \sw_128_module_data_in[1] ,
    \sw_128_module_data_in[0] }),
    .module_data_out({\sw_128_module_data_out[7] ,
    \sw_128_module_data_out[6] ,
    \sw_128_module_data_out[5] ,
    \sw_128_module_data_out[4] ,
    \sw_128_module_data_out[3] ,
    \sw_128_module_data_out[2] ,
    \sw_128_module_data_out[1] ,
    \sw_128_module_data_out[0] }));
 scanchain scanchain_129 (.clk_in(sw_128_clk_out),
    .clk_out(sw_129_clk_out),
    .data_in(sw_128_data_out),
    .data_out(sw_129_data_out),
    .latch_enable_in(sw_128_latch_out),
    .latch_enable_out(sw_129_latch_out),
    .scan_select_in(sw_128_scan_out),
    .scan_select_out(sw_129_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_129_module_data_in[7] ,
    \sw_129_module_data_in[6] ,
    \sw_129_module_data_in[5] ,
    \sw_129_module_data_in[4] ,
    \sw_129_module_data_in[3] ,
    \sw_129_module_data_in[2] ,
    \sw_129_module_data_in[1] ,
    \sw_129_module_data_in[0] }),
    .module_data_out({\sw_129_module_data_out[7] ,
    \sw_129_module_data_out[6] ,
    \sw_129_module_data_out[5] ,
    \sw_129_module_data_out[4] ,
    \sw_129_module_data_out[3] ,
    \sw_129_module_data_out[2] ,
    \sw_129_module_data_out[1] ,
    \sw_129_module_data_out[0] }));
 scanchain scanchain_13 (.clk_in(sw_012_clk_out),
    .clk_out(sw_013_clk_out),
    .data_in(sw_012_data_out),
    .data_out(sw_013_data_out),
    .latch_enable_in(sw_012_latch_out),
    .latch_enable_out(sw_013_latch_out),
    .scan_select_in(sw_012_scan_out),
    .scan_select_out(sw_013_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_013_module_data_in[7] ,
    \sw_013_module_data_in[6] ,
    \sw_013_module_data_in[5] ,
    \sw_013_module_data_in[4] ,
    \sw_013_module_data_in[3] ,
    \sw_013_module_data_in[2] ,
    \sw_013_module_data_in[1] ,
    \sw_013_module_data_in[0] }),
    .module_data_out({\sw_013_module_data_out[7] ,
    \sw_013_module_data_out[6] ,
    \sw_013_module_data_out[5] ,
    \sw_013_module_data_out[4] ,
    \sw_013_module_data_out[3] ,
    \sw_013_module_data_out[2] ,
    \sw_013_module_data_out[1] ,
    \sw_013_module_data_out[0] }));
 scanchain scanchain_130 (.clk_in(sw_129_clk_out),
    .clk_out(sw_130_clk_out),
    .data_in(sw_129_data_out),
    .data_out(sw_130_data_out),
    .latch_enable_in(sw_129_latch_out),
    .latch_enable_out(sw_130_latch_out),
    .scan_select_in(sw_129_scan_out),
    .scan_select_out(sw_130_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_130_module_data_in[7] ,
    \sw_130_module_data_in[6] ,
    \sw_130_module_data_in[5] ,
    \sw_130_module_data_in[4] ,
    \sw_130_module_data_in[3] ,
    \sw_130_module_data_in[2] ,
    \sw_130_module_data_in[1] ,
    \sw_130_module_data_in[0] }),
    .module_data_out({\sw_130_module_data_out[7] ,
    \sw_130_module_data_out[6] ,
    \sw_130_module_data_out[5] ,
    \sw_130_module_data_out[4] ,
    \sw_130_module_data_out[3] ,
    \sw_130_module_data_out[2] ,
    \sw_130_module_data_out[1] ,
    \sw_130_module_data_out[0] }));
 scanchain scanchain_131 (.clk_in(sw_130_clk_out),
    .clk_out(sw_131_clk_out),
    .data_in(sw_130_data_out),
    .data_out(sw_131_data_out),
    .latch_enable_in(sw_130_latch_out),
    .latch_enable_out(sw_131_latch_out),
    .scan_select_in(sw_130_scan_out),
    .scan_select_out(sw_131_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_131_module_data_in[7] ,
    \sw_131_module_data_in[6] ,
    \sw_131_module_data_in[5] ,
    \sw_131_module_data_in[4] ,
    \sw_131_module_data_in[3] ,
    \sw_131_module_data_in[2] ,
    \sw_131_module_data_in[1] ,
    \sw_131_module_data_in[0] }),
    .module_data_out({\sw_131_module_data_out[7] ,
    \sw_131_module_data_out[6] ,
    \sw_131_module_data_out[5] ,
    \sw_131_module_data_out[4] ,
    \sw_131_module_data_out[3] ,
    \sw_131_module_data_out[2] ,
    \sw_131_module_data_out[1] ,
    \sw_131_module_data_out[0] }));
 scanchain scanchain_132 (.clk_in(sw_131_clk_out),
    .clk_out(sw_132_clk_out),
    .data_in(sw_131_data_out),
    .data_out(sw_132_data_out),
    .latch_enable_in(sw_131_latch_out),
    .latch_enable_out(sw_132_latch_out),
    .scan_select_in(sw_131_scan_out),
    .scan_select_out(sw_132_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_132_module_data_in[7] ,
    \sw_132_module_data_in[6] ,
    \sw_132_module_data_in[5] ,
    \sw_132_module_data_in[4] ,
    \sw_132_module_data_in[3] ,
    \sw_132_module_data_in[2] ,
    \sw_132_module_data_in[1] ,
    \sw_132_module_data_in[0] }),
    .module_data_out({\sw_132_module_data_out[7] ,
    \sw_132_module_data_out[6] ,
    \sw_132_module_data_out[5] ,
    \sw_132_module_data_out[4] ,
    \sw_132_module_data_out[3] ,
    \sw_132_module_data_out[2] ,
    \sw_132_module_data_out[1] ,
    \sw_132_module_data_out[0] }));
 scanchain scanchain_133 (.clk_in(sw_132_clk_out),
    .clk_out(sw_133_clk_out),
    .data_in(sw_132_data_out),
    .data_out(sw_133_data_out),
    .latch_enable_in(sw_132_latch_out),
    .latch_enable_out(sw_133_latch_out),
    .scan_select_in(sw_132_scan_out),
    .scan_select_out(sw_133_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_133_module_data_in[7] ,
    \sw_133_module_data_in[6] ,
    \sw_133_module_data_in[5] ,
    \sw_133_module_data_in[4] ,
    \sw_133_module_data_in[3] ,
    \sw_133_module_data_in[2] ,
    \sw_133_module_data_in[1] ,
    \sw_133_module_data_in[0] }),
    .module_data_out({\sw_133_module_data_out[7] ,
    \sw_133_module_data_out[6] ,
    \sw_133_module_data_out[5] ,
    \sw_133_module_data_out[4] ,
    \sw_133_module_data_out[3] ,
    \sw_133_module_data_out[2] ,
    \sw_133_module_data_out[1] ,
    \sw_133_module_data_out[0] }));
 scanchain scanchain_134 (.clk_in(sw_133_clk_out),
    .clk_out(sw_134_clk_out),
    .data_in(sw_133_data_out),
    .data_out(sw_134_data_out),
    .latch_enable_in(sw_133_latch_out),
    .latch_enable_out(sw_134_latch_out),
    .scan_select_in(sw_133_scan_out),
    .scan_select_out(sw_134_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_134_module_data_in[7] ,
    \sw_134_module_data_in[6] ,
    \sw_134_module_data_in[5] ,
    \sw_134_module_data_in[4] ,
    \sw_134_module_data_in[3] ,
    \sw_134_module_data_in[2] ,
    \sw_134_module_data_in[1] ,
    \sw_134_module_data_in[0] }),
    .module_data_out({\sw_134_module_data_out[7] ,
    \sw_134_module_data_out[6] ,
    \sw_134_module_data_out[5] ,
    \sw_134_module_data_out[4] ,
    \sw_134_module_data_out[3] ,
    \sw_134_module_data_out[2] ,
    \sw_134_module_data_out[1] ,
    \sw_134_module_data_out[0] }));
 scanchain scanchain_135 (.clk_in(sw_134_clk_out),
    .clk_out(sw_135_clk_out),
    .data_in(sw_134_data_out),
    .data_out(sw_135_data_out),
    .latch_enable_in(sw_134_latch_out),
    .latch_enable_out(sw_135_latch_out),
    .scan_select_in(sw_134_scan_out),
    .scan_select_out(sw_135_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_135_module_data_in[7] ,
    \sw_135_module_data_in[6] ,
    \sw_135_module_data_in[5] ,
    \sw_135_module_data_in[4] ,
    \sw_135_module_data_in[3] ,
    \sw_135_module_data_in[2] ,
    \sw_135_module_data_in[1] ,
    \sw_135_module_data_in[0] }),
    .module_data_out({\sw_135_module_data_out[7] ,
    \sw_135_module_data_out[6] ,
    \sw_135_module_data_out[5] ,
    \sw_135_module_data_out[4] ,
    \sw_135_module_data_out[3] ,
    \sw_135_module_data_out[2] ,
    \sw_135_module_data_out[1] ,
    \sw_135_module_data_out[0] }));
 scanchain scanchain_136 (.clk_in(sw_135_clk_out),
    .clk_out(sw_136_clk_out),
    .data_in(sw_135_data_out),
    .data_out(sw_136_data_out),
    .latch_enable_in(sw_135_latch_out),
    .latch_enable_out(sw_136_latch_out),
    .scan_select_in(sw_135_scan_out),
    .scan_select_out(sw_136_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_136_module_data_in[7] ,
    \sw_136_module_data_in[6] ,
    \sw_136_module_data_in[5] ,
    \sw_136_module_data_in[4] ,
    \sw_136_module_data_in[3] ,
    \sw_136_module_data_in[2] ,
    \sw_136_module_data_in[1] ,
    \sw_136_module_data_in[0] }),
    .module_data_out({\sw_136_module_data_out[7] ,
    \sw_136_module_data_out[6] ,
    \sw_136_module_data_out[5] ,
    \sw_136_module_data_out[4] ,
    \sw_136_module_data_out[3] ,
    \sw_136_module_data_out[2] ,
    \sw_136_module_data_out[1] ,
    \sw_136_module_data_out[0] }));
 scanchain scanchain_137 (.clk_in(sw_136_clk_out),
    .clk_out(sw_137_clk_out),
    .data_in(sw_136_data_out),
    .data_out(sw_137_data_out),
    .latch_enable_in(sw_136_latch_out),
    .latch_enable_out(sw_137_latch_out),
    .scan_select_in(sw_136_scan_out),
    .scan_select_out(sw_137_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_137_module_data_in[7] ,
    \sw_137_module_data_in[6] ,
    \sw_137_module_data_in[5] ,
    \sw_137_module_data_in[4] ,
    \sw_137_module_data_in[3] ,
    \sw_137_module_data_in[2] ,
    \sw_137_module_data_in[1] ,
    \sw_137_module_data_in[0] }),
    .module_data_out({\sw_137_module_data_out[7] ,
    \sw_137_module_data_out[6] ,
    \sw_137_module_data_out[5] ,
    \sw_137_module_data_out[4] ,
    \sw_137_module_data_out[3] ,
    \sw_137_module_data_out[2] ,
    \sw_137_module_data_out[1] ,
    \sw_137_module_data_out[0] }));
 scanchain scanchain_138 (.clk_in(sw_137_clk_out),
    .clk_out(sw_138_clk_out),
    .data_in(sw_137_data_out),
    .data_out(sw_138_data_out),
    .latch_enable_in(sw_137_latch_out),
    .latch_enable_out(sw_138_latch_out),
    .scan_select_in(sw_137_scan_out),
    .scan_select_out(sw_138_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_138_module_data_in[7] ,
    \sw_138_module_data_in[6] ,
    \sw_138_module_data_in[5] ,
    \sw_138_module_data_in[4] ,
    \sw_138_module_data_in[3] ,
    \sw_138_module_data_in[2] ,
    \sw_138_module_data_in[1] ,
    \sw_138_module_data_in[0] }),
    .module_data_out({\sw_138_module_data_out[7] ,
    \sw_138_module_data_out[6] ,
    \sw_138_module_data_out[5] ,
    \sw_138_module_data_out[4] ,
    \sw_138_module_data_out[3] ,
    \sw_138_module_data_out[2] ,
    \sw_138_module_data_out[1] ,
    \sw_138_module_data_out[0] }));
 scanchain scanchain_139 (.clk_in(sw_138_clk_out),
    .clk_out(sw_139_clk_out),
    .data_in(sw_138_data_out),
    .data_out(sw_139_data_out),
    .latch_enable_in(sw_138_latch_out),
    .latch_enable_out(sw_139_latch_out),
    .scan_select_in(sw_138_scan_out),
    .scan_select_out(sw_139_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_139_module_data_in[7] ,
    \sw_139_module_data_in[6] ,
    \sw_139_module_data_in[5] ,
    \sw_139_module_data_in[4] ,
    \sw_139_module_data_in[3] ,
    \sw_139_module_data_in[2] ,
    \sw_139_module_data_in[1] ,
    \sw_139_module_data_in[0] }),
    .module_data_out({\sw_139_module_data_out[7] ,
    \sw_139_module_data_out[6] ,
    \sw_139_module_data_out[5] ,
    \sw_139_module_data_out[4] ,
    \sw_139_module_data_out[3] ,
    \sw_139_module_data_out[2] ,
    \sw_139_module_data_out[1] ,
    \sw_139_module_data_out[0] }));
 scanchain scanchain_14 (.clk_in(sw_013_clk_out),
    .clk_out(sw_014_clk_out),
    .data_in(sw_013_data_out),
    .data_out(sw_014_data_out),
    .latch_enable_in(sw_013_latch_out),
    .latch_enable_out(sw_014_latch_out),
    .scan_select_in(sw_013_scan_out),
    .scan_select_out(sw_014_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_014_module_data_in[7] ,
    \sw_014_module_data_in[6] ,
    \sw_014_module_data_in[5] ,
    \sw_014_module_data_in[4] ,
    \sw_014_module_data_in[3] ,
    \sw_014_module_data_in[2] ,
    \sw_014_module_data_in[1] ,
    \sw_014_module_data_in[0] }),
    .module_data_out({\sw_014_module_data_out[7] ,
    \sw_014_module_data_out[6] ,
    \sw_014_module_data_out[5] ,
    \sw_014_module_data_out[4] ,
    \sw_014_module_data_out[3] ,
    \sw_014_module_data_out[2] ,
    \sw_014_module_data_out[1] ,
    \sw_014_module_data_out[0] }));
 scanchain scanchain_140 (.clk_in(sw_139_clk_out),
    .clk_out(sw_140_clk_out),
    .data_in(sw_139_data_out),
    .data_out(sw_140_data_out),
    .latch_enable_in(sw_139_latch_out),
    .latch_enable_out(sw_140_latch_out),
    .scan_select_in(sw_139_scan_out),
    .scan_select_out(sw_140_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_140_module_data_in[7] ,
    \sw_140_module_data_in[6] ,
    \sw_140_module_data_in[5] ,
    \sw_140_module_data_in[4] ,
    \sw_140_module_data_in[3] ,
    \sw_140_module_data_in[2] ,
    \sw_140_module_data_in[1] ,
    \sw_140_module_data_in[0] }),
    .module_data_out({\sw_140_module_data_out[7] ,
    \sw_140_module_data_out[6] ,
    \sw_140_module_data_out[5] ,
    \sw_140_module_data_out[4] ,
    \sw_140_module_data_out[3] ,
    \sw_140_module_data_out[2] ,
    \sw_140_module_data_out[1] ,
    \sw_140_module_data_out[0] }));
 scanchain scanchain_141 (.clk_in(sw_140_clk_out),
    .clk_out(sw_141_clk_out),
    .data_in(sw_140_data_out),
    .data_out(sw_141_data_out),
    .latch_enable_in(sw_140_latch_out),
    .latch_enable_out(sw_141_latch_out),
    .scan_select_in(sw_140_scan_out),
    .scan_select_out(sw_141_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_141_module_data_in[7] ,
    \sw_141_module_data_in[6] ,
    \sw_141_module_data_in[5] ,
    \sw_141_module_data_in[4] ,
    \sw_141_module_data_in[3] ,
    \sw_141_module_data_in[2] ,
    \sw_141_module_data_in[1] ,
    \sw_141_module_data_in[0] }),
    .module_data_out({\sw_141_module_data_out[7] ,
    \sw_141_module_data_out[6] ,
    \sw_141_module_data_out[5] ,
    \sw_141_module_data_out[4] ,
    \sw_141_module_data_out[3] ,
    \sw_141_module_data_out[2] ,
    \sw_141_module_data_out[1] ,
    \sw_141_module_data_out[0] }));
 scanchain scanchain_142 (.clk_in(sw_141_clk_out),
    .clk_out(sw_142_clk_out),
    .data_in(sw_141_data_out),
    .data_out(sw_142_data_out),
    .latch_enable_in(sw_141_latch_out),
    .latch_enable_out(sw_142_latch_out),
    .scan_select_in(sw_141_scan_out),
    .scan_select_out(sw_142_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_142_module_data_in[7] ,
    \sw_142_module_data_in[6] ,
    \sw_142_module_data_in[5] ,
    \sw_142_module_data_in[4] ,
    \sw_142_module_data_in[3] ,
    \sw_142_module_data_in[2] ,
    \sw_142_module_data_in[1] ,
    \sw_142_module_data_in[0] }),
    .module_data_out({\sw_142_module_data_out[7] ,
    \sw_142_module_data_out[6] ,
    \sw_142_module_data_out[5] ,
    \sw_142_module_data_out[4] ,
    \sw_142_module_data_out[3] ,
    \sw_142_module_data_out[2] ,
    \sw_142_module_data_out[1] ,
    \sw_142_module_data_out[0] }));
 scanchain scanchain_143 (.clk_in(sw_142_clk_out),
    .clk_out(sw_143_clk_out),
    .data_in(sw_142_data_out),
    .data_out(sw_143_data_out),
    .latch_enable_in(sw_142_latch_out),
    .latch_enable_out(sw_143_latch_out),
    .scan_select_in(sw_142_scan_out),
    .scan_select_out(sw_143_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_143_module_data_in[7] ,
    \sw_143_module_data_in[6] ,
    \sw_143_module_data_in[5] ,
    \sw_143_module_data_in[4] ,
    \sw_143_module_data_in[3] ,
    \sw_143_module_data_in[2] ,
    \sw_143_module_data_in[1] ,
    \sw_143_module_data_in[0] }),
    .module_data_out({\sw_143_module_data_out[7] ,
    \sw_143_module_data_out[6] ,
    \sw_143_module_data_out[5] ,
    \sw_143_module_data_out[4] ,
    \sw_143_module_data_out[3] ,
    \sw_143_module_data_out[2] ,
    \sw_143_module_data_out[1] ,
    \sw_143_module_data_out[0] }));
 scanchain scanchain_144 (.clk_in(sw_143_clk_out),
    .clk_out(sw_144_clk_out),
    .data_in(sw_143_data_out),
    .data_out(sw_144_data_out),
    .latch_enable_in(sw_143_latch_out),
    .latch_enable_out(sw_144_latch_out),
    .scan_select_in(sw_143_scan_out),
    .scan_select_out(sw_144_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_144_module_data_in[7] ,
    \sw_144_module_data_in[6] ,
    \sw_144_module_data_in[5] ,
    \sw_144_module_data_in[4] ,
    \sw_144_module_data_in[3] ,
    \sw_144_module_data_in[2] ,
    \sw_144_module_data_in[1] ,
    \sw_144_module_data_in[0] }),
    .module_data_out({\sw_144_module_data_out[7] ,
    \sw_144_module_data_out[6] ,
    \sw_144_module_data_out[5] ,
    \sw_144_module_data_out[4] ,
    \sw_144_module_data_out[3] ,
    \sw_144_module_data_out[2] ,
    \sw_144_module_data_out[1] ,
    \sw_144_module_data_out[0] }));
 scanchain scanchain_145 (.clk_in(sw_144_clk_out),
    .clk_out(sw_145_clk_out),
    .data_in(sw_144_data_out),
    .data_out(sw_145_data_out),
    .latch_enable_in(sw_144_latch_out),
    .latch_enable_out(sw_145_latch_out),
    .scan_select_in(sw_144_scan_out),
    .scan_select_out(sw_145_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_145_module_data_in[7] ,
    \sw_145_module_data_in[6] ,
    \sw_145_module_data_in[5] ,
    \sw_145_module_data_in[4] ,
    \sw_145_module_data_in[3] ,
    \sw_145_module_data_in[2] ,
    \sw_145_module_data_in[1] ,
    \sw_145_module_data_in[0] }),
    .module_data_out({\sw_145_module_data_out[7] ,
    \sw_145_module_data_out[6] ,
    \sw_145_module_data_out[5] ,
    \sw_145_module_data_out[4] ,
    \sw_145_module_data_out[3] ,
    \sw_145_module_data_out[2] ,
    \sw_145_module_data_out[1] ,
    \sw_145_module_data_out[0] }));
 scanchain scanchain_146 (.clk_in(sw_145_clk_out),
    .clk_out(sw_146_clk_out),
    .data_in(sw_145_data_out),
    .data_out(sw_146_data_out),
    .latch_enable_in(sw_145_latch_out),
    .latch_enable_out(sw_146_latch_out),
    .scan_select_in(sw_145_scan_out),
    .scan_select_out(sw_146_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_146_module_data_in[7] ,
    \sw_146_module_data_in[6] ,
    \sw_146_module_data_in[5] ,
    \sw_146_module_data_in[4] ,
    \sw_146_module_data_in[3] ,
    \sw_146_module_data_in[2] ,
    \sw_146_module_data_in[1] ,
    \sw_146_module_data_in[0] }),
    .module_data_out({\sw_146_module_data_out[7] ,
    \sw_146_module_data_out[6] ,
    \sw_146_module_data_out[5] ,
    \sw_146_module_data_out[4] ,
    \sw_146_module_data_out[3] ,
    \sw_146_module_data_out[2] ,
    \sw_146_module_data_out[1] ,
    \sw_146_module_data_out[0] }));
 scanchain scanchain_147 (.clk_in(sw_146_clk_out),
    .clk_out(sw_147_clk_out),
    .data_in(sw_146_data_out),
    .data_out(sw_147_data_out),
    .latch_enable_in(sw_146_latch_out),
    .latch_enable_out(sw_147_latch_out),
    .scan_select_in(sw_146_scan_out),
    .scan_select_out(sw_147_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_147_module_data_in[7] ,
    \sw_147_module_data_in[6] ,
    \sw_147_module_data_in[5] ,
    \sw_147_module_data_in[4] ,
    \sw_147_module_data_in[3] ,
    \sw_147_module_data_in[2] ,
    \sw_147_module_data_in[1] ,
    \sw_147_module_data_in[0] }),
    .module_data_out({\sw_147_module_data_out[7] ,
    \sw_147_module_data_out[6] ,
    \sw_147_module_data_out[5] ,
    \sw_147_module_data_out[4] ,
    \sw_147_module_data_out[3] ,
    \sw_147_module_data_out[2] ,
    \sw_147_module_data_out[1] ,
    \sw_147_module_data_out[0] }));
 scanchain scanchain_148 (.clk_in(sw_147_clk_out),
    .clk_out(sw_148_clk_out),
    .data_in(sw_147_data_out),
    .data_out(sw_148_data_out),
    .latch_enable_in(sw_147_latch_out),
    .latch_enable_out(sw_148_latch_out),
    .scan_select_in(sw_147_scan_out),
    .scan_select_out(sw_148_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_148_module_data_in[7] ,
    \sw_148_module_data_in[6] ,
    \sw_148_module_data_in[5] ,
    \sw_148_module_data_in[4] ,
    \sw_148_module_data_in[3] ,
    \sw_148_module_data_in[2] ,
    \sw_148_module_data_in[1] ,
    \sw_148_module_data_in[0] }),
    .module_data_out({\sw_148_module_data_out[7] ,
    \sw_148_module_data_out[6] ,
    \sw_148_module_data_out[5] ,
    \sw_148_module_data_out[4] ,
    \sw_148_module_data_out[3] ,
    \sw_148_module_data_out[2] ,
    \sw_148_module_data_out[1] ,
    \sw_148_module_data_out[0] }));
 scanchain scanchain_149 (.clk_in(sw_148_clk_out),
    .clk_out(sw_149_clk_out),
    .data_in(sw_148_data_out),
    .data_out(sw_149_data_out),
    .latch_enable_in(sw_148_latch_out),
    .latch_enable_out(sw_149_latch_out),
    .scan_select_in(sw_148_scan_out),
    .scan_select_out(sw_149_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_149_module_data_in[7] ,
    \sw_149_module_data_in[6] ,
    \sw_149_module_data_in[5] ,
    \sw_149_module_data_in[4] ,
    \sw_149_module_data_in[3] ,
    \sw_149_module_data_in[2] ,
    \sw_149_module_data_in[1] ,
    \sw_149_module_data_in[0] }),
    .module_data_out({\sw_149_module_data_out[7] ,
    \sw_149_module_data_out[6] ,
    \sw_149_module_data_out[5] ,
    \sw_149_module_data_out[4] ,
    \sw_149_module_data_out[3] ,
    \sw_149_module_data_out[2] ,
    \sw_149_module_data_out[1] ,
    \sw_149_module_data_out[0] }));
 scanchain scanchain_15 (.clk_in(sw_014_clk_out),
    .clk_out(sw_015_clk_out),
    .data_in(sw_014_data_out),
    .data_out(sw_015_data_out),
    .latch_enable_in(sw_014_latch_out),
    .latch_enable_out(sw_015_latch_out),
    .scan_select_in(sw_014_scan_out),
    .scan_select_out(sw_015_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_015_module_data_in[7] ,
    \sw_015_module_data_in[6] ,
    \sw_015_module_data_in[5] ,
    \sw_015_module_data_in[4] ,
    \sw_015_module_data_in[3] ,
    \sw_015_module_data_in[2] ,
    \sw_015_module_data_in[1] ,
    \sw_015_module_data_in[0] }),
    .module_data_out({\sw_015_module_data_out[7] ,
    \sw_015_module_data_out[6] ,
    \sw_015_module_data_out[5] ,
    \sw_015_module_data_out[4] ,
    \sw_015_module_data_out[3] ,
    \sw_015_module_data_out[2] ,
    \sw_015_module_data_out[1] ,
    \sw_015_module_data_out[0] }));
 scanchain scanchain_150 (.clk_in(sw_149_clk_out),
    .clk_out(sw_150_clk_out),
    .data_in(sw_149_data_out),
    .data_out(sw_150_data_out),
    .latch_enable_in(sw_149_latch_out),
    .latch_enable_out(sw_150_latch_out),
    .scan_select_in(sw_149_scan_out),
    .scan_select_out(sw_150_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_150_module_data_in[7] ,
    \sw_150_module_data_in[6] ,
    \sw_150_module_data_in[5] ,
    \sw_150_module_data_in[4] ,
    \sw_150_module_data_in[3] ,
    \sw_150_module_data_in[2] ,
    \sw_150_module_data_in[1] ,
    \sw_150_module_data_in[0] }),
    .module_data_out({\sw_150_module_data_out[7] ,
    \sw_150_module_data_out[6] ,
    \sw_150_module_data_out[5] ,
    \sw_150_module_data_out[4] ,
    \sw_150_module_data_out[3] ,
    \sw_150_module_data_out[2] ,
    \sw_150_module_data_out[1] ,
    \sw_150_module_data_out[0] }));
 scanchain scanchain_151 (.clk_in(sw_150_clk_out),
    .clk_out(sw_151_clk_out),
    .data_in(sw_150_data_out),
    .data_out(sw_151_data_out),
    .latch_enable_in(sw_150_latch_out),
    .latch_enable_out(sw_151_latch_out),
    .scan_select_in(sw_150_scan_out),
    .scan_select_out(sw_151_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_151_module_data_in[7] ,
    \sw_151_module_data_in[6] ,
    \sw_151_module_data_in[5] ,
    \sw_151_module_data_in[4] ,
    \sw_151_module_data_in[3] ,
    \sw_151_module_data_in[2] ,
    \sw_151_module_data_in[1] ,
    \sw_151_module_data_in[0] }),
    .module_data_out({\sw_151_module_data_out[7] ,
    \sw_151_module_data_out[6] ,
    \sw_151_module_data_out[5] ,
    \sw_151_module_data_out[4] ,
    \sw_151_module_data_out[3] ,
    \sw_151_module_data_out[2] ,
    \sw_151_module_data_out[1] ,
    \sw_151_module_data_out[0] }));
 scanchain scanchain_152 (.clk_in(sw_151_clk_out),
    .clk_out(sw_152_clk_out),
    .data_in(sw_151_data_out),
    .data_out(sw_152_data_out),
    .latch_enable_in(sw_151_latch_out),
    .latch_enable_out(sw_152_latch_out),
    .scan_select_in(sw_151_scan_out),
    .scan_select_out(sw_152_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_152_module_data_in[7] ,
    \sw_152_module_data_in[6] ,
    \sw_152_module_data_in[5] ,
    \sw_152_module_data_in[4] ,
    \sw_152_module_data_in[3] ,
    \sw_152_module_data_in[2] ,
    \sw_152_module_data_in[1] ,
    \sw_152_module_data_in[0] }),
    .module_data_out({\sw_152_module_data_out[7] ,
    \sw_152_module_data_out[6] ,
    \sw_152_module_data_out[5] ,
    \sw_152_module_data_out[4] ,
    \sw_152_module_data_out[3] ,
    \sw_152_module_data_out[2] ,
    \sw_152_module_data_out[1] ,
    \sw_152_module_data_out[0] }));
 scanchain scanchain_153 (.clk_in(sw_152_clk_out),
    .clk_out(sw_153_clk_out),
    .data_in(sw_152_data_out),
    .data_out(sw_153_data_out),
    .latch_enable_in(sw_152_latch_out),
    .latch_enable_out(sw_153_latch_out),
    .scan_select_in(sw_152_scan_out),
    .scan_select_out(sw_153_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_153_module_data_in[7] ,
    \sw_153_module_data_in[6] ,
    \sw_153_module_data_in[5] ,
    \sw_153_module_data_in[4] ,
    \sw_153_module_data_in[3] ,
    \sw_153_module_data_in[2] ,
    \sw_153_module_data_in[1] ,
    \sw_153_module_data_in[0] }),
    .module_data_out({\sw_153_module_data_out[7] ,
    \sw_153_module_data_out[6] ,
    \sw_153_module_data_out[5] ,
    \sw_153_module_data_out[4] ,
    \sw_153_module_data_out[3] ,
    \sw_153_module_data_out[2] ,
    \sw_153_module_data_out[1] ,
    \sw_153_module_data_out[0] }));
 scanchain scanchain_154 (.clk_in(sw_153_clk_out),
    .clk_out(sw_154_clk_out),
    .data_in(sw_153_data_out),
    .data_out(sw_154_data_out),
    .latch_enable_in(sw_153_latch_out),
    .latch_enable_out(sw_154_latch_out),
    .scan_select_in(sw_153_scan_out),
    .scan_select_out(sw_154_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_154_module_data_in[7] ,
    \sw_154_module_data_in[6] ,
    \sw_154_module_data_in[5] ,
    \sw_154_module_data_in[4] ,
    \sw_154_module_data_in[3] ,
    \sw_154_module_data_in[2] ,
    \sw_154_module_data_in[1] ,
    \sw_154_module_data_in[0] }),
    .module_data_out({\sw_154_module_data_out[7] ,
    \sw_154_module_data_out[6] ,
    \sw_154_module_data_out[5] ,
    \sw_154_module_data_out[4] ,
    \sw_154_module_data_out[3] ,
    \sw_154_module_data_out[2] ,
    \sw_154_module_data_out[1] ,
    \sw_154_module_data_out[0] }));
 scanchain scanchain_155 (.clk_in(sw_154_clk_out),
    .clk_out(sw_155_clk_out),
    .data_in(sw_154_data_out),
    .data_out(sw_155_data_out),
    .latch_enable_in(sw_154_latch_out),
    .latch_enable_out(sw_155_latch_out),
    .scan_select_in(sw_154_scan_out),
    .scan_select_out(sw_155_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_155_module_data_in[7] ,
    \sw_155_module_data_in[6] ,
    \sw_155_module_data_in[5] ,
    \sw_155_module_data_in[4] ,
    \sw_155_module_data_in[3] ,
    \sw_155_module_data_in[2] ,
    \sw_155_module_data_in[1] ,
    \sw_155_module_data_in[0] }),
    .module_data_out({\sw_155_module_data_out[7] ,
    \sw_155_module_data_out[6] ,
    \sw_155_module_data_out[5] ,
    \sw_155_module_data_out[4] ,
    \sw_155_module_data_out[3] ,
    \sw_155_module_data_out[2] ,
    \sw_155_module_data_out[1] ,
    \sw_155_module_data_out[0] }));
 scanchain scanchain_156 (.clk_in(sw_155_clk_out),
    .clk_out(sw_156_clk_out),
    .data_in(sw_155_data_out),
    .data_out(sw_156_data_out),
    .latch_enable_in(sw_155_latch_out),
    .latch_enable_out(sw_156_latch_out),
    .scan_select_in(sw_155_scan_out),
    .scan_select_out(sw_156_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_156_module_data_in[7] ,
    \sw_156_module_data_in[6] ,
    \sw_156_module_data_in[5] ,
    \sw_156_module_data_in[4] ,
    \sw_156_module_data_in[3] ,
    \sw_156_module_data_in[2] ,
    \sw_156_module_data_in[1] ,
    \sw_156_module_data_in[0] }),
    .module_data_out({\sw_156_module_data_out[7] ,
    \sw_156_module_data_out[6] ,
    \sw_156_module_data_out[5] ,
    \sw_156_module_data_out[4] ,
    \sw_156_module_data_out[3] ,
    \sw_156_module_data_out[2] ,
    \sw_156_module_data_out[1] ,
    \sw_156_module_data_out[0] }));
 scanchain scanchain_157 (.clk_in(sw_156_clk_out),
    .clk_out(sw_157_clk_out),
    .data_in(sw_156_data_out),
    .data_out(sw_157_data_out),
    .latch_enable_in(sw_156_latch_out),
    .latch_enable_out(sw_157_latch_out),
    .scan_select_in(sw_156_scan_out),
    .scan_select_out(sw_157_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_157_module_data_in[7] ,
    \sw_157_module_data_in[6] ,
    \sw_157_module_data_in[5] ,
    \sw_157_module_data_in[4] ,
    \sw_157_module_data_in[3] ,
    \sw_157_module_data_in[2] ,
    \sw_157_module_data_in[1] ,
    \sw_157_module_data_in[0] }),
    .module_data_out({\sw_157_module_data_out[7] ,
    \sw_157_module_data_out[6] ,
    \sw_157_module_data_out[5] ,
    \sw_157_module_data_out[4] ,
    \sw_157_module_data_out[3] ,
    \sw_157_module_data_out[2] ,
    \sw_157_module_data_out[1] ,
    \sw_157_module_data_out[0] }));
 scanchain scanchain_158 (.clk_in(sw_157_clk_out),
    .clk_out(sw_158_clk_out),
    .data_in(sw_157_data_out),
    .data_out(sw_158_data_out),
    .latch_enable_in(sw_157_latch_out),
    .latch_enable_out(sw_158_latch_out),
    .scan_select_in(sw_157_scan_out),
    .scan_select_out(sw_158_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_158_module_data_in[7] ,
    \sw_158_module_data_in[6] ,
    \sw_158_module_data_in[5] ,
    \sw_158_module_data_in[4] ,
    \sw_158_module_data_in[3] ,
    \sw_158_module_data_in[2] ,
    \sw_158_module_data_in[1] ,
    \sw_158_module_data_in[0] }),
    .module_data_out({\sw_158_module_data_out[7] ,
    \sw_158_module_data_out[6] ,
    \sw_158_module_data_out[5] ,
    \sw_158_module_data_out[4] ,
    \sw_158_module_data_out[3] ,
    \sw_158_module_data_out[2] ,
    \sw_158_module_data_out[1] ,
    \sw_158_module_data_out[0] }));
 scanchain scanchain_159 (.clk_in(sw_158_clk_out),
    .clk_out(sw_159_clk_out),
    .data_in(sw_158_data_out),
    .data_out(sw_159_data_out),
    .latch_enable_in(sw_158_latch_out),
    .latch_enable_out(sw_159_latch_out),
    .scan_select_in(sw_158_scan_out),
    .scan_select_out(sw_159_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_159_module_data_in[7] ,
    \sw_159_module_data_in[6] ,
    \sw_159_module_data_in[5] ,
    \sw_159_module_data_in[4] ,
    \sw_159_module_data_in[3] ,
    \sw_159_module_data_in[2] ,
    \sw_159_module_data_in[1] ,
    \sw_159_module_data_in[0] }),
    .module_data_out({\sw_159_module_data_out[7] ,
    \sw_159_module_data_out[6] ,
    \sw_159_module_data_out[5] ,
    \sw_159_module_data_out[4] ,
    \sw_159_module_data_out[3] ,
    \sw_159_module_data_out[2] ,
    \sw_159_module_data_out[1] ,
    \sw_159_module_data_out[0] }));
 scanchain scanchain_16 (.clk_in(sw_015_clk_out),
    .clk_out(sw_016_clk_out),
    .data_in(sw_015_data_out),
    .data_out(sw_016_data_out),
    .latch_enable_in(sw_015_latch_out),
    .latch_enable_out(sw_016_latch_out),
    .scan_select_in(sw_015_scan_out),
    .scan_select_out(sw_016_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_016_module_data_in[7] ,
    \sw_016_module_data_in[6] ,
    \sw_016_module_data_in[5] ,
    \sw_016_module_data_in[4] ,
    \sw_016_module_data_in[3] ,
    \sw_016_module_data_in[2] ,
    \sw_016_module_data_in[1] ,
    \sw_016_module_data_in[0] }),
    .module_data_out({\sw_016_module_data_out[7] ,
    \sw_016_module_data_out[6] ,
    \sw_016_module_data_out[5] ,
    \sw_016_module_data_out[4] ,
    \sw_016_module_data_out[3] ,
    \sw_016_module_data_out[2] ,
    \sw_016_module_data_out[1] ,
    \sw_016_module_data_out[0] }));
 scanchain scanchain_160 (.clk_in(sw_159_clk_out),
    .clk_out(sw_160_clk_out),
    .data_in(sw_159_data_out),
    .data_out(sw_160_data_out),
    .latch_enable_in(sw_159_latch_out),
    .latch_enable_out(sw_160_latch_out),
    .scan_select_in(sw_159_scan_out),
    .scan_select_out(sw_160_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_160_module_data_in[7] ,
    \sw_160_module_data_in[6] ,
    \sw_160_module_data_in[5] ,
    \sw_160_module_data_in[4] ,
    \sw_160_module_data_in[3] ,
    \sw_160_module_data_in[2] ,
    \sw_160_module_data_in[1] ,
    \sw_160_module_data_in[0] }),
    .module_data_out({\sw_160_module_data_out[7] ,
    \sw_160_module_data_out[6] ,
    \sw_160_module_data_out[5] ,
    \sw_160_module_data_out[4] ,
    \sw_160_module_data_out[3] ,
    \sw_160_module_data_out[2] ,
    \sw_160_module_data_out[1] ,
    \sw_160_module_data_out[0] }));
 scanchain scanchain_161 (.clk_in(sw_160_clk_out),
    .clk_out(sw_161_clk_out),
    .data_in(sw_160_data_out),
    .data_out(sw_161_data_out),
    .latch_enable_in(sw_160_latch_out),
    .latch_enable_out(sw_161_latch_out),
    .scan_select_in(sw_160_scan_out),
    .scan_select_out(sw_161_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_161_module_data_in[7] ,
    \sw_161_module_data_in[6] ,
    \sw_161_module_data_in[5] ,
    \sw_161_module_data_in[4] ,
    \sw_161_module_data_in[3] ,
    \sw_161_module_data_in[2] ,
    \sw_161_module_data_in[1] ,
    \sw_161_module_data_in[0] }),
    .module_data_out({\sw_161_module_data_out[7] ,
    \sw_161_module_data_out[6] ,
    \sw_161_module_data_out[5] ,
    \sw_161_module_data_out[4] ,
    \sw_161_module_data_out[3] ,
    \sw_161_module_data_out[2] ,
    \sw_161_module_data_out[1] ,
    \sw_161_module_data_out[0] }));
 scanchain scanchain_162 (.clk_in(sw_161_clk_out),
    .clk_out(sw_162_clk_out),
    .data_in(sw_161_data_out),
    .data_out(sw_162_data_out),
    .latch_enable_in(sw_161_latch_out),
    .latch_enable_out(sw_162_latch_out),
    .scan_select_in(sw_161_scan_out),
    .scan_select_out(sw_162_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_162_module_data_in[7] ,
    \sw_162_module_data_in[6] ,
    \sw_162_module_data_in[5] ,
    \sw_162_module_data_in[4] ,
    \sw_162_module_data_in[3] ,
    \sw_162_module_data_in[2] ,
    \sw_162_module_data_in[1] ,
    \sw_162_module_data_in[0] }),
    .module_data_out({\sw_162_module_data_out[7] ,
    \sw_162_module_data_out[6] ,
    \sw_162_module_data_out[5] ,
    \sw_162_module_data_out[4] ,
    \sw_162_module_data_out[3] ,
    \sw_162_module_data_out[2] ,
    \sw_162_module_data_out[1] ,
    \sw_162_module_data_out[0] }));
 scanchain scanchain_163 (.clk_in(sw_162_clk_out),
    .clk_out(sw_163_clk_out),
    .data_in(sw_162_data_out),
    .data_out(sw_163_data_out),
    .latch_enable_in(sw_162_latch_out),
    .latch_enable_out(sw_163_latch_out),
    .scan_select_in(sw_162_scan_out),
    .scan_select_out(sw_163_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_163_module_data_in[7] ,
    \sw_163_module_data_in[6] ,
    \sw_163_module_data_in[5] ,
    \sw_163_module_data_in[4] ,
    \sw_163_module_data_in[3] ,
    \sw_163_module_data_in[2] ,
    \sw_163_module_data_in[1] ,
    \sw_163_module_data_in[0] }),
    .module_data_out({\sw_163_module_data_out[7] ,
    \sw_163_module_data_out[6] ,
    \sw_163_module_data_out[5] ,
    \sw_163_module_data_out[4] ,
    \sw_163_module_data_out[3] ,
    \sw_163_module_data_out[2] ,
    \sw_163_module_data_out[1] ,
    \sw_163_module_data_out[0] }));
 scanchain scanchain_164 (.clk_in(sw_163_clk_out),
    .clk_out(sw_164_clk_out),
    .data_in(sw_163_data_out),
    .data_out(sw_164_data_out),
    .latch_enable_in(sw_163_latch_out),
    .latch_enable_out(sw_164_latch_out),
    .scan_select_in(sw_163_scan_out),
    .scan_select_out(sw_164_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_164_module_data_in[7] ,
    \sw_164_module_data_in[6] ,
    \sw_164_module_data_in[5] ,
    \sw_164_module_data_in[4] ,
    \sw_164_module_data_in[3] ,
    \sw_164_module_data_in[2] ,
    \sw_164_module_data_in[1] ,
    \sw_164_module_data_in[0] }),
    .module_data_out({\sw_164_module_data_out[7] ,
    \sw_164_module_data_out[6] ,
    \sw_164_module_data_out[5] ,
    \sw_164_module_data_out[4] ,
    \sw_164_module_data_out[3] ,
    \sw_164_module_data_out[2] ,
    \sw_164_module_data_out[1] ,
    \sw_164_module_data_out[0] }));
 scanchain scanchain_165 (.clk_in(sw_164_clk_out),
    .clk_out(sw_165_clk_out),
    .data_in(sw_164_data_out),
    .data_out(sw_165_data_out),
    .latch_enable_in(sw_164_latch_out),
    .latch_enable_out(sw_165_latch_out),
    .scan_select_in(sw_164_scan_out),
    .scan_select_out(sw_165_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_165_module_data_in[7] ,
    \sw_165_module_data_in[6] ,
    \sw_165_module_data_in[5] ,
    \sw_165_module_data_in[4] ,
    \sw_165_module_data_in[3] ,
    \sw_165_module_data_in[2] ,
    \sw_165_module_data_in[1] ,
    \sw_165_module_data_in[0] }),
    .module_data_out({\sw_165_module_data_out[7] ,
    \sw_165_module_data_out[6] ,
    \sw_165_module_data_out[5] ,
    \sw_165_module_data_out[4] ,
    \sw_165_module_data_out[3] ,
    \sw_165_module_data_out[2] ,
    \sw_165_module_data_out[1] ,
    \sw_165_module_data_out[0] }));
 scanchain scanchain_166 (.clk_in(sw_165_clk_out),
    .clk_out(sw_166_clk_out),
    .data_in(sw_165_data_out),
    .data_out(sw_166_data_out),
    .latch_enable_in(sw_165_latch_out),
    .latch_enable_out(sw_166_latch_out),
    .scan_select_in(sw_165_scan_out),
    .scan_select_out(sw_166_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_166_module_data_in[7] ,
    \sw_166_module_data_in[6] ,
    \sw_166_module_data_in[5] ,
    \sw_166_module_data_in[4] ,
    \sw_166_module_data_in[3] ,
    \sw_166_module_data_in[2] ,
    \sw_166_module_data_in[1] ,
    \sw_166_module_data_in[0] }),
    .module_data_out({\sw_166_module_data_out[7] ,
    \sw_166_module_data_out[6] ,
    \sw_166_module_data_out[5] ,
    \sw_166_module_data_out[4] ,
    \sw_166_module_data_out[3] ,
    \sw_166_module_data_out[2] ,
    \sw_166_module_data_out[1] ,
    \sw_166_module_data_out[0] }));
 scanchain scanchain_167 (.clk_in(sw_166_clk_out),
    .clk_out(sw_167_clk_out),
    .data_in(sw_166_data_out),
    .data_out(sw_167_data_out),
    .latch_enable_in(sw_166_latch_out),
    .latch_enable_out(sw_167_latch_out),
    .scan_select_in(sw_166_scan_out),
    .scan_select_out(sw_167_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_167_module_data_in[7] ,
    \sw_167_module_data_in[6] ,
    \sw_167_module_data_in[5] ,
    \sw_167_module_data_in[4] ,
    \sw_167_module_data_in[3] ,
    \sw_167_module_data_in[2] ,
    \sw_167_module_data_in[1] ,
    \sw_167_module_data_in[0] }),
    .module_data_out({\sw_167_module_data_out[7] ,
    \sw_167_module_data_out[6] ,
    \sw_167_module_data_out[5] ,
    \sw_167_module_data_out[4] ,
    \sw_167_module_data_out[3] ,
    \sw_167_module_data_out[2] ,
    \sw_167_module_data_out[1] ,
    \sw_167_module_data_out[0] }));
 scanchain scanchain_168 (.clk_in(sw_167_clk_out),
    .clk_out(sw_168_clk_out),
    .data_in(sw_167_data_out),
    .data_out(sw_168_data_out),
    .latch_enable_in(sw_167_latch_out),
    .latch_enable_out(sw_168_latch_out),
    .scan_select_in(sw_167_scan_out),
    .scan_select_out(sw_168_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_168_module_data_in[7] ,
    \sw_168_module_data_in[6] ,
    \sw_168_module_data_in[5] ,
    \sw_168_module_data_in[4] ,
    \sw_168_module_data_in[3] ,
    \sw_168_module_data_in[2] ,
    \sw_168_module_data_in[1] ,
    \sw_168_module_data_in[0] }),
    .module_data_out({\sw_168_module_data_out[7] ,
    \sw_168_module_data_out[6] ,
    \sw_168_module_data_out[5] ,
    \sw_168_module_data_out[4] ,
    \sw_168_module_data_out[3] ,
    \sw_168_module_data_out[2] ,
    \sw_168_module_data_out[1] ,
    \sw_168_module_data_out[0] }));
 scanchain scanchain_169 (.clk_in(sw_168_clk_out),
    .clk_out(sw_169_clk_out),
    .data_in(sw_168_data_out),
    .data_out(sw_169_data_out),
    .latch_enable_in(sw_168_latch_out),
    .latch_enable_out(sw_169_latch_out),
    .scan_select_in(sw_168_scan_out),
    .scan_select_out(sw_169_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_169_module_data_in[7] ,
    \sw_169_module_data_in[6] ,
    \sw_169_module_data_in[5] ,
    \sw_169_module_data_in[4] ,
    \sw_169_module_data_in[3] ,
    \sw_169_module_data_in[2] ,
    \sw_169_module_data_in[1] ,
    \sw_169_module_data_in[0] }),
    .module_data_out({\sw_169_module_data_out[7] ,
    \sw_169_module_data_out[6] ,
    \sw_169_module_data_out[5] ,
    \sw_169_module_data_out[4] ,
    \sw_169_module_data_out[3] ,
    \sw_169_module_data_out[2] ,
    \sw_169_module_data_out[1] ,
    \sw_169_module_data_out[0] }));
 scanchain scanchain_17 (.clk_in(sw_016_clk_out),
    .clk_out(sw_017_clk_out),
    .data_in(sw_016_data_out),
    .data_out(sw_017_data_out),
    .latch_enable_in(sw_016_latch_out),
    .latch_enable_out(sw_017_latch_out),
    .scan_select_in(sw_016_scan_out),
    .scan_select_out(sw_017_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_017_module_data_in[7] ,
    \sw_017_module_data_in[6] ,
    \sw_017_module_data_in[5] ,
    \sw_017_module_data_in[4] ,
    \sw_017_module_data_in[3] ,
    \sw_017_module_data_in[2] ,
    \sw_017_module_data_in[1] ,
    \sw_017_module_data_in[0] }),
    .module_data_out({\sw_017_module_data_out[7] ,
    \sw_017_module_data_out[6] ,
    \sw_017_module_data_out[5] ,
    \sw_017_module_data_out[4] ,
    \sw_017_module_data_out[3] ,
    \sw_017_module_data_out[2] ,
    \sw_017_module_data_out[1] ,
    \sw_017_module_data_out[0] }));
 scanchain scanchain_170 (.clk_in(sw_169_clk_out),
    .clk_out(sw_170_clk_out),
    .data_in(sw_169_data_out),
    .data_out(sw_170_data_out),
    .latch_enable_in(sw_169_latch_out),
    .latch_enable_out(sw_170_latch_out),
    .scan_select_in(sw_169_scan_out),
    .scan_select_out(sw_170_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_170_module_data_in[7] ,
    \sw_170_module_data_in[6] ,
    \sw_170_module_data_in[5] ,
    \sw_170_module_data_in[4] ,
    \sw_170_module_data_in[3] ,
    \sw_170_module_data_in[2] ,
    \sw_170_module_data_in[1] ,
    \sw_170_module_data_in[0] }),
    .module_data_out({\sw_170_module_data_out[7] ,
    \sw_170_module_data_out[6] ,
    \sw_170_module_data_out[5] ,
    \sw_170_module_data_out[4] ,
    \sw_170_module_data_out[3] ,
    \sw_170_module_data_out[2] ,
    \sw_170_module_data_out[1] ,
    \sw_170_module_data_out[0] }));
 scanchain scanchain_171 (.clk_in(sw_170_clk_out),
    .clk_out(sw_171_clk_out),
    .data_in(sw_170_data_out),
    .data_out(sw_171_data_out),
    .latch_enable_in(sw_170_latch_out),
    .latch_enable_out(sw_171_latch_out),
    .scan_select_in(sw_170_scan_out),
    .scan_select_out(sw_171_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_171_module_data_in[7] ,
    \sw_171_module_data_in[6] ,
    \sw_171_module_data_in[5] ,
    \sw_171_module_data_in[4] ,
    \sw_171_module_data_in[3] ,
    \sw_171_module_data_in[2] ,
    \sw_171_module_data_in[1] ,
    \sw_171_module_data_in[0] }),
    .module_data_out({\sw_171_module_data_out[7] ,
    \sw_171_module_data_out[6] ,
    \sw_171_module_data_out[5] ,
    \sw_171_module_data_out[4] ,
    \sw_171_module_data_out[3] ,
    \sw_171_module_data_out[2] ,
    \sw_171_module_data_out[1] ,
    \sw_171_module_data_out[0] }));
 scanchain scanchain_172 (.clk_in(sw_171_clk_out),
    .clk_out(sw_172_clk_out),
    .data_in(sw_171_data_out),
    .data_out(sw_172_data_out),
    .latch_enable_in(sw_171_latch_out),
    .latch_enable_out(sw_172_latch_out),
    .scan_select_in(sw_171_scan_out),
    .scan_select_out(sw_172_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_172_module_data_in[7] ,
    \sw_172_module_data_in[6] ,
    \sw_172_module_data_in[5] ,
    \sw_172_module_data_in[4] ,
    \sw_172_module_data_in[3] ,
    \sw_172_module_data_in[2] ,
    \sw_172_module_data_in[1] ,
    \sw_172_module_data_in[0] }),
    .module_data_out({\sw_172_module_data_out[7] ,
    \sw_172_module_data_out[6] ,
    \sw_172_module_data_out[5] ,
    \sw_172_module_data_out[4] ,
    \sw_172_module_data_out[3] ,
    \sw_172_module_data_out[2] ,
    \sw_172_module_data_out[1] ,
    \sw_172_module_data_out[0] }));
 scanchain scanchain_173 (.clk_in(sw_172_clk_out),
    .clk_out(sw_173_clk_out),
    .data_in(sw_172_data_out),
    .data_out(sw_173_data_out),
    .latch_enable_in(sw_172_latch_out),
    .latch_enable_out(sw_173_latch_out),
    .scan_select_in(sw_172_scan_out),
    .scan_select_out(sw_173_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_173_module_data_in[7] ,
    \sw_173_module_data_in[6] ,
    \sw_173_module_data_in[5] ,
    \sw_173_module_data_in[4] ,
    \sw_173_module_data_in[3] ,
    \sw_173_module_data_in[2] ,
    \sw_173_module_data_in[1] ,
    \sw_173_module_data_in[0] }),
    .module_data_out({\sw_173_module_data_out[7] ,
    \sw_173_module_data_out[6] ,
    \sw_173_module_data_out[5] ,
    \sw_173_module_data_out[4] ,
    \sw_173_module_data_out[3] ,
    \sw_173_module_data_out[2] ,
    \sw_173_module_data_out[1] ,
    \sw_173_module_data_out[0] }));
 scanchain scanchain_174 (.clk_in(sw_173_clk_out),
    .clk_out(sw_174_clk_out),
    .data_in(sw_173_data_out),
    .data_out(sw_174_data_out),
    .latch_enable_in(sw_173_latch_out),
    .latch_enable_out(sw_174_latch_out),
    .scan_select_in(sw_173_scan_out),
    .scan_select_out(sw_174_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_174_module_data_in[7] ,
    \sw_174_module_data_in[6] ,
    \sw_174_module_data_in[5] ,
    \sw_174_module_data_in[4] ,
    \sw_174_module_data_in[3] ,
    \sw_174_module_data_in[2] ,
    \sw_174_module_data_in[1] ,
    \sw_174_module_data_in[0] }),
    .module_data_out({\sw_174_module_data_out[7] ,
    \sw_174_module_data_out[6] ,
    \sw_174_module_data_out[5] ,
    \sw_174_module_data_out[4] ,
    \sw_174_module_data_out[3] ,
    \sw_174_module_data_out[2] ,
    \sw_174_module_data_out[1] ,
    \sw_174_module_data_out[0] }));
 scanchain scanchain_175 (.clk_in(sw_174_clk_out),
    .clk_out(sw_175_clk_out),
    .data_in(sw_174_data_out),
    .data_out(sw_175_data_out),
    .latch_enable_in(sw_174_latch_out),
    .latch_enable_out(sw_175_latch_out),
    .scan_select_in(sw_174_scan_out),
    .scan_select_out(sw_175_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_175_module_data_in[7] ,
    \sw_175_module_data_in[6] ,
    \sw_175_module_data_in[5] ,
    \sw_175_module_data_in[4] ,
    \sw_175_module_data_in[3] ,
    \sw_175_module_data_in[2] ,
    \sw_175_module_data_in[1] ,
    \sw_175_module_data_in[0] }),
    .module_data_out({\sw_175_module_data_out[7] ,
    \sw_175_module_data_out[6] ,
    \sw_175_module_data_out[5] ,
    \sw_175_module_data_out[4] ,
    \sw_175_module_data_out[3] ,
    \sw_175_module_data_out[2] ,
    \sw_175_module_data_out[1] ,
    \sw_175_module_data_out[0] }));
 scanchain scanchain_176 (.clk_in(sw_175_clk_out),
    .clk_out(sw_176_clk_out),
    .data_in(sw_175_data_out),
    .data_out(sw_176_data_out),
    .latch_enable_in(sw_175_latch_out),
    .latch_enable_out(sw_176_latch_out),
    .scan_select_in(sw_175_scan_out),
    .scan_select_out(sw_176_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_176_module_data_in[7] ,
    \sw_176_module_data_in[6] ,
    \sw_176_module_data_in[5] ,
    \sw_176_module_data_in[4] ,
    \sw_176_module_data_in[3] ,
    \sw_176_module_data_in[2] ,
    \sw_176_module_data_in[1] ,
    \sw_176_module_data_in[0] }),
    .module_data_out({\sw_176_module_data_out[7] ,
    \sw_176_module_data_out[6] ,
    \sw_176_module_data_out[5] ,
    \sw_176_module_data_out[4] ,
    \sw_176_module_data_out[3] ,
    \sw_176_module_data_out[2] ,
    \sw_176_module_data_out[1] ,
    \sw_176_module_data_out[0] }));
 scanchain scanchain_177 (.clk_in(sw_176_clk_out),
    .clk_out(sw_177_clk_out),
    .data_in(sw_176_data_out),
    .data_out(sw_177_data_out),
    .latch_enable_in(sw_176_latch_out),
    .latch_enable_out(sw_177_latch_out),
    .scan_select_in(sw_176_scan_out),
    .scan_select_out(sw_177_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_177_module_data_in[7] ,
    \sw_177_module_data_in[6] ,
    \sw_177_module_data_in[5] ,
    \sw_177_module_data_in[4] ,
    \sw_177_module_data_in[3] ,
    \sw_177_module_data_in[2] ,
    \sw_177_module_data_in[1] ,
    \sw_177_module_data_in[0] }),
    .module_data_out({\sw_177_module_data_out[7] ,
    \sw_177_module_data_out[6] ,
    \sw_177_module_data_out[5] ,
    \sw_177_module_data_out[4] ,
    \sw_177_module_data_out[3] ,
    \sw_177_module_data_out[2] ,
    \sw_177_module_data_out[1] ,
    \sw_177_module_data_out[0] }));
 scanchain scanchain_178 (.clk_in(sw_177_clk_out),
    .clk_out(sw_178_clk_out),
    .data_in(sw_177_data_out),
    .data_out(sw_178_data_out),
    .latch_enable_in(sw_177_latch_out),
    .latch_enable_out(sw_178_latch_out),
    .scan_select_in(sw_177_scan_out),
    .scan_select_out(sw_178_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_178_module_data_in[7] ,
    \sw_178_module_data_in[6] ,
    \sw_178_module_data_in[5] ,
    \sw_178_module_data_in[4] ,
    \sw_178_module_data_in[3] ,
    \sw_178_module_data_in[2] ,
    \sw_178_module_data_in[1] ,
    \sw_178_module_data_in[0] }),
    .module_data_out({\sw_178_module_data_out[7] ,
    \sw_178_module_data_out[6] ,
    \sw_178_module_data_out[5] ,
    \sw_178_module_data_out[4] ,
    \sw_178_module_data_out[3] ,
    \sw_178_module_data_out[2] ,
    \sw_178_module_data_out[1] ,
    \sw_178_module_data_out[0] }));
 scanchain scanchain_179 (.clk_in(sw_178_clk_out),
    .clk_out(sw_179_clk_out),
    .data_in(sw_178_data_out),
    .data_out(sw_179_data_out),
    .latch_enable_in(sw_178_latch_out),
    .latch_enable_out(sw_179_latch_out),
    .scan_select_in(sw_178_scan_out),
    .scan_select_out(sw_179_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_179_module_data_in[7] ,
    \sw_179_module_data_in[6] ,
    \sw_179_module_data_in[5] ,
    \sw_179_module_data_in[4] ,
    \sw_179_module_data_in[3] ,
    \sw_179_module_data_in[2] ,
    \sw_179_module_data_in[1] ,
    \sw_179_module_data_in[0] }),
    .module_data_out({\sw_179_module_data_out[7] ,
    \sw_179_module_data_out[6] ,
    \sw_179_module_data_out[5] ,
    \sw_179_module_data_out[4] ,
    \sw_179_module_data_out[3] ,
    \sw_179_module_data_out[2] ,
    \sw_179_module_data_out[1] ,
    \sw_179_module_data_out[0] }));
 scanchain scanchain_18 (.clk_in(sw_017_clk_out),
    .clk_out(sw_018_clk_out),
    .data_in(sw_017_data_out),
    .data_out(sw_018_data_out),
    .latch_enable_in(sw_017_latch_out),
    .latch_enable_out(sw_018_latch_out),
    .scan_select_in(sw_017_scan_out),
    .scan_select_out(sw_018_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_018_module_data_in[7] ,
    \sw_018_module_data_in[6] ,
    \sw_018_module_data_in[5] ,
    \sw_018_module_data_in[4] ,
    \sw_018_module_data_in[3] ,
    \sw_018_module_data_in[2] ,
    \sw_018_module_data_in[1] ,
    \sw_018_module_data_in[0] }),
    .module_data_out({\sw_018_module_data_out[7] ,
    \sw_018_module_data_out[6] ,
    \sw_018_module_data_out[5] ,
    \sw_018_module_data_out[4] ,
    \sw_018_module_data_out[3] ,
    \sw_018_module_data_out[2] ,
    \sw_018_module_data_out[1] ,
    \sw_018_module_data_out[0] }));
 scanchain scanchain_180 (.clk_in(sw_179_clk_out),
    .clk_out(sw_180_clk_out),
    .data_in(sw_179_data_out),
    .data_out(sw_180_data_out),
    .latch_enable_in(sw_179_latch_out),
    .latch_enable_out(sw_180_latch_out),
    .scan_select_in(sw_179_scan_out),
    .scan_select_out(sw_180_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_180_module_data_in[7] ,
    \sw_180_module_data_in[6] ,
    \sw_180_module_data_in[5] ,
    \sw_180_module_data_in[4] ,
    \sw_180_module_data_in[3] ,
    \sw_180_module_data_in[2] ,
    \sw_180_module_data_in[1] ,
    \sw_180_module_data_in[0] }),
    .module_data_out({\sw_180_module_data_out[7] ,
    \sw_180_module_data_out[6] ,
    \sw_180_module_data_out[5] ,
    \sw_180_module_data_out[4] ,
    \sw_180_module_data_out[3] ,
    \sw_180_module_data_out[2] ,
    \sw_180_module_data_out[1] ,
    \sw_180_module_data_out[0] }));
 scanchain scanchain_181 (.clk_in(sw_180_clk_out),
    .clk_out(sw_181_clk_out),
    .data_in(sw_180_data_out),
    .data_out(sw_181_data_out),
    .latch_enable_in(sw_180_latch_out),
    .latch_enable_out(sw_181_latch_out),
    .scan_select_in(sw_180_scan_out),
    .scan_select_out(sw_181_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_181_module_data_in[7] ,
    \sw_181_module_data_in[6] ,
    \sw_181_module_data_in[5] ,
    \sw_181_module_data_in[4] ,
    \sw_181_module_data_in[3] ,
    \sw_181_module_data_in[2] ,
    \sw_181_module_data_in[1] ,
    \sw_181_module_data_in[0] }),
    .module_data_out({\sw_181_module_data_out[7] ,
    \sw_181_module_data_out[6] ,
    \sw_181_module_data_out[5] ,
    \sw_181_module_data_out[4] ,
    \sw_181_module_data_out[3] ,
    \sw_181_module_data_out[2] ,
    \sw_181_module_data_out[1] ,
    \sw_181_module_data_out[0] }));
 scanchain scanchain_182 (.clk_in(sw_181_clk_out),
    .clk_out(sw_182_clk_out),
    .data_in(sw_181_data_out),
    .data_out(sw_182_data_out),
    .latch_enable_in(sw_181_latch_out),
    .latch_enable_out(sw_182_latch_out),
    .scan_select_in(sw_181_scan_out),
    .scan_select_out(sw_182_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_182_module_data_in[7] ,
    \sw_182_module_data_in[6] ,
    \sw_182_module_data_in[5] ,
    \sw_182_module_data_in[4] ,
    \sw_182_module_data_in[3] ,
    \sw_182_module_data_in[2] ,
    \sw_182_module_data_in[1] ,
    \sw_182_module_data_in[0] }),
    .module_data_out({\sw_182_module_data_out[7] ,
    \sw_182_module_data_out[6] ,
    \sw_182_module_data_out[5] ,
    \sw_182_module_data_out[4] ,
    \sw_182_module_data_out[3] ,
    \sw_182_module_data_out[2] ,
    \sw_182_module_data_out[1] ,
    \sw_182_module_data_out[0] }));
 scanchain scanchain_183 (.clk_in(sw_182_clk_out),
    .clk_out(sw_183_clk_out),
    .data_in(sw_182_data_out),
    .data_out(sw_183_data_out),
    .latch_enable_in(sw_182_latch_out),
    .latch_enable_out(sw_183_latch_out),
    .scan_select_in(sw_182_scan_out),
    .scan_select_out(sw_183_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_183_module_data_in[7] ,
    \sw_183_module_data_in[6] ,
    \sw_183_module_data_in[5] ,
    \sw_183_module_data_in[4] ,
    \sw_183_module_data_in[3] ,
    \sw_183_module_data_in[2] ,
    \sw_183_module_data_in[1] ,
    \sw_183_module_data_in[0] }),
    .module_data_out({\sw_183_module_data_out[7] ,
    \sw_183_module_data_out[6] ,
    \sw_183_module_data_out[5] ,
    \sw_183_module_data_out[4] ,
    \sw_183_module_data_out[3] ,
    \sw_183_module_data_out[2] ,
    \sw_183_module_data_out[1] ,
    \sw_183_module_data_out[0] }));
 scanchain scanchain_184 (.clk_in(sw_183_clk_out),
    .clk_out(sw_184_clk_out),
    .data_in(sw_183_data_out),
    .data_out(sw_184_data_out),
    .latch_enable_in(sw_183_latch_out),
    .latch_enable_out(sw_184_latch_out),
    .scan_select_in(sw_183_scan_out),
    .scan_select_out(sw_184_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_184_module_data_in[7] ,
    \sw_184_module_data_in[6] ,
    \sw_184_module_data_in[5] ,
    \sw_184_module_data_in[4] ,
    \sw_184_module_data_in[3] ,
    \sw_184_module_data_in[2] ,
    \sw_184_module_data_in[1] ,
    \sw_184_module_data_in[0] }),
    .module_data_out({\sw_184_module_data_out[7] ,
    \sw_184_module_data_out[6] ,
    \sw_184_module_data_out[5] ,
    \sw_184_module_data_out[4] ,
    \sw_184_module_data_out[3] ,
    \sw_184_module_data_out[2] ,
    \sw_184_module_data_out[1] ,
    \sw_184_module_data_out[0] }));
 scanchain scanchain_185 (.clk_in(sw_184_clk_out),
    .clk_out(sw_185_clk_out),
    .data_in(sw_184_data_out),
    .data_out(sw_185_data_out),
    .latch_enable_in(sw_184_latch_out),
    .latch_enable_out(sw_185_latch_out),
    .scan_select_in(sw_184_scan_out),
    .scan_select_out(sw_185_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_185_module_data_in[7] ,
    \sw_185_module_data_in[6] ,
    \sw_185_module_data_in[5] ,
    \sw_185_module_data_in[4] ,
    \sw_185_module_data_in[3] ,
    \sw_185_module_data_in[2] ,
    \sw_185_module_data_in[1] ,
    \sw_185_module_data_in[0] }),
    .module_data_out({\sw_185_module_data_out[7] ,
    \sw_185_module_data_out[6] ,
    \sw_185_module_data_out[5] ,
    \sw_185_module_data_out[4] ,
    \sw_185_module_data_out[3] ,
    \sw_185_module_data_out[2] ,
    \sw_185_module_data_out[1] ,
    \sw_185_module_data_out[0] }));
 scanchain scanchain_186 (.clk_in(sw_185_clk_out),
    .clk_out(sw_186_clk_out),
    .data_in(sw_185_data_out),
    .data_out(sw_186_data_out),
    .latch_enable_in(sw_185_latch_out),
    .latch_enable_out(sw_186_latch_out),
    .scan_select_in(sw_185_scan_out),
    .scan_select_out(sw_186_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_186_module_data_in[7] ,
    \sw_186_module_data_in[6] ,
    \sw_186_module_data_in[5] ,
    \sw_186_module_data_in[4] ,
    \sw_186_module_data_in[3] ,
    \sw_186_module_data_in[2] ,
    \sw_186_module_data_in[1] ,
    \sw_186_module_data_in[0] }),
    .module_data_out({\sw_186_module_data_out[7] ,
    \sw_186_module_data_out[6] ,
    \sw_186_module_data_out[5] ,
    \sw_186_module_data_out[4] ,
    \sw_186_module_data_out[3] ,
    \sw_186_module_data_out[2] ,
    \sw_186_module_data_out[1] ,
    \sw_186_module_data_out[0] }));
 scanchain scanchain_187 (.clk_in(sw_186_clk_out),
    .clk_out(sw_187_clk_out),
    .data_in(sw_186_data_out),
    .data_out(sw_187_data_out),
    .latch_enable_in(sw_186_latch_out),
    .latch_enable_out(sw_187_latch_out),
    .scan_select_in(sw_186_scan_out),
    .scan_select_out(sw_187_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_187_module_data_in[7] ,
    \sw_187_module_data_in[6] ,
    \sw_187_module_data_in[5] ,
    \sw_187_module_data_in[4] ,
    \sw_187_module_data_in[3] ,
    \sw_187_module_data_in[2] ,
    \sw_187_module_data_in[1] ,
    \sw_187_module_data_in[0] }),
    .module_data_out({\sw_187_module_data_out[7] ,
    \sw_187_module_data_out[6] ,
    \sw_187_module_data_out[5] ,
    \sw_187_module_data_out[4] ,
    \sw_187_module_data_out[3] ,
    \sw_187_module_data_out[2] ,
    \sw_187_module_data_out[1] ,
    \sw_187_module_data_out[0] }));
 scanchain scanchain_188 (.clk_in(sw_187_clk_out),
    .clk_out(sw_188_clk_out),
    .data_in(sw_187_data_out),
    .data_out(sw_188_data_out),
    .latch_enable_in(sw_187_latch_out),
    .latch_enable_out(sw_188_latch_out),
    .scan_select_in(sw_187_scan_out),
    .scan_select_out(sw_188_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_188_module_data_in[7] ,
    \sw_188_module_data_in[6] ,
    \sw_188_module_data_in[5] ,
    \sw_188_module_data_in[4] ,
    \sw_188_module_data_in[3] ,
    \sw_188_module_data_in[2] ,
    \sw_188_module_data_in[1] ,
    \sw_188_module_data_in[0] }),
    .module_data_out({\sw_188_module_data_out[7] ,
    \sw_188_module_data_out[6] ,
    \sw_188_module_data_out[5] ,
    \sw_188_module_data_out[4] ,
    \sw_188_module_data_out[3] ,
    \sw_188_module_data_out[2] ,
    \sw_188_module_data_out[1] ,
    \sw_188_module_data_out[0] }));
 scanchain scanchain_189 (.clk_in(sw_188_clk_out),
    .clk_out(sw_189_clk_out),
    .data_in(sw_188_data_out),
    .data_out(sw_189_data_out),
    .latch_enable_in(sw_188_latch_out),
    .latch_enable_out(sw_189_latch_out),
    .scan_select_in(sw_188_scan_out),
    .scan_select_out(sw_189_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_189_module_data_in[7] ,
    \sw_189_module_data_in[6] ,
    \sw_189_module_data_in[5] ,
    \sw_189_module_data_in[4] ,
    \sw_189_module_data_in[3] ,
    \sw_189_module_data_in[2] ,
    \sw_189_module_data_in[1] ,
    \sw_189_module_data_in[0] }),
    .module_data_out({\sw_189_module_data_out[7] ,
    \sw_189_module_data_out[6] ,
    \sw_189_module_data_out[5] ,
    \sw_189_module_data_out[4] ,
    \sw_189_module_data_out[3] ,
    \sw_189_module_data_out[2] ,
    \sw_189_module_data_out[1] ,
    \sw_189_module_data_out[0] }));
 scanchain scanchain_19 (.clk_in(sw_018_clk_out),
    .clk_out(sw_019_clk_out),
    .data_in(sw_018_data_out),
    .data_out(sw_019_data_out),
    .latch_enable_in(sw_018_latch_out),
    .latch_enable_out(sw_019_latch_out),
    .scan_select_in(sw_018_scan_out),
    .scan_select_out(sw_019_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_019_module_data_in[7] ,
    \sw_019_module_data_in[6] ,
    \sw_019_module_data_in[5] ,
    \sw_019_module_data_in[4] ,
    \sw_019_module_data_in[3] ,
    \sw_019_module_data_in[2] ,
    \sw_019_module_data_in[1] ,
    \sw_019_module_data_in[0] }),
    .module_data_out({\sw_019_module_data_out[7] ,
    \sw_019_module_data_out[6] ,
    \sw_019_module_data_out[5] ,
    \sw_019_module_data_out[4] ,
    \sw_019_module_data_out[3] ,
    \sw_019_module_data_out[2] ,
    \sw_019_module_data_out[1] ,
    \sw_019_module_data_out[0] }));
 scanchain scanchain_190 (.clk_in(sw_189_clk_out),
    .clk_out(sw_190_clk_out),
    .data_in(sw_189_data_out),
    .data_out(sw_190_data_out),
    .latch_enable_in(sw_189_latch_out),
    .latch_enable_out(sw_190_latch_out),
    .scan_select_in(sw_189_scan_out),
    .scan_select_out(sw_190_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_190_module_data_in[7] ,
    \sw_190_module_data_in[6] ,
    \sw_190_module_data_in[5] ,
    \sw_190_module_data_in[4] ,
    \sw_190_module_data_in[3] ,
    \sw_190_module_data_in[2] ,
    \sw_190_module_data_in[1] ,
    \sw_190_module_data_in[0] }),
    .module_data_out({\sw_190_module_data_out[7] ,
    \sw_190_module_data_out[6] ,
    \sw_190_module_data_out[5] ,
    \sw_190_module_data_out[4] ,
    \sw_190_module_data_out[3] ,
    \sw_190_module_data_out[2] ,
    \sw_190_module_data_out[1] ,
    \sw_190_module_data_out[0] }));
 scanchain scanchain_191 (.clk_in(sw_190_clk_out),
    .clk_out(sw_191_clk_out),
    .data_in(sw_190_data_out),
    .data_out(sw_191_data_out),
    .latch_enable_in(sw_190_latch_out),
    .latch_enable_out(sw_191_latch_out),
    .scan_select_in(sw_190_scan_out),
    .scan_select_out(sw_191_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_191_module_data_in[7] ,
    \sw_191_module_data_in[6] ,
    \sw_191_module_data_in[5] ,
    \sw_191_module_data_in[4] ,
    \sw_191_module_data_in[3] ,
    \sw_191_module_data_in[2] ,
    \sw_191_module_data_in[1] ,
    \sw_191_module_data_in[0] }),
    .module_data_out({\sw_191_module_data_out[7] ,
    \sw_191_module_data_out[6] ,
    \sw_191_module_data_out[5] ,
    \sw_191_module_data_out[4] ,
    \sw_191_module_data_out[3] ,
    \sw_191_module_data_out[2] ,
    \sw_191_module_data_out[1] ,
    \sw_191_module_data_out[0] }));
 scanchain scanchain_192 (.clk_in(sw_191_clk_out),
    .clk_out(sw_192_clk_out),
    .data_in(sw_191_data_out),
    .data_out(sw_192_data_out),
    .latch_enable_in(sw_191_latch_out),
    .latch_enable_out(sw_192_latch_out),
    .scan_select_in(sw_191_scan_out),
    .scan_select_out(sw_192_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_192_module_data_in[7] ,
    \sw_192_module_data_in[6] ,
    \sw_192_module_data_in[5] ,
    \sw_192_module_data_in[4] ,
    \sw_192_module_data_in[3] ,
    \sw_192_module_data_in[2] ,
    \sw_192_module_data_in[1] ,
    \sw_192_module_data_in[0] }),
    .module_data_out({\sw_192_module_data_out[7] ,
    \sw_192_module_data_out[6] ,
    \sw_192_module_data_out[5] ,
    \sw_192_module_data_out[4] ,
    \sw_192_module_data_out[3] ,
    \sw_192_module_data_out[2] ,
    \sw_192_module_data_out[1] ,
    \sw_192_module_data_out[0] }));
 scanchain scanchain_193 (.clk_in(sw_192_clk_out),
    .clk_out(sw_193_clk_out),
    .data_in(sw_192_data_out),
    .data_out(sw_193_data_out),
    .latch_enable_in(sw_192_latch_out),
    .latch_enable_out(sw_193_latch_out),
    .scan_select_in(sw_192_scan_out),
    .scan_select_out(sw_193_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_193_module_data_in[7] ,
    \sw_193_module_data_in[6] ,
    \sw_193_module_data_in[5] ,
    \sw_193_module_data_in[4] ,
    \sw_193_module_data_in[3] ,
    \sw_193_module_data_in[2] ,
    \sw_193_module_data_in[1] ,
    \sw_193_module_data_in[0] }),
    .module_data_out({\sw_193_module_data_out[7] ,
    \sw_193_module_data_out[6] ,
    \sw_193_module_data_out[5] ,
    \sw_193_module_data_out[4] ,
    \sw_193_module_data_out[3] ,
    \sw_193_module_data_out[2] ,
    \sw_193_module_data_out[1] ,
    \sw_193_module_data_out[0] }));
 scanchain scanchain_194 (.clk_in(sw_193_clk_out),
    .clk_out(sw_194_clk_out),
    .data_in(sw_193_data_out),
    .data_out(sw_194_data_out),
    .latch_enable_in(sw_193_latch_out),
    .latch_enable_out(sw_194_latch_out),
    .scan_select_in(sw_193_scan_out),
    .scan_select_out(sw_194_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_194_module_data_in[7] ,
    \sw_194_module_data_in[6] ,
    \sw_194_module_data_in[5] ,
    \sw_194_module_data_in[4] ,
    \sw_194_module_data_in[3] ,
    \sw_194_module_data_in[2] ,
    \sw_194_module_data_in[1] ,
    \sw_194_module_data_in[0] }),
    .module_data_out({\sw_194_module_data_out[7] ,
    \sw_194_module_data_out[6] ,
    \sw_194_module_data_out[5] ,
    \sw_194_module_data_out[4] ,
    \sw_194_module_data_out[3] ,
    \sw_194_module_data_out[2] ,
    \sw_194_module_data_out[1] ,
    \sw_194_module_data_out[0] }));
 scanchain scanchain_195 (.clk_in(sw_194_clk_out),
    .clk_out(sw_195_clk_out),
    .data_in(sw_194_data_out),
    .data_out(sw_195_data_out),
    .latch_enable_in(sw_194_latch_out),
    .latch_enable_out(sw_195_latch_out),
    .scan_select_in(sw_194_scan_out),
    .scan_select_out(sw_195_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_195_module_data_in[7] ,
    \sw_195_module_data_in[6] ,
    \sw_195_module_data_in[5] ,
    \sw_195_module_data_in[4] ,
    \sw_195_module_data_in[3] ,
    \sw_195_module_data_in[2] ,
    \sw_195_module_data_in[1] ,
    \sw_195_module_data_in[0] }),
    .module_data_out({\sw_195_module_data_out[7] ,
    \sw_195_module_data_out[6] ,
    \sw_195_module_data_out[5] ,
    \sw_195_module_data_out[4] ,
    \sw_195_module_data_out[3] ,
    \sw_195_module_data_out[2] ,
    \sw_195_module_data_out[1] ,
    \sw_195_module_data_out[0] }));
 scanchain scanchain_196 (.clk_in(sw_195_clk_out),
    .clk_out(sw_196_clk_out),
    .data_in(sw_195_data_out),
    .data_out(sw_196_data_out),
    .latch_enable_in(sw_195_latch_out),
    .latch_enable_out(sw_196_latch_out),
    .scan_select_in(sw_195_scan_out),
    .scan_select_out(sw_196_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_196_module_data_in[7] ,
    \sw_196_module_data_in[6] ,
    \sw_196_module_data_in[5] ,
    \sw_196_module_data_in[4] ,
    \sw_196_module_data_in[3] ,
    \sw_196_module_data_in[2] ,
    \sw_196_module_data_in[1] ,
    \sw_196_module_data_in[0] }),
    .module_data_out({\sw_196_module_data_out[7] ,
    \sw_196_module_data_out[6] ,
    \sw_196_module_data_out[5] ,
    \sw_196_module_data_out[4] ,
    \sw_196_module_data_out[3] ,
    \sw_196_module_data_out[2] ,
    \sw_196_module_data_out[1] ,
    \sw_196_module_data_out[0] }));
 scanchain scanchain_197 (.clk_in(sw_196_clk_out),
    .clk_out(sw_197_clk_out),
    .data_in(sw_196_data_out),
    .data_out(sw_197_data_out),
    .latch_enable_in(sw_196_latch_out),
    .latch_enable_out(sw_197_latch_out),
    .scan_select_in(sw_196_scan_out),
    .scan_select_out(sw_197_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_197_module_data_in[7] ,
    \sw_197_module_data_in[6] ,
    \sw_197_module_data_in[5] ,
    \sw_197_module_data_in[4] ,
    \sw_197_module_data_in[3] ,
    \sw_197_module_data_in[2] ,
    \sw_197_module_data_in[1] ,
    \sw_197_module_data_in[0] }),
    .module_data_out({\sw_197_module_data_out[7] ,
    \sw_197_module_data_out[6] ,
    \sw_197_module_data_out[5] ,
    \sw_197_module_data_out[4] ,
    \sw_197_module_data_out[3] ,
    \sw_197_module_data_out[2] ,
    \sw_197_module_data_out[1] ,
    \sw_197_module_data_out[0] }));
 scanchain scanchain_198 (.clk_in(sw_197_clk_out),
    .clk_out(sw_198_clk_out),
    .data_in(sw_197_data_out),
    .data_out(sw_198_data_out),
    .latch_enable_in(sw_197_latch_out),
    .latch_enable_out(sw_198_latch_out),
    .scan_select_in(sw_197_scan_out),
    .scan_select_out(sw_198_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_198_module_data_in[7] ,
    \sw_198_module_data_in[6] ,
    \sw_198_module_data_in[5] ,
    \sw_198_module_data_in[4] ,
    \sw_198_module_data_in[3] ,
    \sw_198_module_data_in[2] ,
    \sw_198_module_data_in[1] ,
    \sw_198_module_data_in[0] }),
    .module_data_out({\sw_198_module_data_out[7] ,
    \sw_198_module_data_out[6] ,
    \sw_198_module_data_out[5] ,
    \sw_198_module_data_out[4] ,
    \sw_198_module_data_out[3] ,
    \sw_198_module_data_out[2] ,
    \sw_198_module_data_out[1] ,
    \sw_198_module_data_out[0] }));
 scanchain scanchain_199 (.clk_in(sw_198_clk_out),
    .clk_out(sw_199_clk_out),
    .data_in(sw_198_data_out),
    .data_out(sw_199_data_out),
    .latch_enable_in(sw_198_latch_out),
    .latch_enable_out(sw_199_latch_out),
    .scan_select_in(sw_198_scan_out),
    .scan_select_out(sw_199_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_199_module_data_in[7] ,
    \sw_199_module_data_in[6] ,
    \sw_199_module_data_in[5] ,
    \sw_199_module_data_in[4] ,
    \sw_199_module_data_in[3] ,
    \sw_199_module_data_in[2] ,
    \sw_199_module_data_in[1] ,
    \sw_199_module_data_in[0] }),
    .module_data_out({\sw_199_module_data_out[7] ,
    \sw_199_module_data_out[6] ,
    \sw_199_module_data_out[5] ,
    \sw_199_module_data_out[4] ,
    \sw_199_module_data_out[3] ,
    \sw_199_module_data_out[2] ,
    \sw_199_module_data_out[1] ,
    \sw_199_module_data_out[0] }));
 scanchain scanchain_2 (.clk_in(sw_001_clk_out),
    .clk_out(sw_002_clk_out),
    .data_in(sw_001_data_out),
    .data_out(sw_002_data_out),
    .latch_enable_in(sw_001_latch_out),
    .latch_enable_out(sw_002_latch_out),
    .scan_select_in(sw_001_scan_out),
    .scan_select_out(sw_002_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_002_module_data_in[7] ,
    \sw_002_module_data_in[6] ,
    \sw_002_module_data_in[5] ,
    \sw_002_module_data_in[4] ,
    \sw_002_module_data_in[3] ,
    \sw_002_module_data_in[2] ,
    \sw_002_module_data_in[1] ,
    \sw_002_module_data_in[0] }),
    .module_data_out({\sw_002_module_data_out[7] ,
    \sw_002_module_data_out[6] ,
    \sw_002_module_data_out[5] ,
    \sw_002_module_data_out[4] ,
    \sw_002_module_data_out[3] ,
    \sw_002_module_data_out[2] ,
    \sw_002_module_data_out[1] ,
    \sw_002_module_data_out[0] }));
 scanchain scanchain_20 (.clk_in(sw_019_clk_out),
    .clk_out(sw_020_clk_out),
    .data_in(sw_019_data_out),
    .data_out(sw_020_data_out),
    .latch_enable_in(sw_019_latch_out),
    .latch_enable_out(sw_020_latch_out),
    .scan_select_in(sw_019_scan_out),
    .scan_select_out(sw_020_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_020_module_data_in[7] ,
    \sw_020_module_data_in[6] ,
    \sw_020_module_data_in[5] ,
    \sw_020_module_data_in[4] ,
    \sw_020_module_data_in[3] ,
    \sw_020_module_data_in[2] ,
    \sw_020_module_data_in[1] ,
    \sw_020_module_data_in[0] }),
    .module_data_out({\sw_020_module_data_out[7] ,
    \sw_020_module_data_out[6] ,
    \sw_020_module_data_out[5] ,
    \sw_020_module_data_out[4] ,
    \sw_020_module_data_out[3] ,
    \sw_020_module_data_out[2] ,
    \sw_020_module_data_out[1] ,
    \sw_020_module_data_out[0] }));
 scanchain scanchain_200 (.clk_in(sw_199_clk_out),
    .clk_out(sw_200_clk_out),
    .data_in(sw_199_data_out),
    .data_out(sw_200_data_out),
    .latch_enable_in(sw_199_latch_out),
    .latch_enable_out(sw_200_latch_out),
    .scan_select_in(sw_199_scan_out),
    .scan_select_out(sw_200_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_200_module_data_in[7] ,
    \sw_200_module_data_in[6] ,
    \sw_200_module_data_in[5] ,
    \sw_200_module_data_in[4] ,
    \sw_200_module_data_in[3] ,
    \sw_200_module_data_in[2] ,
    \sw_200_module_data_in[1] ,
    \sw_200_module_data_in[0] }),
    .module_data_out({\sw_200_module_data_out[7] ,
    \sw_200_module_data_out[6] ,
    \sw_200_module_data_out[5] ,
    \sw_200_module_data_out[4] ,
    \sw_200_module_data_out[3] ,
    \sw_200_module_data_out[2] ,
    \sw_200_module_data_out[1] ,
    \sw_200_module_data_out[0] }));
 scanchain scanchain_201 (.clk_in(sw_200_clk_out),
    .clk_out(sw_201_clk_out),
    .data_in(sw_200_data_out),
    .data_out(sw_201_data_out),
    .latch_enable_in(sw_200_latch_out),
    .latch_enable_out(sw_201_latch_out),
    .scan_select_in(sw_200_scan_out),
    .scan_select_out(sw_201_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_201_module_data_in[7] ,
    \sw_201_module_data_in[6] ,
    \sw_201_module_data_in[5] ,
    \sw_201_module_data_in[4] ,
    \sw_201_module_data_in[3] ,
    \sw_201_module_data_in[2] ,
    \sw_201_module_data_in[1] ,
    \sw_201_module_data_in[0] }),
    .module_data_out({\sw_201_module_data_out[7] ,
    \sw_201_module_data_out[6] ,
    \sw_201_module_data_out[5] ,
    \sw_201_module_data_out[4] ,
    \sw_201_module_data_out[3] ,
    \sw_201_module_data_out[2] ,
    \sw_201_module_data_out[1] ,
    \sw_201_module_data_out[0] }));
 scanchain scanchain_202 (.clk_in(sw_201_clk_out),
    .clk_out(sw_202_clk_out),
    .data_in(sw_201_data_out),
    .data_out(sw_202_data_out),
    .latch_enable_in(sw_201_latch_out),
    .latch_enable_out(sw_202_latch_out),
    .scan_select_in(sw_201_scan_out),
    .scan_select_out(sw_202_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_202_module_data_in[7] ,
    \sw_202_module_data_in[6] ,
    \sw_202_module_data_in[5] ,
    \sw_202_module_data_in[4] ,
    \sw_202_module_data_in[3] ,
    \sw_202_module_data_in[2] ,
    \sw_202_module_data_in[1] ,
    \sw_202_module_data_in[0] }),
    .module_data_out({\sw_202_module_data_out[7] ,
    \sw_202_module_data_out[6] ,
    \sw_202_module_data_out[5] ,
    \sw_202_module_data_out[4] ,
    \sw_202_module_data_out[3] ,
    \sw_202_module_data_out[2] ,
    \sw_202_module_data_out[1] ,
    \sw_202_module_data_out[0] }));
 scanchain scanchain_203 (.clk_in(sw_202_clk_out),
    .clk_out(sw_203_clk_out),
    .data_in(sw_202_data_out),
    .data_out(sw_203_data_out),
    .latch_enable_in(sw_202_latch_out),
    .latch_enable_out(sw_203_latch_out),
    .scan_select_in(sw_202_scan_out),
    .scan_select_out(sw_203_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_203_module_data_in[7] ,
    \sw_203_module_data_in[6] ,
    \sw_203_module_data_in[5] ,
    \sw_203_module_data_in[4] ,
    \sw_203_module_data_in[3] ,
    \sw_203_module_data_in[2] ,
    \sw_203_module_data_in[1] ,
    \sw_203_module_data_in[0] }),
    .module_data_out({\sw_203_module_data_out[7] ,
    \sw_203_module_data_out[6] ,
    \sw_203_module_data_out[5] ,
    \sw_203_module_data_out[4] ,
    \sw_203_module_data_out[3] ,
    \sw_203_module_data_out[2] ,
    \sw_203_module_data_out[1] ,
    \sw_203_module_data_out[0] }));
 scanchain scanchain_204 (.clk_in(sw_203_clk_out),
    .clk_out(sw_204_clk_out),
    .data_in(sw_203_data_out),
    .data_out(sw_204_data_out),
    .latch_enable_in(sw_203_latch_out),
    .latch_enable_out(sw_204_latch_out),
    .scan_select_in(sw_203_scan_out),
    .scan_select_out(sw_204_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_204_module_data_in[7] ,
    \sw_204_module_data_in[6] ,
    \sw_204_module_data_in[5] ,
    \sw_204_module_data_in[4] ,
    \sw_204_module_data_in[3] ,
    \sw_204_module_data_in[2] ,
    \sw_204_module_data_in[1] ,
    \sw_204_module_data_in[0] }),
    .module_data_out({\sw_204_module_data_out[7] ,
    \sw_204_module_data_out[6] ,
    \sw_204_module_data_out[5] ,
    \sw_204_module_data_out[4] ,
    \sw_204_module_data_out[3] ,
    \sw_204_module_data_out[2] ,
    \sw_204_module_data_out[1] ,
    \sw_204_module_data_out[0] }));
 scanchain scanchain_205 (.clk_in(sw_204_clk_out),
    .clk_out(sw_205_clk_out),
    .data_in(sw_204_data_out),
    .data_out(sw_205_data_out),
    .latch_enable_in(sw_204_latch_out),
    .latch_enable_out(sw_205_latch_out),
    .scan_select_in(sw_204_scan_out),
    .scan_select_out(sw_205_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_205_module_data_in[7] ,
    \sw_205_module_data_in[6] ,
    \sw_205_module_data_in[5] ,
    \sw_205_module_data_in[4] ,
    \sw_205_module_data_in[3] ,
    \sw_205_module_data_in[2] ,
    \sw_205_module_data_in[1] ,
    \sw_205_module_data_in[0] }),
    .module_data_out({\sw_205_module_data_out[7] ,
    \sw_205_module_data_out[6] ,
    \sw_205_module_data_out[5] ,
    \sw_205_module_data_out[4] ,
    \sw_205_module_data_out[3] ,
    \sw_205_module_data_out[2] ,
    \sw_205_module_data_out[1] ,
    \sw_205_module_data_out[0] }));
 scanchain scanchain_206 (.clk_in(sw_205_clk_out),
    .clk_out(sw_206_clk_out),
    .data_in(sw_205_data_out),
    .data_out(sw_206_data_out),
    .latch_enable_in(sw_205_latch_out),
    .latch_enable_out(sw_206_latch_out),
    .scan_select_in(sw_205_scan_out),
    .scan_select_out(sw_206_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_206_module_data_in[7] ,
    \sw_206_module_data_in[6] ,
    \sw_206_module_data_in[5] ,
    \sw_206_module_data_in[4] ,
    \sw_206_module_data_in[3] ,
    \sw_206_module_data_in[2] ,
    \sw_206_module_data_in[1] ,
    \sw_206_module_data_in[0] }),
    .module_data_out({\sw_206_module_data_out[7] ,
    \sw_206_module_data_out[6] ,
    \sw_206_module_data_out[5] ,
    \sw_206_module_data_out[4] ,
    \sw_206_module_data_out[3] ,
    \sw_206_module_data_out[2] ,
    \sw_206_module_data_out[1] ,
    \sw_206_module_data_out[0] }));
 scanchain scanchain_207 (.clk_in(sw_206_clk_out),
    .clk_out(sw_207_clk_out),
    .data_in(sw_206_data_out),
    .data_out(sw_207_data_out),
    .latch_enable_in(sw_206_latch_out),
    .latch_enable_out(sw_207_latch_out),
    .scan_select_in(sw_206_scan_out),
    .scan_select_out(sw_207_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_207_module_data_in[7] ,
    \sw_207_module_data_in[6] ,
    \sw_207_module_data_in[5] ,
    \sw_207_module_data_in[4] ,
    \sw_207_module_data_in[3] ,
    \sw_207_module_data_in[2] ,
    \sw_207_module_data_in[1] ,
    \sw_207_module_data_in[0] }),
    .module_data_out({\sw_207_module_data_out[7] ,
    \sw_207_module_data_out[6] ,
    \sw_207_module_data_out[5] ,
    \sw_207_module_data_out[4] ,
    \sw_207_module_data_out[3] ,
    \sw_207_module_data_out[2] ,
    \sw_207_module_data_out[1] ,
    \sw_207_module_data_out[0] }));
 scanchain scanchain_208 (.clk_in(sw_207_clk_out),
    .clk_out(sw_208_clk_out),
    .data_in(sw_207_data_out),
    .data_out(sw_208_data_out),
    .latch_enable_in(sw_207_latch_out),
    .latch_enable_out(sw_208_latch_out),
    .scan_select_in(sw_207_scan_out),
    .scan_select_out(sw_208_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_208_module_data_in[7] ,
    \sw_208_module_data_in[6] ,
    \sw_208_module_data_in[5] ,
    \sw_208_module_data_in[4] ,
    \sw_208_module_data_in[3] ,
    \sw_208_module_data_in[2] ,
    \sw_208_module_data_in[1] ,
    \sw_208_module_data_in[0] }),
    .module_data_out({\sw_208_module_data_out[7] ,
    \sw_208_module_data_out[6] ,
    \sw_208_module_data_out[5] ,
    \sw_208_module_data_out[4] ,
    \sw_208_module_data_out[3] ,
    \sw_208_module_data_out[2] ,
    \sw_208_module_data_out[1] ,
    \sw_208_module_data_out[0] }));
 scanchain scanchain_209 (.clk_in(sw_208_clk_out),
    .clk_out(sw_209_clk_out),
    .data_in(sw_208_data_out),
    .data_out(sw_209_data_out),
    .latch_enable_in(sw_208_latch_out),
    .latch_enable_out(sw_209_latch_out),
    .scan_select_in(sw_208_scan_out),
    .scan_select_out(sw_209_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_209_module_data_in[7] ,
    \sw_209_module_data_in[6] ,
    \sw_209_module_data_in[5] ,
    \sw_209_module_data_in[4] ,
    \sw_209_module_data_in[3] ,
    \sw_209_module_data_in[2] ,
    \sw_209_module_data_in[1] ,
    \sw_209_module_data_in[0] }),
    .module_data_out({\sw_209_module_data_out[7] ,
    \sw_209_module_data_out[6] ,
    \sw_209_module_data_out[5] ,
    \sw_209_module_data_out[4] ,
    \sw_209_module_data_out[3] ,
    \sw_209_module_data_out[2] ,
    \sw_209_module_data_out[1] ,
    \sw_209_module_data_out[0] }));
 scanchain scanchain_21 (.clk_in(sw_020_clk_out),
    .clk_out(sw_021_clk_out),
    .data_in(sw_020_data_out),
    .data_out(sw_021_data_out),
    .latch_enable_in(sw_020_latch_out),
    .latch_enable_out(sw_021_latch_out),
    .scan_select_in(sw_020_scan_out),
    .scan_select_out(sw_021_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_021_module_data_in[7] ,
    \sw_021_module_data_in[6] ,
    \sw_021_module_data_in[5] ,
    \sw_021_module_data_in[4] ,
    \sw_021_module_data_in[3] ,
    \sw_021_module_data_in[2] ,
    \sw_021_module_data_in[1] ,
    \sw_021_module_data_in[0] }),
    .module_data_out({\sw_021_module_data_out[7] ,
    \sw_021_module_data_out[6] ,
    \sw_021_module_data_out[5] ,
    \sw_021_module_data_out[4] ,
    \sw_021_module_data_out[3] ,
    \sw_021_module_data_out[2] ,
    \sw_021_module_data_out[1] ,
    \sw_021_module_data_out[0] }));
 scanchain scanchain_210 (.clk_in(sw_209_clk_out),
    .clk_out(sw_210_clk_out),
    .data_in(sw_209_data_out),
    .data_out(sw_210_data_out),
    .latch_enable_in(sw_209_latch_out),
    .latch_enable_out(sw_210_latch_out),
    .scan_select_in(sw_209_scan_out),
    .scan_select_out(sw_210_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_210_module_data_in[7] ,
    \sw_210_module_data_in[6] ,
    \sw_210_module_data_in[5] ,
    \sw_210_module_data_in[4] ,
    \sw_210_module_data_in[3] ,
    \sw_210_module_data_in[2] ,
    \sw_210_module_data_in[1] ,
    \sw_210_module_data_in[0] }),
    .module_data_out({\sw_210_module_data_out[7] ,
    \sw_210_module_data_out[6] ,
    \sw_210_module_data_out[5] ,
    \sw_210_module_data_out[4] ,
    \sw_210_module_data_out[3] ,
    \sw_210_module_data_out[2] ,
    \sw_210_module_data_out[1] ,
    \sw_210_module_data_out[0] }));
 scanchain scanchain_211 (.clk_in(sw_210_clk_out),
    .clk_out(sw_211_clk_out),
    .data_in(sw_210_data_out),
    .data_out(sw_211_data_out),
    .latch_enable_in(sw_210_latch_out),
    .latch_enable_out(sw_211_latch_out),
    .scan_select_in(sw_210_scan_out),
    .scan_select_out(sw_211_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_211_module_data_in[7] ,
    \sw_211_module_data_in[6] ,
    \sw_211_module_data_in[5] ,
    \sw_211_module_data_in[4] ,
    \sw_211_module_data_in[3] ,
    \sw_211_module_data_in[2] ,
    \sw_211_module_data_in[1] ,
    \sw_211_module_data_in[0] }),
    .module_data_out({\sw_211_module_data_out[7] ,
    \sw_211_module_data_out[6] ,
    \sw_211_module_data_out[5] ,
    \sw_211_module_data_out[4] ,
    \sw_211_module_data_out[3] ,
    \sw_211_module_data_out[2] ,
    \sw_211_module_data_out[1] ,
    \sw_211_module_data_out[0] }));
 scanchain scanchain_212 (.clk_in(sw_211_clk_out),
    .clk_out(sw_212_clk_out),
    .data_in(sw_211_data_out),
    .data_out(sw_212_data_out),
    .latch_enable_in(sw_211_latch_out),
    .latch_enable_out(sw_212_latch_out),
    .scan_select_in(sw_211_scan_out),
    .scan_select_out(sw_212_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_212_module_data_in[7] ,
    \sw_212_module_data_in[6] ,
    \sw_212_module_data_in[5] ,
    \sw_212_module_data_in[4] ,
    \sw_212_module_data_in[3] ,
    \sw_212_module_data_in[2] ,
    \sw_212_module_data_in[1] ,
    \sw_212_module_data_in[0] }),
    .module_data_out({\sw_212_module_data_out[7] ,
    \sw_212_module_data_out[6] ,
    \sw_212_module_data_out[5] ,
    \sw_212_module_data_out[4] ,
    \sw_212_module_data_out[3] ,
    \sw_212_module_data_out[2] ,
    \sw_212_module_data_out[1] ,
    \sw_212_module_data_out[0] }));
 scanchain scanchain_213 (.clk_in(sw_212_clk_out),
    .clk_out(sw_213_clk_out),
    .data_in(sw_212_data_out),
    .data_out(sw_213_data_out),
    .latch_enable_in(sw_212_latch_out),
    .latch_enable_out(sw_213_latch_out),
    .scan_select_in(sw_212_scan_out),
    .scan_select_out(sw_213_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_213_module_data_in[7] ,
    \sw_213_module_data_in[6] ,
    \sw_213_module_data_in[5] ,
    \sw_213_module_data_in[4] ,
    \sw_213_module_data_in[3] ,
    \sw_213_module_data_in[2] ,
    \sw_213_module_data_in[1] ,
    \sw_213_module_data_in[0] }),
    .module_data_out({\sw_213_module_data_out[7] ,
    \sw_213_module_data_out[6] ,
    \sw_213_module_data_out[5] ,
    \sw_213_module_data_out[4] ,
    \sw_213_module_data_out[3] ,
    \sw_213_module_data_out[2] ,
    \sw_213_module_data_out[1] ,
    \sw_213_module_data_out[0] }));
 scanchain scanchain_214 (.clk_in(sw_213_clk_out),
    .clk_out(sw_214_clk_out),
    .data_in(sw_213_data_out),
    .data_out(sw_214_data_out),
    .latch_enable_in(sw_213_latch_out),
    .latch_enable_out(sw_214_latch_out),
    .scan_select_in(sw_213_scan_out),
    .scan_select_out(sw_214_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_214_module_data_in[7] ,
    \sw_214_module_data_in[6] ,
    \sw_214_module_data_in[5] ,
    \sw_214_module_data_in[4] ,
    \sw_214_module_data_in[3] ,
    \sw_214_module_data_in[2] ,
    \sw_214_module_data_in[1] ,
    \sw_214_module_data_in[0] }),
    .module_data_out({\sw_214_module_data_out[7] ,
    \sw_214_module_data_out[6] ,
    \sw_214_module_data_out[5] ,
    \sw_214_module_data_out[4] ,
    \sw_214_module_data_out[3] ,
    \sw_214_module_data_out[2] ,
    \sw_214_module_data_out[1] ,
    \sw_214_module_data_out[0] }));
 scanchain scanchain_215 (.clk_in(sw_214_clk_out),
    .clk_out(sw_215_clk_out),
    .data_in(sw_214_data_out),
    .data_out(sw_215_data_out),
    .latch_enable_in(sw_214_latch_out),
    .latch_enable_out(sw_215_latch_out),
    .scan_select_in(sw_214_scan_out),
    .scan_select_out(sw_215_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_215_module_data_in[7] ,
    \sw_215_module_data_in[6] ,
    \sw_215_module_data_in[5] ,
    \sw_215_module_data_in[4] ,
    \sw_215_module_data_in[3] ,
    \sw_215_module_data_in[2] ,
    \sw_215_module_data_in[1] ,
    \sw_215_module_data_in[0] }),
    .module_data_out({\sw_215_module_data_out[7] ,
    \sw_215_module_data_out[6] ,
    \sw_215_module_data_out[5] ,
    \sw_215_module_data_out[4] ,
    \sw_215_module_data_out[3] ,
    \sw_215_module_data_out[2] ,
    \sw_215_module_data_out[1] ,
    \sw_215_module_data_out[0] }));
 scanchain scanchain_216 (.clk_in(sw_215_clk_out),
    .clk_out(sw_216_clk_out),
    .data_in(sw_215_data_out),
    .data_out(sw_216_data_out),
    .latch_enable_in(sw_215_latch_out),
    .latch_enable_out(sw_216_latch_out),
    .scan_select_in(sw_215_scan_out),
    .scan_select_out(sw_216_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_216_module_data_in[7] ,
    \sw_216_module_data_in[6] ,
    \sw_216_module_data_in[5] ,
    \sw_216_module_data_in[4] ,
    \sw_216_module_data_in[3] ,
    \sw_216_module_data_in[2] ,
    \sw_216_module_data_in[1] ,
    \sw_216_module_data_in[0] }),
    .module_data_out({\sw_216_module_data_out[7] ,
    \sw_216_module_data_out[6] ,
    \sw_216_module_data_out[5] ,
    \sw_216_module_data_out[4] ,
    \sw_216_module_data_out[3] ,
    \sw_216_module_data_out[2] ,
    \sw_216_module_data_out[1] ,
    \sw_216_module_data_out[0] }));
 scanchain scanchain_217 (.clk_in(sw_216_clk_out),
    .clk_out(sw_217_clk_out),
    .data_in(sw_216_data_out),
    .data_out(sw_217_data_out),
    .latch_enable_in(sw_216_latch_out),
    .latch_enable_out(sw_217_latch_out),
    .scan_select_in(sw_216_scan_out),
    .scan_select_out(sw_217_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_217_module_data_in[7] ,
    \sw_217_module_data_in[6] ,
    \sw_217_module_data_in[5] ,
    \sw_217_module_data_in[4] ,
    \sw_217_module_data_in[3] ,
    \sw_217_module_data_in[2] ,
    \sw_217_module_data_in[1] ,
    \sw_217_module_data_in[0] }),
    .module_data_out({\sw_217_module_data_out[7] ,
    \sw_217_module_data_out[6] ,
    \sw_217_module_data_out[5] ,
    \sw_217_module_data_out[4] ,
    \sw_217_module_data_out[3] ,
    \sw_217_module_data_out[2] ,
    \sw_217_module_data_out[1] ,
    \sw_217_module_data_out[0] }));
 scanchain scanchain_218 (.clk_in(sw_217_clk_out),
    .clk_out(sw_218_clk_out),
    .data_in(sw_217_data_out),
    .data_out(sw_218_data_out),
    .latch_enable_in(sw_217_latch_out),
    .latch_enable_out(sw_218_latch_out),
    .scan_select_in(sw_217_scan_out),
    .scan_select_out(sw_218_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_218_module_data_in[7] ,
    \sw_218_module_data_in[6] ,
    \sw_218_module_data_in[5] ,
    \sw_218_module_data_in[4] ,
    \sw_218_module_data_in[3] ,
    \sw_218_module_data_in[2] ,
    \sw_218_module_data_in[1] ,
    \sw_218_module_data_in[0] }),
    .module_data_out({\sw_218_module_data_out[7] ,
    \sw_218_module_data_out[6] ,
    \sw_218_module_data_out[5] ,
    \sw_218_module_data_out[4] ,
    \sw_218_module_data_out[3] ,
    \sw_218_module_data_out[2] ,
    \sw_218_module_data_out[1] ,
    \sw_218_module_data_out[0] }));
 scanchain scanchain_219 (.clk_in(sw_218_clk_out),
    .clk_out(sw_219_clk_out),
    .data_in(sw_218_data_out),
    .data_out(sw_219_data_out),
    .latch_enable_in(sw_218_latch_out),
    .latch_enable_out(sw_219_latch_out),
    .scan_select_in(sw_218_scan_out),
    .scan_select_out(sw_219_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_219_module_data_in[7] ,
    \sw_219_module_data_in[6] ,
    \sw_219_module_data_in[5] ,
    \sw_219_module_data_in[4] ,
    \sw_219_module_data_in[3] ,
    \sw_219_module_data_in[2] ,
    \sw_219_module_data_in[1] ,
    \sw_219_module_data_in[0] }),
    .module_data_out({\sw_219_module_data_out[7] ,
    \sw_219_module_data_out[6] ,
    \sw_219_module_data_out[5] ,
    \sw_219_module_data_out[4] ,
    \sw_219_module_data_out[3] ,
    \sw_219_module_data_out[2] ,
    \sw_219_module_data_out[1] ,
    \sw_219_module_data_out[0] }));
 scanchain scanchain_22 (.clk_in(sw_021_clk_out),
    .clk_out(sw_022_clk_out),
    .data_in(sw_021_data_out),
    .data_out(sw_022_data_out),
    .latch_enable_in(sw_021_latch_out),
    .latch_enable_out(sw_022_latch_out),
    .scan_select_in(sw_021_scan_out),
    .scan_select_out(sw_022_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_022_module_data_in[7] ,
    \sw_022_module_data_in[6] ,
    \sw_022_module_data_in[5] ,
    \sw_022_module_data_in[4] ,
    \sw_022_module_data_in[3] ,
    \sw_022_module_data_in[2] ,
    \sw_022_module_data_in[1] ,
    \sw_022_module_data_in[0] }),
    .module_data_out({\sw_022_module_data_out[7] ,
    \sw_022_module_data_out[6] ,
    \sw_022_module_data_out[5] ,
    \sw_022_module_data_out[4] ,
    \sw_022_module_data_out[3] ,
    \sw_022_module_data_out[2] ,
    \sw_022_module_data_out[1] ,
    \sw_022_module_data_out[0] }));
 scanchain scanchain_220 (.clk_in(sw_219_clk_out),
    .clk_out(sw_220_clk_out),
    .data_in(sw_219_data_out),
    .data_out(sw_220_data_out),
    .latch_enable_in(sw_219_latch_out),
    .latch_enable_out(sw_220_latch_out),
    .scan_select_in(sw_219_scan_out),
    .scan_select_out(sw_220_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_220_module_data_in[7] ,
    \sw_220_module_data_in[6] ,
    \sw_220_module_data_in[5] ,
    \sw_220_module_data_in[4] ,
    \sw_220_module_data_in[3] ,
    \sw_220_module_data_in[2] ,
    \sw_220_module_data_in[1] ,
    \sw_220_module_data_in[0] }),
    .module_data_out({\sw_220_module_data_out[7] ,
    \sw_220_module_data_out[6] ,
    \sw_220_module_data_out[5] ,
    \sw_220_module_data_out[4] ,
    \sw_220_module_data_out[3] ,
    \sw_220_module_data_out[2] ,
    \sw_220_module_data_out[1] ,
    \sw_220_module_data_out[0] }));
 scanchain scanchain_221 (.clk_in(sw_220_clk_out),
    .clk_out(sw_221_clk_out),
    .data_in(sw_220_data_out),
    .data_out(sw_221_data_out),
    .latch_enable_in(sw_220_latch_out),
    .latch_enable_out(sw_221_latch_out),
    .scan_select_in(sw_220_scan_out),
    .scan_select_out(sw_221_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_221_module_data_in[7] ,
    \sw_221_module_data_in[6] ,
    \sw_221_module_data_in[5] ,
    \sw_221_module_data_in[4] ,
    \sw_221_module_data_in[3] ,
    \sw_221_module_data_in[2] ,
    \sw_221_module_data_in[1] ,
    \sw_221_module_data_in[0] }),
    .module_data_out({\sw_221_module_data_out[7] ,
    \sw_221_module_data_out[6] ,
    \sw_221_module_data_out[5] ,
    \sw_221_module_data_out[4] ,
    \sw_221_module_data_out[3] ,
    \sw_221_module_data_out[2] ,
    \sw_221_module_data_out[1] ,
    \sw_221_module_data_out[0] }));
 scanchain scanchain_222 (.clk_in(sw_221_clk_out),
    .clk_out(sw_222_clk_out),
    .data_in(sw_221_data_out),
    .data_out(sw_222_data_out),
    .latch_enable_in(sw_221_latch_out),
    .latch_enable_out(sw_222_latch_out),
    .scan_select_in(sw_221_scan_out),
    .scan_select_out(sw_222_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_222_module_data_in[7] ,
    \sw_222_module_data_in[6] ,
    \sw_222_module_data_in[5] ,
    \sw_222_module_data_in[4] ,
    \sw_222_module_data_in[3] ,
    \sw_222_module_data_in[2] ,
    \sw_222_module_data_in[1] ,
    \sw_222_module_data_in[0] }),
    .module_data_out({\sw_222_module_data_out[7] ,
    \sw_222_module_data_out[6] ,
    \sw_222_module_data_out[5] ,
    \sw_222_module_data_out[4] ,
    \sw_222_module_data_out[3] ,
    \sw_222_module_data_out[2] ,
    \sw_222_module_data_out[1] ,
    \sw_222_module_data_out[0] }));
 scanchain scanchain_223 (.clk_in(sw_222_clk_out),
    .clk_out(sw_223_clk_out),
    .data_in(sw_222_data_out),
    .data_out(sw_223_data_out),
    .latch_enable_in(sw_222_latch_out),
    .latch_enable_out(sw_223_latch_out),
    .scan_select_in(sw_222_scan_out),
    .scan_select_out(sw_223_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_223_module_data_in[7] ,
    \sw_223_module_data_in[6] ,
    \sw_223_module_data_in[5] ,
    \sw_223_module_data_in[4] ,
    \sw_223_module_data_in[3] ,
    \sw_223_module_data_in[2] ,
    \sw_223_module_data_in[1] ,
    \sw_223_module_data_in[0] }),
    .module_data_out({\sw_223_module_data_out[7] ,
    \sw_223_module_data_out[6] ,
    \sw_223_module_data_out[5] ,
    \sw_223_module_data_out[4] ,
    \sw_223_module_data_out[3] ,
    \sw_223_module_data_out[2] ,
    \sw_223_module_data_out[1] ,
    \sw_223_module_data_out[0] }));
 scanchain scanchain_224 (.clk_in(sw_223_clk_out),
    .clk_out(sw_224_clk_out),
    .data_in(sw_223_data_out),
    .data_out(sw_224_data_out),
    .latch_enable_in(sw_223_latch_out),
    .latch_enable_out(sw_224_latch_out),
    .scan_select_in(sw_223_scan_out),
    .scan_select_out(sw_224_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_224_module_data_in[7] ,
    \sw_224_module_data_in[6] ,
    \sw_224_module_data_in[5] ,
    \sw_224_module_data_in[4] ,
    \sw_224_module_data_in[3] ,
    \sw_224_module_data_in[2] ,
    \sw_224_module_data_in[1] ,
    \sw_224_module_data_in[0] }),
    .module_data_out({\sw_224_module_data_out[7] ,
    \sw_224_module_data_out[6] ,
    \sw_224_module_data_out[5] ,
    \sw_224_module_data_out[4] ,
    \sw_224_module_data_out[3] ,
    \sw_224_module_data_out[2] ,
    \sw_224_module_data_out[1] ,
    \sw_224_module_data_out[0] }));
 scanchain scanchain_225 (.clk_in(sw_224_clk_out),
    .clk_out(sw_225_clk_out),
    .data_in(sw_224_data_out),
    .data_out(sw_225_data_out),
    .latch_enable_in(sw_224_latch_out),
    .latch_enable_out(sw_225_latch_out),
    .scan_select_in(sw_224_scan_out),
    .scan_select_out(sw_225_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_225_module_data_in[7] ,
    \sw_225_module_data_in[6] ,
    \sw_225_module_data_in[5] ,
    \sw_225_module_data_in[4] ,
    \sw_225_module_data_in[3] ,
    \sw_225_module_data_in[2] ,
    \sw_225_module_data_in[1] ,
    \sw_225_module_data_in[0] }),
    .module_data_out({\sw_225_module_data_out[7] ,
    \sw_225_module_data_out[6] ,
    \sw_225_module_data_out[5] ,
    \sw_225_module_data_out[4] ,
    \sw_225_module_data_out[3] ,
    \sw_225_module_data_out[2] ,
    \sw_225_module_data_out[1] ,
    \sw_225_module_data_out[0] }));
 scanchain scanchain_226 (.clk_in(sw_225_clk_out),
    .clk_out(sw_226_clk_out),
    .data_in(sw_225_data_out),
    .data_out(sw_226_data_out),
    .latch_enable_in(sw_225_latch_out),
    .latch_enable_out(sw_226_latch_out),
    .scan_select_in(sw_225_scan_out),
    .scan_select_out(sw_226_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_226_module_data_in[7] ,
    \sw_226_module_data_in[6] ,
    \sw_226_module_data_in[5] ,
    \sw_226_module_data_in[4] ,
    \sw_226_module_data_in[3] ,
    \sw_226_module_data_in[2] ,
    \sw_226_module_data_in[1] ,
    \sw_226_module_data_in[0] }),
    .module_data_out({\sw_226_module_data_out[7] ,
    \sw_226_module_data_out[6] ,
    \sw_226_module_data_out[5] ,
    \sw_226_module_data_out[4] ,
    \sw_226_module_data_out[3] ,
    \sw_226_module_data_out[2] ,
    \sw_226_module_data_out[1] ,
    \sw_226_module_data_out[0] }));
 scanchain scanchain_227 (.clk_in(sw_226_clk_out),
    .clk_out(sw_227_clk_out),
    .data_in(sw_226_data_out),
    .data_out(sw_227_data_out),
    .latch_enable_in(sw_226_latch_out),
    .latch_enable_out(sw_227_latch_out),
    .scan_select_in(sw_226_scan_out),
    .scan_select_out(sw_227_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_227_module_data_in[7] ,
    \sw_227_module_data_in[6] ,
    \sw_227_module_data_in[5] ,
    \sw_227_module_data_in[4] ,
    \sw_227_module_data_in[3] ,
    \sw_227_module_data_in[2] ,
    \sw_227_module_data_in[1] ,
    \sw_227_module_data_in[0] }),
    .module_data_out({\sw_227_module_data_out[7] ,
    \sw_227_module_data_out[6] ,
    \sw_227_module_data_out[5] ,
    \sw_227_module_data_out[4] ,
    \sw_227_module_data_out[3] ,
    \sw_227_module_data_out[2] ,
    \sw_227_module_data_out[1] ,
    \sw_227_module_data_out[0] }));
 scanchain scanchain_228 (.clk_in(sw_227_clk_out),
    .clk_out(sw_228_clk_out),
    .data_in(sw_227_data_out),
    .data_out(sw_228_data_out),
    .latch_enable_in(sw_227_latch_out),
    .latch_enable_out(sw_228_latch_out),
    .scan_select_in(sw_227_scan_out),
    .scan_select_out(sw_228_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_228_module_data_in[7] ,
    \sw_228_module_data_in[6] ,
    \sw_228_module_data_in[5] ,
    \sw_228_module_data_in[4] ,
    \sw_228_module_data_in[3] ,
    \sw_228_module_data_in[2] ,
    \sw_228_module_data_in[1] ,
    \sw_228_module_data_in[0] }),
    .module_data_out({\sw_228_module_data_out[7] ,
    \sw_228_module_data_out[6] ,
    \sw_228_module_data_out[5] ,
    \sw_228_module_data_out[4] ,
    \sw_228_module_data_out[3] ,
    \sw_228_module_data_out[2] ,
    \sw_228_module_data_out[1] ,
    \sw_228_module_data_out[0] }));
 scanchain scanchain_229 (.clk_in(sw_228_clk_out),
    .clk_out(sw_229_clk_out),
    .data_in(sw_228_data_out),
    .data_out(sw_229_data_out),
    .latch_enable_in(sw_228_latch_out),
    .latch_enable_out(sw_229_latch_out),
    .scan_select_in(sw_228_scan_out),
    .scan_select_out(sw_229_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_229_module_data_in[7] ,
    \sw_229_module_data_in[6] ,
    \sw_229_module_data_in[5] ,
    \sw_229_module_data_in[4] ,
    \sw_229_module_data_in[3] ,
    \sw_229_module_data_in[2] ,
    \sw_229_module_data_in[1] ,
    \sw_229_module_data_in[0] }),
    .module_data_out({\sw_229_module_data_out[7] ,
    \sw_229_module_data_out[6] ,
    \sw_229_module_data_out[5] ,
    \sw_229_module_data_out[4] ,
    \sw_229_module_data_out[3] ,
    \sw_229_module_data_out[2] ,
    \sw_229_module_data_out[1] ,
    \sw_229_module_data_out[0] }));
 scanchain scanchain_23 (.clk_in(sw_022_clk_out),
    .clk_out(sw_023_clk_out),
    .data_in(sw_022_data_out),
    .data_out(sw_023_data_out),
    .latch_enable_in(sw_022_latch_out),
    .latch_enable_out(sw_023_latch_out),
    .scan_select_in(sw_022_scan_out),
    .scan_select_out(sw_023_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_023_module_data_in[7] ,
    \sw_023_module_data_in[6] ,
    \sw_023_module_data_in[5] ,
    \sw_023_module_data_in[4] ,
    \sw_023_module_data_in[3] ,
    \sw_023_module_data_in[2] ,
    \sw_023_module_data_in[1] ,
    \sw_023_module_data_in[0] }),
    .module_data_out({\sw_023_module_data_out[7] ,
    \sw_023_module_data_out[6] ,
    \sw_023_module_data_out[5] ,
    \sw_023_module_data_out[4] ,
    \sw_023_module_data_out[3] ,
    \sw_023_module_data_out[2] ,
    \sw_023_module_data_out[1] ,
    \sw_023_module_data_out[0] }));
 scanchain scanchain_230 (.clk_in(sw_229_clk_out),
    .clk_out(sw_230_clk_out),
    .data_in(sw_229_data_out),
    .data_out(sw_230_data_out),
    .latch_enable_in(sw_229_latch_out),
    .latch_enable_out(sw_230_latch_out),
    .scan_select_in(sw_229_scan_out),
    .scan_select_out(sw_230_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_230_module_data_in[7] ,
    \sw_230_module_data_in[6] ,
    \sw_230_module_data_in[5] ,
    \sw_230_module_data_in[4] ,
    \sw_230_module_data_in[3] ,
    \sw_230_module_data_in[2] ,
    \sw_230_module_data_in[1] ,
    \sw_230_module_data_in[0] }),
    .module_data_out({\sw_230_module_data_out[7] ,
    \sw_230_module_data_out[6] ,
    \sw_230_module_data_out[5] ,
    \sw_230_module_data_out[4] ,
    \sw_230_module_data_out[3] ,
    \sw_230_module_data_out[2] ,
    \sw_230_module_data_out[1] ,
    \sw_230_module_data_out[0] }));
 scanchain scanchain_231 (.clk_in(sw_230_clk_out),
    .clk_out(sw_231_clk_out),
    .data_in(sw_230_data_out),
    .data_out(sw_231_data_out),
    .latch_enable_in(sw_230_latch_out),
    .latch_enable_out(sw_231_latch_out),
    .scan_select_in(sw_230_scan_out),
    .scan_select_out(sw_231_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_231_module_data_in[7] ,
    \sw_231_module_data_in[6] ,
    \sw_231_module_data_in[5] ,
    \sw_231_module_data_in[4] ,
    \sw_231_module_data_in[3] ,
    \sw_231_module_data_in[2] ,
    \sw_231_module_data_in[1] ,
    \sw_231_module_data_in[0] }),
    .module_data_out({\sw_231_module_data_out[7] ,
    \sw_231_module_data_out[6] ,
    \sw_231_module_data_out[5] ,
    \sw_231_module_data_out[4] ,
    \sw_231_module_data_out[3] ,
    \sw_231_module_data_out[2] ,
    \sw_231_module_data_out[1] ,
    \sw_231_module_data_out[0] }));
 scanchain scanchain_232 (.clk_in(sw_231_clk_out),
    .clk_out(sw_232_clk_out),
    .data_in(sw_231_data_out),
    .data_out(sw_232_data_out),
    .latch_enable_in(sw_231_latch_out),
    .latch_enable_out(sw_232_latch_out),
    .scan_select_in(sw_231_scan_out),
    .scan_select_out(sw_232_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_232_module_data_in[7] ,
    \sw_232_module_data_in[6] ,
    \sw_232_module_data_in[5] ,
    \sw_232_module_data_in[4] ,
    \sw_232_module_data_in[3] ,
    \sw_232_module_data_in[2] ,
    \sw_232_module_data_in[1] ,
    \sw_232_module_data_in[0] }),
    .module_data_out({\sw_232_module_data_out[7] ,
    \sw_232_module_data_out[6] ,
    \sw_232_module_data_out[5] ,
    \sw_232_module_data_out[4] ,
    \sw_232_module_data_out[3] ,
    \sw_232_module_data_out[2] ,
    \sw_232_module_data_out[1] ,
    \sw_232_module_data_out[0] }));
 scanchain scanchain_233 (.clk_in(sw_232_clk_out),
    .clk_out(sw_233_clk_out),
    .data_in(sw_232_data_out),
    .data_out(sw_233_data_out),
    .latch_enable_in(sw_232_latch_out),
    .latch_enable_out(sw_233_latch_out),
    .scan_select_in(sw_232_scan_out),
    .scan_select_out(sw_233_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_233_module_data_in[7] ,
    \sw_233_module_data_in[6] ,
    \sw_233_module_data_in[5] ,
    \sw_233_module_data_in[4] ,
    \sw_233_module_data_in[3] ,
    \sw_233_module_data_in[2] ,
    \sw_233_module_data_in[1] ,
    \sw_233_module_data_in[0] }),
    .module_data_out({\sw_233_module_data_out[7] ,
    \sw_233_module_data_out[6] ,
    \sw_233_module_data_out[5] ,
    \sw_233_module_data_out[4] ,
    \sw_233_module_data_out[3] ,
    \sw_233_module_data_out[2] ,
    \sw_233_module_data_out[1] ,
    \sw_233_module_data_out[0] }));
 scanchain scanchain_234 (.clk_in(sw_233_clk_out),
    .clk_out(sw_234_clk_out),
    .data_in(sw_233_data_out),
    .data_out(sw_234_data_out),
    .latch_enable_in(sw_233_latch_out),
    .latch_enable_out(sw_234_latch_out),
    .scan_select_in(sw_233_scan_out),
    .scan_select_out(sw_234_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_234_module_data_in[7] ,
    \sw_234_module_data_in[6] ,
    \sw_234_module_data_in[5] ,
    \sw_234_module_data_in[4] ,
    \sw_234_module_data_in[3] ,
    \sw_234_module_data_in[2] ,
    \sw_234_module_data_in[1] ,
    \sw_234_module_data_in[0] }),
    .module_data_out({\sw_234_module_data_out[7] ,
    \sw_234_module_data_out[6] ,
    \sw_234_module_data_out[5] ,
    \sw_234_module_data_out[4] ,
    \sw_234_module_data_out[3] ,
    \sw_234_module_data_out[2] ,
    \sw_234_module_data_out[1] ,
    \sw_234_module_data_out[0] }));
 scanchain scanchain_235 (.clk_in(sw_234_clk_out),
    .clk_out(sw_235_clk_out),
    .data_in(sw_234_data_out),
    .data_out(sw_235_data_out),
    .latch_enable_in(sw_234_latch_out),
    .latch_enable_out(sw_235_latch_out),
    .scan_select_in(sw_234_scan_out),
    .scan_select_out(sw_235_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_235_module_data_in[7] ,
    \sw_235_module_data_in[6] ,
    \sw_235_module_data_in[5] ,
    \sw_235_module_data_in[4] ,
    \sw_235_module_data_in[3] ,
    \sw_235_module_data_in[2] ,
    \sw_235_module_data_in[1] ,
    \sw_235_module_data_in[0] }),
    .module_data_out({\sw_235_module_data_out[7] ,
    \sw_235_module_data_out[6] ,
    \sw_235_module_data_out[5] ,
    \sw_235_module_data_out[4] ,
    \sw_235_module_data_out[3] ,
    \sw_235_module_data_out[2] ,
    \sw_235_module_data_out[1] ,
    \sw_235_module_data_out[0] }));
 scanchain scanchain_236 (.clk_in(sw_235_clk_out),
    .clk_out(sw_236_clk_out),
    .data_in(sw_235_data_out),
    .data_out(sw_236_data_out),
    .latch_enable_in(sw_235_latch_out),
    .latch_enable_out(sw_236_latch_out),
    .scan_select_in(sw_235_scan_out),
    .scan_select_out(sw_236_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_236_module_data_in[7] ,
    \sw_236_module_data_in[6] ,
    \sw_236_module_data_in[5] ,
    \sw_236_module_data_in[4] ,
    \sw_236_module_data_in[3] ,
    \sw_236_module_data_in[2] ,
    \sw_236_module_data_in[1] ,
    \sw_236_module_data_in[0] }),
    .module_data_out({\sw_236_module_data_out[7] ,
    \sw_236_module_data_out[6] ,
    \sw_236_module_data_out[5] ,
    \sw_236_module_data_out[4] ,
    \sw_236_module_data_out[3] ,
    \sw_236_module_data_out[2] ,
    \sw_236_module_data_out[1] ,
    \sw_236_module_data_out[0] }));
 scanchain scanchain_237 (.clk_in(sw_236_clk_out),
    .clk_out(sw_237_clk_out),
    .data_in(sw_236_data_out),
    .data_out(sw_237_data_out),
    .latch_enable_in(sw_236_latch_out),
    .latch_enable_out(sw_237_latch_out),
    .scan_select_in(sw_236_scan_out),
    .scan_select_out(sw_237_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_237_module_data_in[7] ,
    \sw_237_module_data_in[6] ,
    \sw_237_module_data_in[5] ,
    \sw_237_module_data_in[4] ,
    \sw_237_module_data_in[3] ,
    \sw_237_module_data_in[2] ,
    \sw_237_module_data_in[1] ,
    \sw_237_module_data_in[0] }),
    .module_data_out({\sw_237_module_data_out[7] ,
    \sw_237_module_data_out[6] ,
    \sw_237_module_data_out[5] ,
    \sw_237_module_data_out[4] ,
    \sw_237_module_data_out[3] ,
    \sw_237_module_data_out[2] ,
    \sw_237_module_data_out[1] ,
    \sw_237_module_data_out[0] }));
 scanchain scanchain_238 (.clk_in(sw_237_clk_out),
    .clk_out(sw_238_clk_out),
    .data_in(sw_237_data_out),
    .data_out(sw_238_data_out),
    .latch_enable_in(sw_237_latch_out),
    .latch_enable_out(sw_238_latch_out),
    .scan_select_in(sw_237_scan_out),
    .scan_select_out(sw_238_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_238_module_data_in[7] ,
    \sw_238_module_data_in[6] ,
    \sw_238_module_data_in[5] ,
    \sw_238_module_data_in[4] ,
    \sw_238_module_data_in[3] ,
    \sw_238_module_data_in[2] ,
    \sw_238_module_data_in[1] ,
    \sw_238_module_data_in[0] }),
    .module_data_out({\sw_238_module_data_out[7] ,
    \sw_238_module_data_out[6] ,
    \sw_238_module_data_out[5] ,
    \sw_238_module_data_out[4] ,
    \sw_238_module_data_out[3] ,
    \sw_238_module_data_out[2] ,
    \sw_238_module_data_out[1] ,
    \sw_238_module_data_out[0] }));
 scanchain scanchain_239 (.clk_in(sw_238_clk_out),
    .clk_out(sw_239_clk_out),
    .data_in(sw_238_data_out),
    .data_out(sw_239_data_out),
    .latch_enable_in(sw_238_latch_out),
    .latch_enable_out(sw_239_latch_out),
    .scan_select_in(sw_238_scan_out),
    .scan_select_out(sw_239_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_239_module_data_in[7] ,
    \sw_239_module_data_in[6] ,
    \sw_239_module_data_in[5] ,
    \sw_239_module_data_in[4] ,
    \sw_239_module_data_in[3] ,
    \sw_239_module_data_in[2] ,
    \sw_239_module_data_in[1] ,
    \sw_239_module_data_in[0] }),
    .module_data_out({\sw_239_module_data_out[7] ,
    \sw_239_module_data_out[6] ,
    \sw_239_module_data_out[5] ,
    \sw_239_module_data_out[4] ,
    \sw_239_module_data_out[3] ,
    \sw_239_module_data_out[2] ,
    \sw_239_module_data_out[1] ,
    \sw_239_module_data_out[0] }));
 scanchain scanchain_24 (.clk_in(sw_023_clk_out),
    .clk_out(sw_024_clk_out),
    .data_in(sw_023_data_out),
    .data_out(sw_024_data_out),
    .latch_enable_in(sw_023_latch_out),
    .latch_enable_out(sw_024_latch_out),
    .scan_select_in(sw_023_scan_out),
    .scan_select_out(sw_024_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_024_module_data_in[7] ,
    \sw_024_module_data_in[6] ,
    \sw_024_module_data_in[5] ,
    \sw_024_module_data_in[4] ,
    \sw_024_module_data_in[3] ,
    \sw_024_module_data_in[2] ,
    \sw_024_module_data_in[1] ,
    \sw_024_module_data_in[0] }),
    .module_data_out({\sw_024_module_data_out[7] ,
    \sw_024_module_data_out[6] ,
    \sw_024_module_data_out[5] ,
    \sw_024_module_data_out[4] ,
    \sw_024_module_data_out[3] ,
    \sw_024_module_data_out[2] ,
    \sw_024_module_data_out[1] ,
    \sw_024_module_data_out[0] }));
 scanchain scanchain_240 (.clk_in(sw_239_clk_out),
    .clk_out(sw_240_clk_out),
    .data_in(sw_239_data_out),
    .data_out(sw_240_data_out),
    .latch_enable_in(sw_239_latch_out),
    .latch_enable_out(sw_240_latch_out),
    .scan_select_in(sw_239_scan_out),
    .scan_select_out(sw_240_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_240_module_data_in[7] ,
    \sw_240_module_data_in[6] ,
    \sw_240_module_data_in[5] ,
    \sw_240_module_data_in[4] ,
    \sw_240_module_data_in[3] ,
    \sw_240_module_data_in[2] ,
    \sw_240_module_data_in[1] ,
    \sw_240_module_data_in[0] }),
    .module_data_out({\sw_240_module_data_out[7] ,
    \sw_240_module_data_out[6] ,
    \sw_240_module_data_out[5] ,
    \sw_240_module_data_out[4] ,
    \sw_240_module_data_out[3] ,
    \sw_240_module_data_out[2] ,
    \sw_240_module_data_out[1] ,
    \sw_240_module_data_out[0] }));
 scanchain scanchain_241 (.clk_in(sw_240_clk_out),
    .clk_out(sw_241_clk_out),
    .data_in(sw_240_data_out),
    .data_out(sw_241_data_out),
    .latch_enable_in(sw_240_latch_out),
    .latch_enable_out(sw_241_latch_out),
    .scan_select_in(sw_240_scan_out),
    .scan_select_out(sw_241_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_241_module_data_in[7] ,
    \sw_241_module_data_in[6] ,
    \sw_241_module_data_in[5] ,
    \sw_241_module_data_in[4] ,
    \sw_241_module_data_in[3] ,
    \sw_241_module_data_in[2] ,
    \sw_241_module_data_in[1] ,
    \sw_241_module_data_in[0] }),
    .module_data_out({\sw_241_module_data_out[7] ,
    \sw_241_module_data_out[6] ,
    \sw_241_module_data_out[5] ,
    \sw_241_module_data_out[4] ,
    \sw_241_module_data_out[3] ,
    \sw_241_module_data_out[2] ,
    \sw_241_module_data_out[1] ,
    \sw_241_module_data_out[0] }));
 scanchain scanchain_242 (.clk_in(sw_241_clk_out),
    .clk_out(sw_242_clk_out),
    .data_in(sw_241_data_out),
    .data_out(sw_242_data_out),
    .latch_enable_in(sw_241_latch_out),
    .latch_enable_out(sw_242_latch_out),
    .scan_select_in(sw_241_scan_out),
    .scan_select_out(sw_242_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_242_module_data_in[7] ,
    \sw_242_module_data_in[6] ,
    \sw_242_module_data_in[5] ,
    \sw_242_module_data_in[4] ,
    \sw_242_module_data_in[3] ,
    \sw_242_module_data_in[2] ,
    \sw_242_module_data_in[1] ,
    \sw_242_module_data_in[0] }),
    .module_data_out({\sw_242_module_data_out[7] ,
    \sw_242_module_data_out[6] ,
    \sw_242_module_data_out[5] ,
    \sw_242_module_data_out[4] ,
    \sw_242_module_data_out[3] ,
    \sw_242_module_data_out[2] ,
    \sw_242_module_data_out[1] ,
    \sw_242_module_data_out[0] }));
 scanchain scanchain_243 (.clk_in(sw_242_clk_out),
    .clk_out(sw_243_clk_out),
    .data_in(sw_242_data_out),
    .data_out(sw_243_data_out),
    .latch_enable_in(sw_242_latch_out),
    .latch_enable_out(sw_243_latch_out),
    .scan_select_in(sw_242_scan_out),
    .scan_select_out(sw_243_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_243_module_data_in[7] ,
    \sw_243_module_data_in[6] ,
    \sw_243_module_data_in[5] ,
    \sw_243_module_data_in[4] ,
    \sw_243_module_data_in[3] ,
    \sw_243_module_data_in[2] ,
    \sw_243_module_data_in[1] ,
    \sw_243_module_data_in[0] }),
    .module_data_out({\sw_243_module_data_out[7] ,
    \sw_243_module_data_out[6] ,
    \sw_243_module_data_out[5] ,
    \sw_243_module_data_out[4] ,
    \sw_243_module_data_out[3] ,
    \sw_243_module_data_out[2] ,
    \sw_243_module_data_out[1] ,
    \sw_243_module_data_out[0] }));
 scanchain scanchain_244 (.clk_in(sw_243_clk_out),
    .clk_out(sw_244_clk_out),
    .data_in(sw_243_data_out),
    .data_out(sw_244_data_out),
    .latch_enable_in(sw_243_latch_out),
    .latch_enable_out(sw_244_latch_out),
    .scan_select_in(sw_243_scan_out),
    .scan_select_out(sw_244_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_244_module_data_in[7] ,
    \sw_244_module_data_in[6] ,
    \sw_244_module_data_in[5] ,
    \sw_244_module_data_in[4] ,
    \sw_244_module_data_in[3] ,
    \sw_244_module_data_in[2] ,
    \sw_244_module_data_in[1] ,
    \sw_244_module_data_in[0] }),
    .module_data_out({\sw_244_module_data_out[7] ,
    \sw_244_module_data_out[6] ,
    \sw_244_module_data_out[5] ,
    \sw_244_module_data_out[4] ,
    \sw_244_module_data_out[3] ,
    \sw_244_module_data_out[2] ,
    \sw_244_module_data_out[1] ,
    \sw_244_module_data_out[0] }));
 scanchain scanchain_245 (.clk_in(sw_244_clk_out),
    .clk_out(sw_245_clk_out),
    .data_in(sw_244_data_out),
    .data_out(sw_245_data_out),
    .latch_enable_in(sw_244_latch_out),
    .latch_enable_out(sw_245_latch_out),
    .scan_select_in(sw_244_scan_out),
    .scan_select_out(sw_245_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_245_module_data_in[7] ,
    \sw_245_module_data_in[6] ,
    \sw_245_module_data_in[5] ,
    \sw_245_module_data_in[4] ,
    \sw_245_module_data_in[3] ,
    \sw_245_module_data_in[2] ,
    \sw_245_module_data_in[1] ,
    \sw_245_module_data_in[0] }),
    .module_data_out({\sw_245_module_data_out[7] ,
    \sw_245_module_data_out[6] ,
    \sw_245_module_data_out[5] ,
    \sw_245_module_data_out[4] ,
    \sw_245_module_data_out[3] ,
    \sw_245_module_data_out[2] ,
    \sw_245_module_data_out[1] ,
    \sw_245_module_data_out[0] }));
 scanchain scanchain_246 (.clk_in(sw_245_clk_out),
    .clk_out(sw_246_clk_out),
    .data_in(sw_245_data_out),
    .data_out(sw_246_data_out),
    .latch_enable_in(sw_245_latch_out),
    .latch_enable_out(sw_246_latch_out),
    .scan_select_in(sw_245_scan_out),
    .scan_select_out(sw_246_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_246_module_data_in[7] ,
    \sw_246_module_data_in[6] ,
    \sw_246_module_data_in[5] ,
    \sw_246_module_data_in[4] ,
    \sw_246_module_data_in[3] ,
    \sw_246_module_data_in[2] ,
    \sw_246_module_data_in[1] ,
    \sw_246_module_data_in[0] }),
    .module_data_out({\sw_246_module_data_out[7] ,
    \sw_246_module_data_out[6] ,
    \sw_246_module_data_out[5] ,
    \sw_246_module_data_out[4] ,
    \sw_246_module_data_out[3] ,
    \sw_246_module_data_out[2] ,
    \sw_246_module_data_out[1] ,
    \sw_246_module_data_out[0] }));
 scanchain scanchain_247 (.clk_in(sw_246_clk_out),
    .clk_out(sw_247_clk_out),
    .data_in(sw_246_data_out),
    .data_out(sw_247_data_out),
    .latch_enable_in(sw_246_latch_out),
    .latch_enable_out(sw_247_latch_out),
    .scan_select_in(sw_246_scan_out),
    .scan_select_out(sw_247_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_247_module_data_in[7] ,
    \sw_247_module_data_in[6] ,
    \sw_247_module_data_in[5] ,
    \sw_247_module_data_in[4] ,
    \sw_247_module_data_in[3] ,
    \sw_247_module_data_in[2] ,
    \sw_247_module_data_in[1] ,
    \sw_247_module_data_in[0] }),
    .module_data_out({\sw_247_module_data_out[7] ,
    \sw_247_module_data_out[6] ,
    \sw_247_module_data_out[5] ,
    \sw_247_module_data_out[4] ,
    \sw_247_module_data_out[3] ,
    \sw_247_module_data_out[2] ,
    \sw_247_module_data_out[1] ,
    \sw_247_module_data_out[0] }));
 scanchain scanchain_248 (.clk_in(sw_247_clk_out),
    .clk_out(sw_248_clk_out),
    .data_in(sw_247_data_out),
    .data_out(sw_248_data_out),
    .latch_enable_in(sw_247_latch_out),
    .latch_enable_out(sw_248_latch_out),
    .scan_select_in(sw_247_scan_out),
    .scan_select_out(sw_248_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_248_module_data_in[7] ,
    \sw_248_module_data_in[6] ,
    \sw_248_module_data_in[5] ,
    \sw_248_module_data_in[4] ,
    \sw_248_module_data_in[3] ,
    \sw_248_module_data_in[2] ,
    \sw_248_module_data_in[1] ,
    \sw_248_module_data_in[0] }),
    .module_data_out({\sw_248_module_data_out[7] ,
    \sw_248_module_data_out[6] ,
    \sw_248_module_data_out[5] ,
    \sw_248_module_data_out[4] ,
    \sw_248_module_data_out[3] ,
    \sw_248_module_data_out[2] ,
    \sw_248_module_data_out[1] ,
    \sw_248_module_data_out[0] }));
 scanchain scanchain_249 (.clk_in(sw_248_clk_out),
    .clk_out(sw_249_clk_out),
    .data_in(sw_248_data_out),
    .data_out(sw_249_data_out),
    .latch_enable_in(sw_248_latch_out),
    .latch_enable_out(sw_249_latch_out),
    .scan_select_in(sw_248_scan_out),
    .scan_select_out(sw_249_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_249_module_data_in[7] ,
    \sw_249_module_data_in[6] ,
    \sw_249_module_data_in[5] ,
    \sw_249_module_data_in[4] ,
    \sw_249_module_data_in[3] ,
    \sw_249_module_data_in[2] ,
    \sw_249_module_data_in[1] ,
    \sw_249_module_data_in[0] }),
    .module_data_out({\sw_249_module_data_out[7] ,
    \sw_249_module_data_out[6] ,
    \sw_249_module_data_out[5] ,
    \sw_249_module_data_out[4] ,
    \sw_249_module_data_out[3] ,
    \sw_249_module_data_out[2] ,
    \sw_249_module_data_out[1] ,
    \sw_249_module_data_out[0] }));
 scanchain scanchain_25 (.clk_in(sw_024_clk_out),
    .clk_out(sw_025_clk_out),
    .data_in(sw_024_data_out),
    .data_out(sw_025_data_out),
    .latch_enable_in(sw_024_latch_out),
    .latch_enable_out(sw_025_latch_out),
    .scan_select_in(sw_024_scan_out),
    .scan_select_out(sw_025_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_025_module_data_in[7] ,
    \sw_025_module_data_in[6] ,
    \sw_025_module_data_in[5] ,
    \sw_025_module_data_in[4] ,
    \sw_025_module_data_in[3] ,
    \sw_025_module_data_in[2] ,
    \sw_025_module_data_in[1] ,
    \sw_025_module_data_in[0] }),
    .module_data_out({\sw_025_module_data_out[7] ,
    \sw_025_module_data_out[6] ,
    \sw_025_module_data_out[5] ,
    \sw_025_module_data_out[4] ,
    \sw_025_module_data_out[3] ,
    \sw_025_module_data_out[2] ,
    \sw_025_module_data_out[1] ,
    \sw_025_module_data_out[0] }));
 scanchain scanchain_250 (.clk_in(sw_249_clk_out),
    .clk_out(sw_250_clk_out),
    .data_in(sw_249_data_out),
    .data_out(sw_250_data_out),
    .latch_enable_in(sw_249_latch_out),
    .latch_enable_out(sw_250_latch_out),
    .scan_select_in(sw_249_scan_out),
    .scan_select_out(sw_250_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_250_module_data_in[7] ,
    \sw_250_module_data_in[6] ,
    \sw_250_module_data_in[5] ,
    \sw_250_module_data_in[4] ,
    \sw_250_module_data_in[3] ,
    \sw_250_module_data_in[2] ,
    \sw_250_module_data_in[1] ,
    \sw_250_module_data_in[0] }),
    .module_data_out({\sw_250_module_data_out[7] ,
    \sw_250_module_data_out[6] ,
    \sw_250_module_data_out[5] ,
    \sw_250_module_data_out[4] ,
    \sw_250_module_data_out[3] ,
    \sw_250_module_data_out[2] ,
    \sw_250_module_data_out[1] ,
    \sw_250_module_data_out[0] }));
 scanchain scanchain_251 (.clk_in(sw_250_clk_out),
    .clk_out(sw_251_clk_out),
    .data_in(sw_250_data_out),
    .data_out(sw_251_data_out),
    .latch_enable_in(sw_250_latch_out),
    .latch_enable_out(sw_251_latch_out),
    .scan_select_in(sw_250_scan_out),
    .scan_select_out(sw_251_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_251_module_data_in[7] ,
    \sw_251_module_data_in[6] ,
    \sw_251_module_data_in[5] ,
    \sw_251_module_data_in[4] ,
    \sw_251_module_data_in[3] ,
    \sw_251_module_data_in[2] ,
    \sw_251_module_data_in[1] ,
    \sw_251_module_data_in[0] }),
    .module_data_out({\sw_251_module_data_out[7] ,
    \sw_251_module_data_out[6] ,
    \sw_251_module_data_out[5] ,
    \sw_251_module_data_out[4] ,
    \sw_251_module_data_out[3] ,
    \sw_251_module_data_out[2] ,
    \sw_251_module_data_out[1] ,
    \sw_251_module_data_out[0] }));
 scanchain scanchain_252 (.clk_in(sw_251_clk_out),
    .clk_out(sw_252_clk_out),
    .data_in(sw_251_data_out),
    .data_out(sw_252_data_out),
    .latch_enable_in(sw_251_latch_out),
    .latch_enable_out(sw_252_latch_out),
    .scan_select_in(sw_251_scan_out),
    .scan_select_out(sw_252_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_252_module_data_in[7] ,
    \sw_252_module_data_in[6] ,
    \sw_252_module_data_in[5] ,
    \sw_252_module_data_in[4] ,
    \sw_252_module_data_in[3] ,
    \sw_252_module_data_in[2] ,
    \sw_252_module_data_in[1] ,
    \sw_252_module_data_in[0] }),
    .module_data_out({\sw_252_module_data_out[7] ,
    \sw_252_module_data_out[6] ,
    \sw_252_module_data_out[5] ,
    \sw_252_module_data_out[4] ,
    \sw_252_module_data_out[3] ,
    \sw_252_module_data_out[2] ,
    \sw_252_module_data_out[1] ,
    \sw_252_module_data_out[0] }));
 scanchain scanchain_253 (.clk_in(sw_252_clk_out),
    .clk_out(sw_253_clk_out),
    .data_in(sw_252_data_out),
    .data_out(sw_253_data_out),
    .latch_enable_in(sw_252_latch_out),
    .latch_enable_out(sw_253_latch_out),
    .scan_select_in(sw_252_scan_out),
    .scan_select_out(sw_253_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_253_module_data_in[7] ,
    \sw_253_module_data_in[6] ,
    \sw_253_module_data_in[5] ,
    \sw_253_module_data_in[4] ,
    \sw_253_module_data_in[3] ,
    \sw_253_module_data_in[2] ,
    \sw_253_module_data_in[1] ,
    \sw_253_module_data_in[0] }),
    .module_data_out({\sw_253_module_data_out[7] ,
    \sw_253_module_data_out[6] ,
    \sw_253_module_data_out[5] ,
    \sw_253_module_data_out[4] ,
    \sw_253_module_data_out[3] ,
    \sw_253_module_data_out[2] ,
    \sw_253_module_data_out[1] ,
    \sw_253_module_data_out[0] }));
 scanchain scanchain_254 (.clk_in(sw_253_clk_out),
    .clk_out(sw_254_clk_out),
    .data_in(sw_253_data_out),
    .data_out(sw_254_data_out),
    .latch_enable_in(sw_253_latch_out),
    .latch_enable_out(sw_254_latch_out),
    .scan_select_in(sw_253_scan_out),
    .scan_select_out(sw_254_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_254_module_data_in[7] ,
    \sw_254_module_data_in[6] ,
    \sw_254_module_data_in[5] ,
    \sw_254_module_data_in[4] ,
    \sw_254_module_data_in[3] ,
    \sw_254_module_data_in[2] ,
    \sw_254_module_data_in[1] ,
    \sw_254_module_data_in[0] }),
    .module_data_out({\sw_254_module_data_out[7] ,
    \sw_254_module_data_out[6] ,
    \sw_254_module_data_out[5] ,
    \sw_254_module_data_out[4] ,
    \sw_254_module_data_out[3] ,
    \sw_254_module_data_out[2] ,
    \sw_254_module_data_out[1] ,
    \sw_254_module_data_out[0] }));
 scanchain scanchain_255 (.clk_in(sw_254_clk_out),
    .clk_out(sw_255_clk_out),
    .data_in(sw_254_data_out),
    .data_out(sw_255_data_out),
    .latch_enable_in(sw_254_latch_out),
    .latch_enable_out(sw_255_latch_out),
    .scan_select_in(sw_254_scan_out),
    .scan_select_out(sw_255_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_255_module_data_in[7] ,
    \sw_255_module_data_in[6] ,
    \sw_255_module_data_in[5] ,
    \sw_255_module_data_in[4] ,
    \sw_255_module_data_in[3] ,
    \sw_255_module_data_in[2] ,
    \sw_255_module_data_in[1] ,
    \sw_255_module_data_in[0] }),
    .module_data_out({\sw_255_module_data_out[7] ,
    \sw_255_module_data_out[6] ,
    \sw_255_module_data_out[5] ,
    \sw_255_module_data_out[4] ,
    \sw_255_module_data_out[3] ,
    \sw_255_module_data_out[2] ,
    \sw_255_module_data_out[1] ,
    \sw_255_module_data_out[0] }));
 scanchain scanchain_256 (.clk_in(sw_255_clk_out),
    .clk_out(sw_256_clk_out),
    .data_in(sw_255_data_out),
    .data_out(sw_256_data_out),
    .latch_enable_in(sw_255_latch_out),
    .latch_enable_out(sw_256_latch_out),
    .scan_select_in(sw_255_scan_out),
    .scan_select_out(sw_256_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_256_module_data_in[7] ,
    \sw_256_module_data_in[6] ,
    \sw_256_module_data_in[5] ,
    \sw_256_module_data_in[4] ,
    \sw_256_module_data_in[3] ,
    \sw_256_module_data_in[2] ,
    \sw_256_module_data_in[1] ,
    \sw_256_module_data_in[0] }),
    .module_data_out({\sw_256_module_data_out[7] ,
    \sw_256_module_data_out[6] ,
    \sw_256_module_data_out[5] ,
    \sw_256_module_data_out[4] ,
    \sw_256_module_data_out[3] ,
    \sw_256_module_data_out[2] ,
    \sw_256_module_data_out[1] ,
    \sw_256_module_data_out[0] }));
 scanchain scanchain_257 (.clk_in(sw_256_clk_out),
    .clk_out(sw_257_clk_out),
    .data_in(sw_256_data_out),
    .data_out(sw_257_data_out),
    .latch_enable_in(sw_256_latch_out),
    .latch_enable_out(sw_257_latch_out),
    .scan_select_in(sw_256_scan_out),
    .scan_select_out(sw_257_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_257_module_data_in[7] ,
    \sw_257_module_data_in[6] ,
    \sw_257_module_data_in[5] ,
    \sw_257_module_data_in[4] ,
    \sw_257_module_data_in[3] ,
    \sw_257_module_data_in[2] ,
    \sw_257_module_data_in[1] ,
    \sw_257_module_data_in[0] }),
    .module_data_out({\sw_257_module_data_out[7] ,
    \sw_257_module_data_out[6] ,
    \sw_257_module_data_out[5] ,
    \sw_257_module_data_out[4] ,
    \sw_257_module_data_out[3] ,
    \sw_257_module_data_out[2] ,
    \sw_257_module_data_out[1] ,
    \sw_257_module_data_out[0] }));
 scanchain scanchain_258 (.clk_in(sw_257_clk_out),
    .clk_out(sw_258_clk_out),
    .data_in(sw_257_data_out),
    .data_out(sw_258_data_out),
    .latch_enable_in(sw_257_latch_out),
    .latch_enable_out(sw_258_latch_out),
    .scan_select_in(sw_257_scan_out),
    .scan_select_out(sw_258_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_258_module_data_in[7] ,
    \sw_258_module_data_in[6] ,
    \sw_258_module_data_in[5] ,
    \sw_258_module_data_in[4] ,
    \sw_258_module_data_in[3] ,
    \sw_258_module_data_in[2] ,
    \sw_258_module_data_in[1] ,
    \sw_258_module_data_in[0] }),
    .module_data_out({\sw_258_module_data_out[7] ,
    \sw_258_module_data_out[6] ,
    \sw_258_module_data_out[5] ,
    \sw_258_module_data_out[4] ,
    \sw_258_module_data_out[3] ,
    \sw_258_module_data_out[2] ,
    \sw_258_module_data_out[1] ,
    \sw_258_module_data_out[0] }));
 scanchain scanchain_259 (.clk_in(sw_258_clk_out),
    .clk_out(sw_259_clk_out),
    .data_in(sw_258_data_out),
    .data_out(sw_259_data_out),
    .latch_enable_in(sw_258_latch_out),
    .latch_enable_out(sw_259_latch_out),
    .scan_select_in(sw_258_scan_out),
    .scan_select_out(sw_259_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_259_module_data_in[7] ,
    \sw_259_module_data_in[6] ,
    \sw_259_module_data_in[5] ,
    \sw_259_module_data_in[4] ,
    \sw_259_module_data_in[3] ,
    \sw_259_module_data_in[2] ,
    \sw_259_module_data_in[1] ,
    \sw_259_module_data_in[0] }),
    .module_data_out({\sw_259_module_data_out[7] ,
    \sw_259_module_data_out[6] ,
    \sw_259_module_data_out[5] ,
    \sw_259_module_data_out[4] ,
    \sw_259_module_data_out[3] ,
    \sw_259_module_data_out[2] ,
    \sw_259_module_data_out[1] ,
    \sw_259_module_data_out[0] }));
 scanchain scanchain_26 (.clk_in(sw_025_clk_out),
    .clk_out(sw_026_clk_out),
    .data_in(sw_025_data_out),
    .data_out(sw_026_data_out),
    .latch_enable_in(sw_025_latch_out),
    .latch_enable_out(sw_026_latch_out),
    .scan_select_in(sw_025_scan_out),
    .scan_select_out(sw_026_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_026_module_data_in[7] ,
    \sw_026_module_data_in[6] ,
    \sw_026_module_data_in[5] ,
    \sw_026_module_data_in[4] ,
    \sw_026_module_data_in[3] ,
    \sw_026_module_data_in[2] ,
    \sw_026_module_data_in[1] ,
    \sw_026_module_data_in[0] }),
    .module_data_out({\sw_026_module_data_out[7] ,
    \sw_026_module_data_out[6] ,
    \sw_026_module_data_out[5] ,
    \sw_026_module_data_out[4] ,
    \sw_026_module_data_out[3] ,
    \sw_026_module_data_out[2] ,
    \sw_026_module_data_out[1] ,
    \sw_026_module_data_out[0] }));
 scanchain scanchain_260 (.clk_in(sw_259_clk_out),
    .clk_out(sw_260_clk_out),
    .data_in(sw_259_data_out),
    .data_out(sw_260_data_out),
    .latch_enable_in(sw_259_latch_out),
    .latch_enable_out(sw_260_latch_out),
    .scan_select_in(sw_259_scan_out),
    .scan_select_out(sw_260_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_260_module_data_in[7] ,
    \sw_260_module_data_in[6] ,
    \sw_260_module_data_in[5] ,
    \sw_260_module_data_in[4] ,
    \sw_260_module_data_in[3] ,
    \sw_260_module_data_in[2] ,
    \sw_260_module_data_in[1] ,
    \sw_260_module_data_in[0] }),
    .module_data_out({\sw_260_module_data_out[7] ,
    \sw_260_module_data_out[6] ,
    \sw_260_module_data_out[5] ,
    \sw_260_module_data_out[4] ,
    \sw_260_module_data_out[3] ,
    \sw_260_module_data_out[2] ,
    \sw_260_module_data_out[1] ,
    \sw_260_module_data_out[0] }));
 scanchain scanchain_261 (.clk_in(sw_260_clk_out),
    .clk_out(sw_261_clk_out),
    .data_in(sw_260_data_out),
    .data_out(sw_261_data_out),
    .latch_enable_in(sw_260_latch_out),
    .latch_enable_out(sw_261_latch_out),
    .scan_select_in(sw_260_scan_out),
    .scan_select_out(sw_261_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_261_module_data_in[7] ,
    \sw_261_module_data_in[6] ,
    \sw_261_module_data_in[5] ,
    \sw_261_module_data_in[4] ,
    \sw_261_module_data_in[3] ,
    \sw_261_module_data_in[2] ,
    \sw_261_module_data_in[1] ,
    \sw_261_module_data_in[0] }),
    .module_data_out({\sw_261_module_data_out[7] ,
    \sw_261_module_data_out[6] ,
    \sw_261_module_data_out[5] ,
    \sw_261_module_data_out[4] ,
    \sw_261_module_data_out[3] ,
    \sw_261_module_data_out[2] ,
    \sw_261_module_data_out[1] ,
    \sw_261_module_data_out[0] }));
 scanchain scanchain_262 (.clk_in(sw_261_clk_out),
    .clk_out(sw_262_clk_out),
    .data_in(sw_261_data_out),
    .data_out(sw_262_data_out),
    .latch_enable_in(sw_261_latch_out),
    .latch_enable_out(sw_262_latch_out),
    .scan_select_in(sw_261_scan_out),
    .scan_select_out(sw_262_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_262_module_data_in[7] ,
    \sw_262_module_data_in[6] ,
    \sw_262_module_data_in[5] ,
    \sw_262_module_data_in[4] ,
    \sw_262_module_data_in[3] ,
    \sw_262_module_data_in[2] ,
    \sw_262_module_data_in[1] ,
    \sw_262_module_data_in[0] }),
    .module_data_out({\sw_262_module_data_out[7] ,
    \sw_262_module_data_out[6] ,
    \sw_262_module_data_out[5] ,
    \sw_262_module_data_out[4] ,
    \sw_262_module_data_out[3] ,
    \sw_262_module_data_out[2] ,
    \sw_262_module_data_out[1] ,
    \sw_262_module_data_out[0] }));
 scanchain scanchain_263 (.clk_in(sw_262_clk_out),
    .clk_out(sw_263_clk_out),
    .data_in(sw_262_data_out),
    .data_out(sw_263_data_out),
    .latch_enable_in(sw_262_latch_out),
    .latch_enable_out(sw_263_latch_out),
    .scan_select_in(sw_262_scan_out),
    .scan_select_out(sw_263_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_263_module_data_in[7] ,
    \sw_263_module_data_in[6] ,
    \sw_263_module_data_in[5] ,
    \sw_263_module_data_in[4] ,
    \sw_263_module_data_in[3] ,
    \sw_263_module_data_in[2] ,
    \sw_263_module_data_in[1] ,
    \sw_263_module_data_in[0] }),
    .module_data_out({\sw_263_module_data_out[7] ,
    \sw_263_module_data_out[6] ,
    \sw_263_module_data_out[5] ,
    \sw_263_module_data_out[4] ,
    \sw_263_module_data_out[3] ,
    \sw_263_module_data_out[2] ,
    \sw_263_module_data_out[1] ,
    \sw_263_module_data_out[0] }));
 scanchain scanchain_264 (.clk_in(sw_263_clk_out),
    .clk_out(sw_264_clk_out),
    .data_in(sw_263_data_out),
    .data_out(sw_264_data_out),
    .latch_enable_in(sw_263_latch_out),
    .latch_enable_out(sw_264_latch_out),
    .scan_select_in(sw_263_scan_out),
    .scan_select_out(sw_264_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_264_module_data_in[7] ,
    \sw_264_module_data_in[6] ,
    \sw_264_module_data_in[5] ,
    \sw_264_module_data_in[4] ,
    \sw_264_module_data_in[3] ,
    \sw_264_module_data_in[2] ,
    \sw_264_module_data_in[1] ,
    \sw_264_module_data_in[0] }),
    .module_data_out({\sw_264_module_data_out[7] ,
    \sw_264_module_data_out[6] ,
    \sw_264_module_data_out[5] ,
    \sw_264_module_data_out[4] ,
    \sw_264_module_data_out[3] ,
    \sw_264_module_data_out[2] ,
    \sw_264_module_data_out[1] ,
    \sw_264_module_data_out[0] }));
 scanchain scanchain_265 (.clk_in(sw_264_clk_out),
    .clk_out(sw_265_clk_out),
    .data_in(sw_264_data_out),
    .data_out(sw_265_data_out),
    .latch_enable_in(sw_264_latch_out),
    .latch_enable_out(sw_265_latch_out),
    .scan_select_in(sw_264_scan_out),
    .scan_select_out(sw_265_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_265_module_data_in[7] ,
    \sw_265_module_data_in[6] ,
    \sw_265_module_data_in[5] ,
    \sw_265_module_data_in[4] ,
    \sw_265_module_data_in[3] ,
    \sw_265_module_data_in[2] ,
    \sw_265_module_data_in[1] ,
    \sw_265_module_data_in[0] }),
    .module_data_out({\sw_265_module_data_out[7] ,
    \sw_265_module_data_out[6] ,
    \sw_265_module_data_out[5] ,
    \sw_265_module_data_out[4] ,
    \sw_265_module_data_out[3] ,
    \sw_265_module_data_out[2] ,
    \sw_265_module_data_out[1] ,
    \sw_265_module_data_out[0] }));
 scanchain scanchain_266 (.clk_in(sw_265_clk_out),
    .clk_out(sw_266_clk_out),
    .data_in(sw_265_data_out),
    .data_out(sw_266_data_out),
    .latch_enable_in(sw_265_latch_out),
    .latch_enable_out(sw_266_latch_out),
    .scan_select_in(sw_265_scan_out),
    .scan_select_out(sw_266_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_266_module_data_in[7] ,
    \sw_266_module_data_in[6] ,
    \sw_266_module_data_in[5] ,
    \sw_266_module_data_in[4] ,
    \sw_266_module_data_in[3] ,
    \sw_266_module_data_in[2] ,
    \sw_266_module_data_in[1] ,
    \sw_266_module_data_in[0] }),
    .module_data_out({\sw_266_module_data_out[7] ,
    \sw_266_module_data_out[6] ,
    \sw_266_module_data_out[5] ,
    \sw_266_module_data_out[4] ,
    \sw_266_module_data_out[3] ,
    \sw_266_module_data_out[2] ,
    \sw_266_module_data_out[1] ,
    \sw_266_module_data_out[0] }));
 scanchain scanchain_267 (.clk_in(sw_266_clk_out),
    .clk_out(sw_267_clk_out),
    .data_in(sw_266_data_out),
    .data_out(sw_267_data_out),
    .latch_enable_in(sw_266_latch_out),
    .latch_enable_out(sw_267_latch_out),
    .scan_select_in(sw_266_scan_out),
    .scan_select_out(sw_267_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_267_module_data_in[7] ,
    \sw_267_module_data_in[6] ,
    \sw_267_module_data_in[5] ,
    \sw_267_module_data_in[4] ,
    \sw_267_module_data_in[3] ,
    \sw_267_module_data_in[2] ,
    \sw_267_module_data_in[1] ,
    \sw_267_module_data_in[0] }),
    .module_data_out({\sw_267_module_data_out[7] ,
    \sw_267_module_data_out[6] ,
    \sw_267_module_data_out[5] ,
    \sw_267_module_data_out[4] ,
    \sw_267_module_data_out[3] ,
    \sw_267_module_data_out[2] ,
    \sw_267_module_data_out[1] ,
    \sw_267_module_data_out[0] }));
 scanchain scanchain_268 (.clk_in(sw_267_clk_out),
    .clk_out(sw_268_clk_out),
    .data_in(sw_267_data_out),
    .data_out(sw_268_data_out),
    .latch_enable_in(sw_267_latch_out),
    .latch_enable_out(sw_268_latch_out),
    .scan_select_in(sw_267_scan_out),
    .scan_select_out(sw_268_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_268_module_data_in[7] ,
    \sw_268_module_data_in[6] ,
    \sw_268_module_data_in[5] ,
    \sw_268_module_data_in[4] ,
    \sw_268_module_data_in[3] ,
    \sw_268_module_data_in[2] ,
    \sw_268_module_data_in[1] ,
    \sw_268_module_data_in[0] }),
    .module_data_out({\sw_268_module_data_out[7] ,
    \sw_268_module_data_out[6] ,
    \sw_268_module_data_out[5] ,
    \sw_268_module_data_out[4] ,
    \sw_268_module_data_out[3] ,
    \sw_268_module_data_out[2] ,
    \sw_268_module_data_out[1] ,
    \sw_268_module_data_out[0] }));
 scanchain scanchain_269 (.clk_in(sw_268_clk_out),
    .clk_out(sw_269_clk_out),
    .data_in(sw_268_data_out),
    .data_out(sw_269_data_out),
    .latch_enable_in(sw_268_latch_out),
    .latch_enable_out(sw_269_latch_out),
    .scan_select_in(sw_268_scan_out),
    .scan_select_out(sw_269_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_269_module_data_in[7] ,
    \sw_269_module_data_in[6] ,
    \sw_269_module_data_in[5] ,
    \sw_269_module_data_in[4] ,
    \sw_269_module_data_in[3] ,
    \sw_269_module_data_in[2] ,
    \sw_269_module_data_in[1] ,
    \sw_269_module_data_in[0] }),
    .module_data_out({\sw_269_module_data_out[7] ,
    \sw_269_module_data_out[6] ,
    \sw_269_module_data_out[5] ,
    \sw_269_module_data_out[4] ,
    \sw_269_module_data_out[3] ,
    \sw_269_module_data_out[2] ,
    \sw_269_module_data_out[1] ,
    \sw_269_module_data_out[0] }));
 scanchain scanchain_27 (.clk_in(sw_026_clk_out),
    .clk_out(sw_027_clk_out),
    .data_in(sw_026_data_out),
    .data_out(sw_027_data_out),
    .latch_enable_in(sw_026_latch_out),
    .latch_enable_out(sw_027_latch_out),
    .scan_select_in(sw_026_scan_out),
    .scan_select_out(sw_027_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_027_module_data_in[7] ,
    \sw_027_module_data_in[6] ,
    \sw_027_module_data_in[5] ,
    \sw_027_module_data_in[4] ,
    \sw_027_module_data_in[3] ,
    \sw_027_module_data_in[2] ,
    \sw_027_module_data_in[1] ,
    \sw_027_module_data_in[0] }),
    .module_data_out({\sw_027_module_data_out[7] ,
    \sw_027_module_data_out[6] ,
    \sw_027_module_data_out[5] ,
    \sw_027_module_data_out[4] ,
    \sw_027_module_data_out[3] ,
    \sw_027_module_data_out[2] ,
    \sw_027_module_data_out[1] ,
    \sw_027_module_data_out[0] }));
 scanchain scanchain_270 (.clk_in(sw_269_clk_out),
    .clk_out(sw_270_clk_out),
    .data_in(sw_269_data_out),
    .data_out(sw_270_data_out),
    .latch_enable_in(sw_269_latch_out),
    .latch_enable_out(sw_270_latch_out),
    .scan_select_in(sw_269_scan_out),
    .scan_select_out(sw_270_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_270_module_data_in[7] ,
    \sw_270_module_data_in[6] ,
    \sw_270_module_data_in[5] ,
    \sw_270_module_data_in[4] ,
    \sw_270_module_data_in[3] ,
    \sw_270_module_data_in[2] ,
    \sw_270_module_data_in[1] ,
    \sw_270_module_data_in[0] }),
    .module_data_out({\sw_270_module_data_out[7] ,
    \sw_270_module_data_out[6] ,
    \sw_270_module_data_out[5] ,
    \sw_270_module_data_out[4] ,
    \sw_270_module_data_out[3] ,
    \sw_270_module_data_out[2] ,
    \sw_270_module_data_out[1] ,
    \sw_270_module_data_out[0] }));
 scanchain scanchain_271 (.clk_in(sw_270_clk_out),
    .clk_out(sw_271_clk_out),
    .data_in(sw_270_data_out),
    .data_out(sw_271_data_out),
    .latch_enable_in(sw_270_latch_out),
    .latch_enable_out(sw_271_latch_out),
    .scan_select_in(sw_270_scan_out),
    .scan_select_out(sw_271_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_271_module_data_in[7] ,
    \sw_271_module_data_in[6] ,
    \sw_271_module_data_in[5] ,
    \sw_271_module_data_in[4] ,
    \sw_271_module_data_in[3] ,
    \sw_271_module_data_in[2] ,
    \sw_271_module_data_in[1] ,
    \sw_271_module_data_in[0] }),
    .module_data_out({\sw_271_module_data_out[7] ,
    \sw_271_module_data_out[6] ,
    \sw_271_module_data_out[5] ,
    \sw_271_module_data_out[4] ,
    \sw_271_module_data_out[3] ,
    \sw_271_module_data_out[2] ,
    \sw_271_module_data_out[1] ,
    \sw_271_module_data_out[0] }));
 scanchain scanchain_272 (.clk_in(sw_271_clk_out),
    .clk_out(sw_272_clk_out),
    .data_in(sw_271_data_out),
    .data_out(sw_272_data_out),
    .latch_enable_in(sw_271_latch_out),
    .latch_enable_out(sw_272_latch_out),
    .scan_select_in(sw_271_scan_out),
    .scan_select_out(sw_272_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_272_module_data_in[7] ,
    \sw_272_module_data_in[6] ,
    \sw_272_module_data_in[5] ,
    \sw_272_module_data_in[4] ,
    \sw_272_module_data_in[3] ,
    \sw_272_module_data_in[2] ,
    \sw_272_module_data_in[1] ,
    \sw_272_module_data_in[0] }),
    .module_data_out({\sw_272_module_data_out[7] ,
    \sw_272_module_data_out[6] ,
    \sw_272_module_data_out[5] ,
    \sw_272_module_data_out[4] ,
    \sw_272_module_data_out[3] ,
    \sw_272_module_data_out[2] ,
    \sw_272_module_data_out[1] ,
    \sw_272_module_data_out[0] }));
 scanchain scanchain_273 (.clk_in(sw_272_clk_out),
    .clk_out(sw_273_clk_out),
    .data_in(sw_272_data_out),
    .data_out(sw_273_data_out),
    .latch_enable_in(sw_272_latch_out),
    .latch_enable_out(sw_273_latch_out),
    .scan_select_in(sw_272_scan_out),
    .scan_select_out(sw_273_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_273_module_data_in[7] ,
    \sw_273_module_data_in[6] ,
    \sw_273_module_data_in[5] ,
    \sw_273_module_data_in[4] ,
    \sw_273_module_data_in[3] ,
    \sw_273_module_data_in[2] ,
    \sw_273_module_data_in[1] ,
    \sw_273_module_data_in[0] }),
    .module_data_out({\sw_273_module_data_out[7] ,
    \sw_273_module_data_out[6] ,
    \sw_273_module_data_out[5] ,
    \sw_273_module_data_out[4] ,
    \sw_273_module_data_out[3] ,
    \sw_273_module_data_out[2] ,
    \sw_273_module_data_out[1] ,
    \sw_273_module_data_out[0] }));
 scanchain scanchain_274 (.clk_in(sw_273_clk_out),
    .clk_out(sw_274_clk_out),
    .data_in(sw_273_data_out),
    .data_out(sw_274_data_out),
    .latch_enable_in(sw_273_latch_out),
    .latch_enable_out(sw_274_latch_out),
    .scan_select_in(sw_273_scan_out),
    .scan_select_out(sw_274_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_274_module_data_in[7] ,
    \sw_274_module_data_in[6] ,
    \sw_274_module_data_in[5] ,
    \sw_274_module_data_in[4] ,
    \sw_274_module_data_in[3] ,
    \sw_274_module_data_in[2] ,
    \sw_274_module_data_in[1] ,
    \sw_274_module_data_in[0] }),
    .module_data_out({\sw_274_module_data_out[7] ,
    \sw_274_module_data_out[6] ,
    \sw_274_module_data_out[5] ,
    \sw_274_module_data_out[4] ,
    \sw_274_module_data_out[3] ,
    \sw_274_module_data_out[2] ,
    \sw_274_module_data_out[1] ,
    \sw_274_module_data_out[0] }));
 scanchain scanchain_275 (.clk_in(sw_274_clk_out),
    .clk_out(sw_275_clk_out),
    .data_in(sw_274_data_out),
    .data_out(sw_275_data_out),
    .latch_enable_in(sw_274_latch_out),
    .latch_enable_out(sw_275_latch_out),
    .scan_select_in(sw_274_scan_out),
    .scan_select_out(sw_275_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_275_module_data_in[7] ,
    \sw_275_module_data_in[6] ,
    \sw_275_module_data_in[5] ,
    \sw_275_module_data_in[4] ,
    \sw_275_module_data_in[3] ,
    \sw_275_module_data_in[2] ,
    \sw_275_module_data_in[1] ,
    \sw_275_module_data_in[0] }),
    .module_data_out({\sw_275_module_data_out[7] ,
    \sw_275_module_data_out[6] ,
    \sw_275_module_data_out[5] ,
    \sw_275_module_data_out[4] ,
    \sw_275_module_data_out[3] ,
    \sw_275_module_data_out[2] ,
    \sw_275_module_data_out[1] ,
    \sw_275_module_data_out[0] }));
 scanchain scanchain_276 (.clk_in(sw_275_clk_out),
    .clk_out(sw_276_clk_out),
    .data_in(sw_275_data_out),
    .data_out(sw_276_data_out),
    .latch_enable_in(sw_275_latch_out),
    .latch_enable_out(sw_276_latch_out),
    .scan_select_in(sw_275_scan_out),
    .scan_select_out(sw_276_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_276_module_data_in[7] ,
    \sw_276_module_data_in[6] ,
    \sw_276_module_data_in[5] ,
    \sw_276_module_data_in[4] ,
    \sw_276_module_data_in[3] ,
    \sw_276_module_data_in[2] ,
    \sw_276_module_data_in[1] ,
    \sw_276_module_data_in[0] }),
    .module_data_out({\sw_276_module_data_out[7] ,
    \sw_276_module_data_out[6] ,
    \sw_276_module_data_out[5] ,
    \sw_276_module_data_out[4] ,
    \sw_276_module_data_out[3] ,
    \sw_276_module_data_out[2] ,
    \sw_276_module_data_out[1] ,
    \sw_276_module_data_out[0] }));
 scanchain scanchain_277 (.clk_in(sw_276_clk_out),
    .clk_out(sw_277_clk_out),
    .data_in(sw_276_data_out),
    .data_out(sw_277_data_out),
    .latch_enable_in(sw_276_latch_out),
    .latch_enable_out(sw_277_latch_out),
    .scan_select_in(sw_276_scan_out),
    .scan_select_out(sw_277_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_277_module_data_in[7] ,
    \sw_277_module_data_in[6] ,
    \sw_277_module_data_in[5] ,
    \sw_277_module_data_in[4] ,
    \sw_277_module_data_in[3] ,
    \sw_277_module_data_in[2] ,
    \sw_277_module_data_in[1] ,
    \sw_277_module_data_in[0] }),
    .module_data_out({\sw_277_module_data_out[7] ,
    \sw_277_module_data_out[6] ,
    \sw_277_module_data_out[5] ,
    \sw_277_module_data_out[4] ,
    \sw_277_module_data_out[3] ,
    \sw_277_module_data_out[2] ,
    \sw_277_module_data_out[1] ,
    \sw_277_module_data_out[0] }));
 scanchain scanchain_278 (.clk_in(sw_277_clk_out),
    .clk_out(sw_278_clk_out),
    .data_in(sw_277_data_out),
    .data_out(sw_278_data_out),
    .latch_enable_in(sw_277_latch_out),
    .latch_enable_out(sw_278_latch_out),
    .scan_select_in(sw_277_scan_out),
    .scan_select_out(sw_278_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_278_module_data_in[7] ,
    \sw_278_module_data_in[6] ,
    \sw_278_module_data_in[5] ,
    \sw_278_module_data_in[4] ,
    \sw_278_module_data_in[3] ,
    \sw_278_module_data_in[2] ,
    \sw_278_module_data_in[1] ,
    \sw_278_module_data_in[0] }),
    .module_data_out({\sw_278_module_data_out[7] ,
    \sw_278_module_data_out[6] ,
    \sw_278_module_data_out[5] ,
    \sw_278_module_data_out[4] ,
    \sw_278_module_data_out[3] ,
    \sw_278_module_data_out[2] ,
    \sw_278_module_data_out[1] ,
    \sw_278_module_data_out[0] }));
 scanchain scanchain_279 (.clk_in(sw_278_clk_out),
    .clk_out(sw_279_clk_out),
    .data_in(sw_278_data_out),
    .data_out(sw_279_data_out),
    .latch_enable_in(sw_278_latch_out),
    .latch_enable_out(sw_279_latch_out),
    .scan_select_in(sw_278_scan_out),
    .scan_select_out(sw_279_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_279_module_data_in[7] ,
    \sw_279_module_data_in[6] ,
    \sw_279_module_data_in[5] ,
    \sw_279_module_data_in[4] ,
    \sw_279_module_data_in[3] ,
    \sw_279_module_data_in[2] ,
    \sw_279_module_data_in[1] ,
    \sw_279_module_data_in[0] }),
    .module_data_out({\sw_279_module_data_out[7] ,
    \sw_279_module_data_out[6] ,
    \sw_279_module_data_out[5] ,
    \sw_279_module_data_out[4] ,
    \sw_279_module_data_out[3] ,
    \sw_279_module_data_out[2] ,
    \sw_279_module_data_out[1] ,
    \sw_279_module_data_out[0] }));
 scanchain scanchain_28 (.clk_in(sw_027_clk_out),
    .clk_out(sw_028_clk_out),
    .data_in(sw_027_data_out),
    .data_out(sw_028_data_out),
    .latch_enable_in(sw_027_latch_out),
    .latch_enable_out(sw_028_latch_out),
    .scan_select_in(sw_027_scan_out),
    .scan_select_out(sw_028_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_028_module_data_in[7] ,
    \sw_028_module_data_in[6] ,
    \sw_028_module_data_in[5] ,
    \sw_028_module_data_in[4] ,
    \sw_028_module_data_in[3] ,
    \sw_028_module_data_in[2] ,
    \sw_028_module_data_in[1] ,
    \sw_028_module_data_in[0] }),
    .module_data_out({\sw_028_module_data_out[7] ,
    \sw_028_module_data_out[6] ,
    \sw_028_module_data_out[5] ,
    \sw_028_module_data_out[4] ,
    \sw_028_module_data_out[3] ,
    \sw_028_module_data_out[2] ,
    \sw_028_module_data_out[1] ,
    \sw_028_module_data_out[0] }));
 scanchain scanchain_280 (.clk_in(sw_279_clk_out),
    .clk_out(sw_280_clk_out),
    .data_in(sw_279_data_out),
    .data_out(sw_280_data_out),
    .latch_enable_in(sw_279_latch_out),
    .latch_enable_out(sw_280_latch_out),
    .scan_select_in(sw_279_scan_out),
    .scan_select_out(sw_280_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_280_module_data_in[7] ,
    \sw_280_module_data_in[6] ,
    \sw_280_module_data_in[5] ,
    \sw_280_module_data_in[4] ,
    \sw_280_module_data_in[3] ,
    \sw_280_module_data_in[2] ,
    \sw_280_module_data_in[1] ,
    \sw_280_module_data_in[0] }),
    .module_data_out({\sw_280_module_data_out[7] ,
    \sw_280_module_data_out[6] ,
    \sw_280_module_data_out[5] ,
    \sw_280_module_data_out[4] ,
    \sw_280_module_data_out[3] ,
    \sw_280_module_data_out[2] ,
    \sw_280_module_data_out[1] ,
    \sw_280_module_data_out[0] }));
 scanchain scanchain_281 (.clk_in(sw_280_clk_out),
    .clk_out(sw_281_clk_out),
    .data_in(sw_280_data_out),
    .data_out(sw_281_data_out),
    .latch_enable_in(sw_280_latch_out),
    .latch_enable_out(sw_281_latch_out),
    .scan_select_in(sw_280_scan_out),
    .scan_select_out(sw_281_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_281_module_data_in[7] ,
    \sw_281_module_data_in[6] ,
    \sw_281_module_data_in[5] ,
    \sw_281_module_data_in[4] ,
    \sw_281_module_data_in[3] ,
    \sw_281_module_data_in[2] ,
    \sw_281_module_data_in[1] ,
    \sw_281_module_data_in[0] }),
    .module_data_out({\sw_281_module_data_out[7] ,
    \sw_281_module_data_out[6] ,
    \sw_281_module_data_out[5] ,
    \sw_281_module_data_out[4] ,
    \sw_281_module_data_out[3] ,
    \sw_281_module_data_out[2] ,
    \sw_281_module_data_out[1] ,
    \sw_281_module_data_out[0] }));
 scanchain scanchain_282 (.clk_in(sw_281_clk_out),
    .clk_out(sw_282_clk_out),
    .data_in(sw_281_data_out),
    .data_out(sw_282_data_out),
    .latch_enable_in(sw_281_latch_out),
    .latch_enable_out(sw_282_latch_out),
    .scan_select_in(sw_281_scan_out),
    .scan_select_out(sw_282_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_282_module_data_in[7] ,
    \sw_282_module_data_in[6] ,
    \sw_282_module_data_in[5] ,
    \sw_282_module_data_in[4] ,
    \sw_282_module_data_in[3] ,
    \sw_282_module_data_in[2] ,
    \sw_282_module_data_in[1] ,
    \sw_282_module_data_in[0] }),
    .module_data_out({\sw_282_module_data_out[7] ,
    \sw_282_module_data_out[6] ,
    \sw_282_module_data_out[5] ,
    \sw_282_module_data_out[4] ,
    \sw_282_module_data_out[3] ,
    \sw_282_module_data_out[2] ,
    \sw_282_module_data_out[1] ,
    \sw_282_module_data_out[0] }));
 scanchain scanchain_283 (.clk_in(sw_282_clk_out),
    .clk_out(sw_283_clk_out),
    .data_in(sw_282_data_out),
    .data_out(sw_283_data_out),
    .latch_enable_in(sw_282_latch_out),
    .latch_enable_out(sw_283_latch_out),
    .scan_select_in(sw_282_scan_out),
    .scan_select_out(sw_283_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_283_module_data_in[7] ,
    \sw_283_module_data_in[6] ,
    \sw_283_module_data_in[5] ,
    \sw_283_module_data_in[4] ,
    \sw_283_module_data_in[3] ,
    \sw_283_module_data_in[2] ,
    \sw_283_module_data_in[1] ,
    \sw_283_module_data_in[0] }),
    .module_data_out({\sw_283_module_data_out[7] ,
    \sw_283_module_data_out[6] ,
    \sw_283_module_data_out[5] ,
    \sw_283_module_data_out[4] ,
    \sw_283_module_data_out[3] ,
    \sw_283_module_data_out[2] ,
    \sw_283_module_data_out[1] ,
    \sw_283_module_data_out[0] }));
 scanchain scanchain_284 (.clk_in(sw_283_clk_out),
    .clk_out(sw_284_clk_out),
    .data_in(sw_283_data_out),
    .data_out(sw_284_data_out),
    .latch_enable_in(sw_283_latch_out),
    .latch_enable_out(sw_284_latch_out),
    .scan_select_in(sw_283_scan_out),
    .scan_select_out(sw_284_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_284_module_data_in[7] ,
    \sw_284_module_data_in[6] ,
    \sw_284_module_data_in[5] ,
    \sw_284_module_data_in[4] ,
    \sw_284_module_data_in[3] ,
    \sw_284_module_data_in[2] ,
    \sw_284_module_data_in[1] ,
    \sw_284_module_data_in[0] }),
    .module_data_out({\sw_284_module_data_out[7] ,
    \sw_284_module_data_out[6] ,
    \sw_284_module_data_out[5] ,
    \sw_284_module_data_out[4] ,
    \sw_284_module_data_out[3] ,
    \sw_284_module_data_out[2] ,
    \sw_284_module_data_out[1] ,
    \sw_284_module_data_out[0] }));
 scanchain scanchain_285 (.clk_in(sw_284_clk_out),
    .clk_out(sw_285_clk_out),
    .data_in(sw_284_data_out),
    .data_out(sw_285_data_out),
    .latch_enable_in(sw_284_latch_out),
    .latch_enable_out(sw_285_latch_out),
    .scan_select_in(sw_284_scan_out),
    .scan_select_out(sw_285_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_285_module_data_in[7] ,
    \sw_285_module_data_in[6] ,
    \sw_285_module_data_in[5] ,
    \sw_285_module_data_in[4] ,
    \sw_285_module_data_in[3] ,
    \sw_285_module_data_in[2] ,
    \sw_285_module_data_in[1] ,
    \sw_285_module_data_in[0] }),
    .module_data_out({\sw_285_module_data_out[7] ,
    \sw_285_module_data_out[6] ,
    \sw_285_module_data_out[5] ,
    \sw_285_module_data_out[4] ,
    \sw_285_module_data_out[3] ,
    \sw_285_module_data_out[2] ,
    \sw_285_module_data_out[1] ,
    \sw_285_module_data_out[0] }));
 scanchain scanchain_286 (.clk_in(sw_285_clk_out),
    .clk_out(sw_286_clk_out),
    .data_in(sw_285_data_out),
    .data_out(sw_286_data_out),
    .latch_enable_in(sw_285_latch_out),
    .latch_enable_out(sw_286_latch_out),
    .scan_select_in(sw_285_scan_out),
    .scan_select_out(sw_286_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_286_module_data_in[7] ,
    \sw_286_module_data_in[6] ,
    \sw_286_module_data_in[5] ,
    \sw_286_module_data_in[4] ,
    \sw_286_module_data_in[3] ,
    \sw_286_module_data_in[2] ,
    \sw_286_module_data_in[1] ,
    \sw_286_module_data_in[0] }),
    .module_data_out({\sw_286_module_data_out[7] ,
    \sw_286_module_data_out[6] ,
    \sw_286_module_data_out[5] ,
    \sw_286_module_data_out[4] ,
    \sw_286_module_data_out[3] ,
    \sw_286_module_data_out[2] ,
    \sw_286_module_data_out[1] ,
    \sw_286_module_data_out[0] }));
 scanchain scanchain_287 (.clk_in(sw_286_clk_out),
    .clk_out(sw_287_clk_out),
    .data_in(sw_286_data_out),
    .data_out(sw_287_data_out),
    .latch_enable_in(sw_286_latch_out),
    .latch_enable_out(sw_287_latch_out),
    .scan_select_in(sw_286_scan_out),
    .scan_select_out(sw_287_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_287_module_data_in[7] ,
    \sw_287_module_data_in[6] ,
    \sw_287_module_data_in[5] ,
    \sw_287_module_data_in[4] ,
    \sw_287_module_data_in[3] ,
    \sw_287_module_data_in[2] ,
    \sw_287_module_data_in[1] ,
    \sw_287_module_data_in[0] }),
    .module_data_out({\sw_287_module_data_out[7] ,
    \sw_287_module_data_out[6] ,
    \sw_287_module_data_out[5] ,
    \sw_287_module_data_out[4] ,
    \sw_287_module_data_out[3] ,
    \sw_287_module_data_out[2] ,
    \sw_287_module_data_out[1] ,
    \sw_287_module_data_out[0] }));
 scanchain scanchain_288 (.clk_in(sw_287_clk_out),
    .clk_out(sw_288_clk_out),
    .data_in(sw_287_data_out),
    .data_out(sw_288_data_out),
    .latch_enable_in(sw_287_latch_out),
    .latch_enable_out(sw_288_latch_out),
    .scan_select_in(sw_287_scan_out),
    .scan_select_out(sw_288_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_288_module_data_in[7] ,
    \sw_288_module_data_in[6] ,
    \sw_288_module_data_in[5] ,
    \sw_288_module_data_in[4] ,
    \sw_288_module_data_in[3] ,
    \sw_288_module_data_in[2] ,
    \sw_288_module_data_in[1] ,
    \sw_288_module_data_in[0] }),
    .module_data_out({\sw_288_module_data_out[7] ,
    \sw_288_module_data_out[6] ,
    \sw_288_module_data_out[5] ,
    \sw_288_module_data_out[4] ,
    \sw_288_module_data_out[3] ,
    \sw_288_module_data_out[2] ,
    \sw_288_module_data_out[1] ,
    \sw_288_module_data_out[0] }));
 scanchain scanchain_289 (.clk_in(sw_288_clk_out),
    .clk_out(sw_289_clk_out),
    .data_in(sw_288_data_out),
    .data_out(sw_289_data_out),
    .latch_enable_in(sw_288_latch_out),
    .latch_enable_out(sw_289_latch_out),
    .scan_select_in(sw_288_scan_out),
    .scan_select_out(sw_289_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_289_module_data_in[7] ,
    \sw_289_module_data_in[6] ,
    \sw_289_module_data_in[5] ,
    \sw_289_module_data_in[4] ,
    \sw_289_module_data_in[3] ,
    \sw_289_module_data_in[2] ,
    \sw_289_module_data_in[1] ,
    \sw_289_module_data_in[0] }),
    .module_data_out({\sw_289_module_data_out[7] ,
    \sw_289_module_data_out[6] ,
    \sw_289_module_data_out[5] ,
    \sw_289_module_data_out[4] ,
    \sw_289_module_data_out[3] ,
    \sw_289_module_data_out[2] ,
    \sw_289_module_data_out[1] ,
    \sw_289_module_data_out[0] }));
 scanchain scanchain_29 (.clk_in(sw_028_clk_out),
    .clk_out(sw_029_clk_out),
    .data_in(sw_028_data_out),
    .data_out(sw_029_data_out),
    .latch_enable_in(sw_028_latch_out),
    .latch_enable_out(sw_029_latch_out),
    .scan_select_in(sw_028_scan_out),
    .scan_select_out(sw_029_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_029_module_data_in[7] ,
    \sw_029_module_data_in[6] ,
    \sw_029_module_data_in[5] ,
    \sw_029_module_data_in[4] ,
    \sw_029_module_data_in[3] ,
    \sw_029_module_data_in[2] ,
    \sw_029_module_data_in[1] ,
    \sw_029_module_data_in[0] }),
    .module_data_out({\sw_029_module_data_out[7] ,
    \sw_029_module_data_out[6] ,
    \sw_029_module_data_out[5] ,
    \sw_029_module_data_out[4] ,
    \sw_029_module_data_out[3] ,
    \sw_029_module_data_out[2] ,
    \sw_029_module_data_out[1] ,
    \sw_029_module_data_out[0] }));
 scanchain scanchain_290 (.clk_in(sw_289_clk_out),
    .clk_out(sw_290_clk_out),
    .data_in(sw_289_data_out),
    .data_out(sw_290_data_out),
    .latch_enable_in(sw_289_latch_out),
    .latch_enable_out(sw_290_latch_out),
    .scan_select_in(sw_289_scan_out),
    .scan_select_out(sw_290_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_290_module_data_in[7] ,
    \sw_290_module_data_in[6] ,
    \sw_290_module_data_in[5] ,
    \sw_290_module_data_in[4] ,
    \sw_290_module_data_in[3] ,
    \sw_290_module_data_in[2] ,
    \sw_290_module_data_in[1] ,
    \sw_290_module_data_in[0] }),
    .module_data_out({\sw_290_module_data_out[7] ,
    \sw_290_module_data_out[6] ,
    \sw_290_module_data_out[5] ,
    \sw_290_module_data_out[4] ,
    \sw_290_module_data_out[3] ,
    \sw_290_module_data_out[2] ,
    \sw_290_module_data_out[1] ,
    \sw_290_module_data_out[0] }));
 scanchain scanchain_291 (.clk_in(sw_290_clk_out),
    .clk_out(sw_291_clk_out),
    .data_in(sw_290_data_out),
    .data_out(sw_291_data_out),
    .latch_enable_in(sw_290_latch_out),
    .latch_enable_out(sw_291_latch_out),
    .scan_select_in(sw_290_scan_out),
    .scan_select_out(sw_291_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_291_module_data_in[7] ,
    \sw_291_module_data_in[6] ,
    \sw_291_module_data_in[5] ,
    \sw_291_module_data_in[4] ,
    \sw_291_module_data_in[3] ,
    \sw_291_module_data_in[2] ,
    \sw_291_module_data_in[1] ,
    \sw_291_module_data_in[0] }),
    .module_data_out({\sw_291_module_data_out[7] ,
    \sw_291_module_data_out[6] ,
    \sw_291_module_data_out[5] ,
    \sw_291_module_data_out[4] ,
    \sw_291_module_data_out[3] ,
    \sw_291_module_data_out[2] ,
    \sw_291_module_data_out[1] ,
    \sw_291_module_data_out[0] }));
 scanchain scanchain_292 (.clk_in(sw_291_clk_out),
    .clk_out(sw_292_clk_out),
    .data_in(sw_291_data_out),
    .data_out(sw_292_data_out),
    .latch_enable_in(sw_291_latch_out),
    .latch_enable_out(sw_292_latch_out),
    .scan_select_in(sw_291_scan_out),
    .scan_select_out(sw_292_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_292_module_data_in[7] ,
    \sw_292_module_data_in[6] ,
    \sw_292_module_data_in[5] ,
    \sw_292_module_data_in[4] ,
    \sw_292_module_data_in[3] ,
    \sw_292_module_data_in[2] ,
    \sw_292_module_data_in[1] ,
    \sw_292_module_data_in[0] }),
    .module_data_out({\sw_292_module_data_out[7] ,
    \sw_292_module_data_out[6] ,
    \sw_292_module_data_out[5] ,
    \sw_292_module_data_out[4] ,
    \sw_292_module_data_out[3] ,
    \sw_292_module_data_out[2] ,
    \sw_292_module_data_out[1] ,
    \sw_292_module_data_out[0] }));
 scanchain scanchain_293 (.clk_in(sw_292_clk_out),
    .clk_out(sw_293_clk_out),
    .data_in(sw_292_data_out),
    .data_out(sw_293_data_out),
    .latch_enable_in(sw_292_latch_out),
    .latch_enable_out(sw_293_latch_out),
    .scan_select_in(sw_292_scan_out),
    .scan_select_out(sw_293_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_293_module_data_in[7] ,
    \sw_293_module_data_in[6] ,
    \sw_293_module_data_in[5] ,
    \sw_293_module_data_in[4] ,
    \sw_293_module_data_in[3] ,
    \sw_293_module_data_in[2] ,
    \sw_293_module_data_in[1] ,
    \sw_293_module_data_in[0] }),
    .module_data_out({\sw_293_module_data_out[7] ,
    \sw_293_module_data_out[6] ,
    \sw_293_module_data_out[5] ,
    \sw_293_module_data_out[4] ,
    \sw_293_module_data_out[3] ,
    \sw_293_module_data_out[2] ,
    \sw_293_module_data_out[1] ,
    \sw_293_module_data_out[0] }));
 scanchain scanchain_294 (.clk_in(sw_293_clk_out),
    .clk_out(sw_294_clk_out),
    .data_in(sw_293_data_out),
    .data_out(sw_294_data_out),
    .latch_enable_in(sw_293_latch_out),
    .latch_enable_out(sw_294_latch_out),
    .scan_select_in(sw_293_scan_out),
    .scan_select_out(sw_294_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_294_module_data_in[7] ,
    \sw_294_module_data_in[6] ,
    \sw_294_module_data_in[5] ,
    \sw_294_module_data_in[4] ,
    \sw_294_module_data_in[3] ,
    \sw_294_module_data_in[2] ,
    \sw_294_module_data_in[1] ,
    \sw_294_module_data_in[0] }),
    .module_data_out({\sw_294_module_data_out[7] ,
    \sw_294_module_data_out[6] ,
    \sw_294_module_data_out[5] ,
    \sw_294_module_data_out[4] ,
    \sw_294_module_data_out[3] ,
    \sw_294_module_data_out[2] ,
    \sw_294_module_data_out[1] ,
    \sw_294_module_data_out[0] }));
 scanchain scanchain_295 (.clk_in(sw_294_clk_out),
    .clk_out(sw_295_clk_out),
    .data_in(sw_294_data_out),
    .data_out(sw_295_data_out),
    .latch_enable_in(sw_294_latch_out),
    .latch_enable_out(sw_295_latch_out),
    .scan_select_in(sw_294_scan_out),
    .scan_select_out(sw_295_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_295_module_data_in[7] ,
    \sw_295_module_data_in[6] ,
    \sw_295_module_data_in[5] ,
    \sw_295_module_data_in[4] ,
    \sw_295_module_data_in[3] ,
    \sw_295_module_data_in[2] ,
    \sw_295_module_data_in[1] ,
    \sw_295_module_data_in[0] }),
    .module_data_out({\sw_295_module_data_out[7] ,
    \sw_295_module_data_out[6] ,
    \sw_295_module_data_out[5] ,
    \sw_295_module_data_out[4] ,
    \sw_295_module_data_out[3] ,
    \sw_295_module_data_out[2] ,
    \sw_295_module_data_out[1] ,
    \sw_295_module_data_out[0] }));
 scanchain scanchain_296 (.clk_in(sw_295_clk_out),
    .clk_out(sw_296_clk_out),
    .data_in(sw_295_data_out),
    .data_out(sw_296_data_out),
    .latch_enable_in(sw_295_latch_out),
    .latch_enable_out(sw_296_latch_out),
    .scan_select_in(sw_295_scan_out),
    .scan_select_out(sw_296_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_296_module_data_in[7] ,
    \sw_296_module_data_in[6] ,
    \sw_296_module_data_in[5] ,
    \sw_296_module_data_in[4] ,
    \sw_296_module_data_in[3] ,
    \sw_296_module_data_in[2] ,
    \sw_296_module_data_in[1] ,
    \sw_296_module_data_in[0] }),
    .module_data_out({\sw_296_module_data_out[7] ,
    \sw_296_module_data_out[6] ,
    \sw_296_module_data_out[5] ,
    \sw_296_module_data_out[4] ,
    \sw_296_module_data_out[3] ,
    \sw_296_module_data_out[2] ,
    \sw_296_module_data_out[1] ,
    \sw_296_module_data_out[0] }));
 scanchain scanchain_297 (.clk_in(sw_296_clk_out),
    .clk_out(sw_297_clk_out),
    .data_in(sw_296_data_out),
    .data_out(sw_297_data_out),
    .latch_enable_in(sw_296_latch_out),
    .latch_enable_out(sw_297_latch_out),
    .scan_select_in(sw_296_scan_out),
    .scan_select_out(sw_297_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_297_module_data_in[7] ,
    \sw_297_module_data_in[6] ,
    \sw_297_module_data_in[5] ,
    \sw_297_module_data_in[4] ,
    \sw_297_module_data_in[3] ,
    \sw_297_module_data_in[2] ,
    \sw_297_module_data_in[1] ,
    \sw_297_module_data_in[0] }),
    .module_data_out({\sw_297_module_data_out[7] ,
    \sw_297_module_data_out[6] ,
    \sw_297_module_data_out[5] ,
    \sw_297_module_data_out[4] ,
    \sw_297_module_data_out[3] ,
    \sw_297_module_data_out[2] ,
    \sw_297_module_data_out[1] ,
    \sw_297_module_data_out[0] }));
 scanchain scanchain_298 (.clk_in(sw_297_clk_out),
    .clk_out(sw_298_clk_out),
    .data_in(sw_297_data_out),
    .data_out(sw_298_data_out),
    .latch_enable_in(sw_297_latch_out),
    .latch_enable_out(sw_298_latch_out),
    .scan_select_in(sw_297_scan_out),
    .scan_select_out(sw_298_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_298_module_data_in[7] ,
    \sw_298_module_data_in[6] ,
    \sw_298_module_data_in[5] ,
    \sw_298_module_data_in[4] ,
    \sw_298_module_data_in[3] ,
    \sw_298_module_data_in[2] ,
    \sw_298_module_data_in[1] ,
    \sw_298_module_data_in[0] }),
    .module_data_out({\sw_298_module_data_out[7] ,
    \sw_298_module_data_out[6] ,
    \sw_298_module_data_out[5] ,
    \sw_298_module_data_out[4] ,
    \sw_298_module_data_out[3] ,
    \sw_298_module_data_out[2] ,
    \sw_298_module_data_out[1] ,
    \sw_298_module_data_out[0] }));
 scanchain scanchain_299 (.clk_in(sw_298_clk_out),
    .clk_out(sw_299_clk_out),
    .data_in(sw_298_data_out),
    .data_out(sw_299_data_out),
    .latch_enable_in(sw_298_latch_out),
    .latch_enable_out(sw_299_latch_out),
    .scan_select_in(sw_298_scan_out),
    .scan_select_out(sw_299_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_299_module_data_in[7] ,
    \sw_299_module_data_in[6] ,
    \sw_299_module_data_in[5] ,
    \sw_299_module_data_in[4] ,
    \sw_299_module_data_in[3] ,
    \sw_299_module_data_in[2] ,
    \sw_299_module_data_in[1] ,
    \sw_299_module_data_in[0] }),
    .module_data_out({\sw_299_module_data_out[7] ,
    \sw_299_module_data_out[6] ,
    \sw_299_module_data_out[5] ,
    \sw_299_module_data_out[4] ,
    \sw_299_module_data_out[3] ,
    \sw_299_module_data_out[2] ,
    \sw_299_module_data_out[1] ,
    \sw_299_module_data_out[0] }));
 scanchain scanchain_3 (.clk_in(sw_002_clk_out),
    .clk_out(sw_003_clk_out),
    .data_in(sw_002_data_out),
    .data_out(sw_003_data_out),
    .latch_enable_in(sw_002_latch_out),
    .latch_enable_out(sw_003_latch_out),
    .scan_select_in(sw_002_scan_out),
    .scan_select_out(sw_003_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_003_module_data_in[7] ,
    \sw_003_module_data_in[6] ,
    \sw_003_module_data_in[5] ,
    \sw_003_module_data_in[4] ,
    \sw_003_module_data_in[3] ,
    \sw_003_module_data_in[2] ,
    \sw_003_module_data_in[1] ,
    \sw_003_module_data_in[0] }),
    .module_data_out({\sw_003_module_data_out[7] ,
    \sw_003_module_data_out[6] ,
    \sw_003_module_data_out[5] ,
    \sw_003_module_data_out[4] ,
    \sw_003_module_data_out[3] ,
    \sw_003_module_data_out[2] ,
    \sw_003_module_data_out[1] ,
    \sw_003_module_data_out[0] }));
 scanchain scanchain_30 (.clk_in(sw_029_clk_out),
    .clk_out(sw_030_clk_out),
    .data_in(sw_029_data_out),
    .data_out(sw_030_data_out),
    .latch_enable_in(sw_029_latch_out),
    .latch_enable_out(sw_030_latch_out),
    .scan_select_in(sw_029_scan_out),
    .scan_select_out(sw_030_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_030_module_data_in[7] ,
    \sw_030_module_data_in[6] ,
    \sw_030_module_data_in[5] ,
    \sw_030_module_data_in[4] ,
    \sw_030_module_data_in[3] ,
    \sw_030_module_data_in[2] ,
    \sw_030_module_data_in[1] ,
    \sw_030_module_data_in[0] }),
    .module_data_out({\sw_030_module_data_out[7] ,
    \sw_030_module_data_out[6] ,
    \sw_030_module_data_out[5] ,
    \sw_030_module_data_out[4] ,
    \sw_030_module_data_out[3] ,
    \sw_030_module_data_out[2] ,
    \sw_030_module_data_out[1] ,
    \sw_030_module_data_out[0] }));
 scanchain scanchain_300 (.clk_in(sw_299_clk_out),
    .clk_out(sw_300_clk_out),
    .data_in(sw_299_data_out),
    .data_out(sw_300_data_out),
    .latch_enable_in(sw_299_latch_out),
    .latch_enable_out(sw_300_latch_out),
    .scan_select_in(sw_299_scan_out),
    .scan_select_out(sw_300_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_300_module_data_in[7] ,
    \sw_300_module_data_in[6] ,
    \sw_300_module_data_in[5] ,
    \sw_300_module_data_in[4] ,
    \sw_300_module_data_in[3] ,
    \sw_300_module_data_in[2] ,
    \sw_300_module_data_in[1] ,
    \sw_300_module_data_in[0] }),
    .module_data_out({\sw_300_module_data_out[7] ,
    \sw_300_module_data_out[6] ,
    \sw_300_module_data_out[5] ,
    \sw_300_module_data_out[4] ,
    \sw_300_module_data_out[3] ,
    \sw_300_module_data_out[2] ,
    \sw_300_module_data_out[1] ,
    \sw_300_module_data_out[0] }));
 scanchain scanchain_301 (.clk_in(sw_300_clk_out),
    .clk_out(sw_301_clk_out),
    .data_in(sw_300_data_out),
    .data_out(sw_301_data_out),
    .latch_enable_in(sw_300_latch_out),
    .latch_enable_out(sw_301_latch_out),
    .scan_select_in(sw_300_scan_out),
    .scan_select_out(sw_301_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_301_module_data_in[7] ,
    \sw_301_module_data_in[6] ,
    \sw_301_module_data_in[5] ,
    \sw_301_module_data_in[4] ,
    \sw_301_module_data_in[3] ,
    \sw_301_module_data_in[2] ,
    \sw_301_module_data_in[1] ,
    \sw_301_module_data_in[0] }),
    .module_data_out({\sw_301_module_data_out[7] ,
    \sw_301_module_data_out[6] ,
    \sw_301_module_data_out[5] ,
    \sw_301_module_data_out[4] ,
    \sw_301_module_data_out[3] ,
    \sw_301_module_data_out[2] ,
    \sw_301_module_data_out[1] ,
    \sw_301_module_data_out[0] }));
 scanchain scanchain_302 (.clk_in(sw_301_clk_out),
    .clk_out(sw_302_clk_out),
    .data_in(sw_301_data_out),
    .data_out(sw_302_data_out),
    .latch_enable_in(sw_301_latch_out),
    .latch_enable_out(sw_302_latch_out),
    .scan_select_in(sw_301_scan_out),
    .scan_select_out(sw_302_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_302_module_data_in[7] ,
    \sw_302_module_data_in[6] ,
    \sw_302_module_data_in[5] ,
    \sw_302_module_data_in[4] ,
    \sw_302_module_data_in[3] ,
    \sw_302_module_data_in[2] ,
    \sw_302_module_data_in[1] ,
    \sw_302_module_data_in[0] }),
    .module_data_out({\sw_302_module_data_out[7] ,
    \sw_302_module_data_out[6] ,
    \sw_302_module_data_out[5] ,
    \sw_302_module_data_out[4] ,
    \sw_302_module_data_out[3] ,
    \sw_302_module_data_out[2] ,
    \sw_302_module_data_out[1] ,
    \sw_302_module_data_out[0] }));
 scanchain scanchain_303 (.clk_in(sw_302_clk_out),
    .clk_out(sw_303_clk_out),
    .data_in(sw_302_data_out),
    .data_out(sw_303_data_out),
    .latch_enable_in(sw_302_latch_out),
    .latch_enable_out(sw_303_latch_out),
    .scan_select_in(sw_302_scan_out),
    .scan_select_out(sw_303_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_303_module_data_in[7] ,
    \sw_303_module_data_in[6] ,
    \sw_303_module_data_in[5] ,
    \sw_303_module_data_in[4] ,
    \sw_303_module_data_in[3] ,
    \sw_303_module_data_in[2] ,
    \sw_303_module_data_in[1] ,
    \sw_303_module_data_in[0] }),
    .module_data_out({\sw_303_module_data_out[7] ,
    \sw_303_module_data_out[6] ,
    \sw_303_module_data_out[5] ,
    \sw_303_module_data_out[4] ,
    \sw_303_module_data_out[3] ,
    \sw_303_module_data_out[2] ,
    \sw_303_module_data_out[1] ,
    \sw_303_module_data_out[0] }));
 scanchain scanchain_304 (.clk_in(sw_303_clk_out),
    .clk_out(sw_304_clk_out),
    .data_in(sw_303_data_out),
    .data_out(sw_304_data_out),
    .latch_enable_in(sw_303_latch_out),
    .latch_enable_out(sw_304_latch_out),
    .scan_select_in(sw_303_scan_out),
    .scan_select_out(sw_304_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_304_module_data_in[7] ,
    \sw_304_module_data_in[6] ,
    \sw_304_module_data_in[5] ,
    \sw_304_module_data_in[4] ,
    \sw_304_module_data_in[3] ,
    \sw_304_module_data_in[2] ,
    \sw_304_module_data_in[1] ,
    \sw_304_module_data_in[0] }),
    .module_data_out({\sw_304_module_data_out[7] ,
    \sw_304_module_data_out[6] ,
    \sw_304_module_data_out[5] ,
    \sw_304_module_data_out[4] ,
    \sw_304_module_data_out[3] ,
    \sw_304_module_data_out[2] ,
    \sw_304_module_data_out[1] ,
    \sw_304_module_data_out[0] }));
 scanchain scanchain_305 (.clk_in(sw_304_clk_out),
    .clk_out(sw_305_clk_out),
    .data_in(sw_304_data_out),
    .data_out(sw_305_data_out),
    .latch_enable_in(sw_304_latch_out),
    .latch_enable_out(sw_305_latch_out),
    .scan_select_in(sw_304_scan_out),
    .scan_select_out(sw_305_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_305_module_data_in[7] ,
    \sw_305_module_data_in[6] ,
    \sw_305_module_data_in[5] ,
    \sw_305_module_data_in[4] ,
    \sw_305_module_data_in[3] ,
    \sw_305_module_data_in[2] ,
    \sw_305_module_data_in[1] ,
    \sw_305_module_data_in[0] }),
    .module_data_out({\sw_305_module_data_out[7] ,
    \sw_305_module_data_out[6] ,
    \sw_305_module_data_out[5] ,
    \sw_305_module_data_out[4] ,
    \sw_305_module_data_out[3] ,
    \sw_305_module_data_out[2] ,
    \sw_305_module_data_out[1] ,
    \sw_305_module_data_out[0] }));
 scanchain scanchain_306 (.clk_in(sw_305_clk_out),
    .clk_out(sw_306_clk_out),
    .data_in(sw_305_data_out),
    .data_out(sw_306_data_out),
    .latch_enable_in(sw_305_latch_out),
    .latch_enable_out(sw_306_latch_out),
    .scan_select_in(sw_305_scan_out),
    .scan_select_out(sw_306_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_306_module_data_in[7] ,
    \sw_306_module_data_in[6] ,
    \sw_306_module_data_in[5] ,
    \sw_306_module_data_in[4] ,
    \sw_306_module_data_in[3] ,
    \sw_306_module_data_in[2] ,
    \sw_306_module_data_in[1] ,
    \sw_306_module_data_in[0] }),
    .module_data_out({\sw_306_module_data_out[7] ,
    \sw_306_module_data_out[6] ,
    \sw_306_module_data_out[5] ,
    \sw_306_module_data_out[4] ,
    \sw_306_module_data_out[3] ,
    \sw_306_module_data_out[2] ,
    \sw_306_module_data_out[1] ,
    \sw_306_module_data_out[0] }));
 scanchain scanchain_307 (.clk_in(sw_306_clk_out),
    .clk_out(sw_307_clk_out),
    .data_in(sw_306_data_out),
    .data_out(sw_307_data_out),
    .latch_enable_in(sw_306_latch_out),
    .latch_enable_out(sw_307_latch_out),
    .scan_select_in(sw_306_scan_out),
    .scan_select_out(sw_307_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_307_module_data_in[7] ,
    \sw_307_module_data_in[6] ,
    \sw_307_module_data_in[5] ,
    \sw_307_module_data_in[4] ,
    \sw_307_module_data_in[3] ,
    \sw_307_module_data_in[2] ,
    \sw_307_module_data_in[1] ,
    \sw_307_module_data_in[0] }),
    .module_data_out({\sw_307_module_data_out[7] ,
    \sw_307_module_data_out[6] ,
    \sw_307_module_data_out[5] ,
    \sw_307_module_data_out[4] ,
    \sw_307_module_data_out[3] ,
    \sw_307_module_data_out[2] ,
    \sw_307_module_data_out[1] ,
    \sw_307_module_data_out[0] }));
 scanchain scanchain_308 (.clk_in(sw_307_clk_out),
    .clk_out(sw_308_clk_out),
    .data_in(sw_307_data_out),
    .data_out(sw_308_data_out),
    .latch_enable_in(sw_307_latch_out),
    .latch_enable_out(sw_308_latch_out),
    .scan_select_in(sw_307_scan_out),
    .scan_select_out(sw_308_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_308_module_data_in[7] ,
    \sw_308_module_data_in[6] ,
    \sw_308_module_data_in[5] ,
    \sw_308_module_data_in[4] ,
    \sw_308_module_data_in[3] ,
    \sw_308_module_data_in[2] ,
    \sw_308_module_data_in[1] ,
    \sw_308_module_data_in[0] }),
    .module_data_out({\sw_308_module_data_out[7] ,
    \sw_308_module_data_out[6] ,
    \sw_308_module_data_out[5] ,
    \sw_308_module_data_out[4] ,
    \sw_308_module_data_out[3] ,
    \sw_308_module_data_out[2] ,
    \sw_308_module_data_out[1] ,
    \sw_308_module_data_out[0] }));
 scanchain scanchain_309 (.clk_in(sw_308_clk_out),
    .clk_out(sw_309_clk_out),
    .data_in(sw_308_data_out),
    .data_out(sw_309_data_out),
    .latch_enable_in(sw_308_latch_out),
    .latch_enable_out(sw_309_latch_out),
    .scan_select_in(sw_308_scan_out),
    .scan_select_out(sw_309_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_309_module_data_in[7] ,
    \sw_309_module_data_in[6] ,
    \sw_309_module_data_in[5] ,
    \sw_309_module_data_in[4] ,
    \sw_309_module_data_in[3] ,
    \sw_309_module_data_in[2] ,
    \sw_309_module_data_in[1] ,
    \sw_309_module_data_in[0] }),
    .module_data_out({\sw_309_module_data_out[7] ,
    \sw_309_module_data_out[6] ,
    \sw_309_module_data_out[5] ,
    \sw_309_module_data_out[4] ,
    \sw_309_module_data_out[3] ,
    \sw_309_module_data_out[2] ,
    \sw_309_module_data_out[1] ,
    \sw_309_module_data_out[0] }));
 scanchain scanchain_31 (.clk_in(sw_030_clk_out),
    .clk_out(sw_031_clk_out),
    .data_in(sw_030_data_out),
    .data_out(sw_031_data_out),
    .latch_enable_in(sw_030_latch_out),
    .latch_enable_out(sw_031_latch_out),
    .scan_select_in(sw_030_scan_out),
    .scan_select_out(sw_031_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_031_module_data_in[7] ,
    \sw_031_module_data_in[6] ,
    \sw_031_module_data_in[5] ,
    \sw_031_module_data_in[4] ,
    \sw_031_module_data_in[3] ,
    \sw_031_module_data_in[2] ,
    \sw_031_module_data_in[1] ,
    \sw_031_module_data_in[0] }),
    .module_data_out({\sw_031_module_data_out[7] ,
    \sw_031_module_data_out[6] ,
    \sw_031_module_data_out[5] ,
    \sw_031_module_data_out[4] ,
    \sw_031_module_data_out[3] ,
    \sw_031_module_data_out[2] ,
    \sw_031_module_data_out[1] ,
    \sw_031_module_data_out[0] }));
 scanchain scanchain_310 (.clk_in(sw_309_clk_out),
    .clk_out(sw_310_clk_out),
    .data_in(sw_309_data_out),
    .data_out(sw_310_data_out),
    .latch_enable_in(sw_309_latch_out),
    .latch_enable_out(sw_310_latch_out),
    .scan_select_in(sw_309_scan_out),
    .scan_select_out(sw_310_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_310_module_data_in[7] ,
    \sw_310_module_data_in[6] ,
    \sw_310_module_data_in[5] ,
    \sw_310_module_data_in[4] ,
    \sw_310_module_data_in[3] ,
    \sw_310_module_data_in[2] ,
    \sw_310_module_data_in[1] ,
    \sw_310_module_data_in[0] }),
    .module_data_out({\sw_310_module_data_out[7] ,
    \sw_310_module_data_out[6] ,
    \sw_310_module_data_out[5] ,
    \sw_310_module_data_out[4] ,
    \sw_310_module_data_out[3] ,
    \sw_310_module_data_out[2] ,
    \sw_310_module_data_out[1] ,
    \sw_310_module_data_out[0] }));
 scanchain scanchain_311 (.clk_in(sw_310_clk_out),
    .clk_out(sw_311_clk_out),
    .data_in(sw_310_data_out),
    .data_out(sw_311_data_out),
    .latch_enable_in(sw_310_latch_out),
    .latch_enable_out(sw_311_latch_out),
    .scan_select_in(sw_310_scan_out),
    .scan_select_out(sw_311_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_311_module_data_in[7] ,
    \sw_311_module_data_in[6] ,
    \sw_311_module_data_in[5] ,
    \sw_311_module_data_in[4] ,
    \sw_311_module_data_in[3] ,
    \sw_311_module_data_in[2] ,
    \sw_311_module_data_in[1] ,
    \sw_311_module_data_in[0] }),
    .module_data_out({\sw_311_module_data_out[7] ,
    \sw_311_module_data_out[6] ,
    \sw_311_module_data_out[5] ,
    \sw_311_module_data_out[4] ,
    \sw_311_module_data_out[3] ,
    \sw_311_module_data_out[2] ,
    \sw_311_module_data_out[1] ,
    \sw_311_module_data_out[0] }));
 scanchain scanchain_312 (.clk_in(sw_311_clk_out),
    .clk_out(sw_312_clk_out),
    .data_in(sw_311_data_out),
    .data_out(sw_312_data_out),
    .latch_enable_in(sw_311_latch_out),
    .latch_enable_out(sw_312_latch_out),
    .scan_select_in(sw_311_scan_out),
    .scan_select_out(sw_312_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_312_module_data_in[7] ,
    \sw_312_module_data_in[6] ,
    \sw_312_module_data_in[5] ,
    \sw_312_module_data_in[4] ,
    \sw_312_module_data_in[3] ,
    \sw_312_module_data_in[2] ,
    \sw_312_module_data_in[1] ,
    \sw_312_module_data_in[0] }),
    .module_data_out({\sw_312_module_data_out[7] ,
    \sw_312_module_data_out[6] ,
    \sw_312_module_data_out[5] ,
    \sw_312_module_data_out[4] ,
    \sw_312_module_data_out[3] ,
    \sw_312_module_data_out[2] ,
    \sw_312_module_data_out[1] ,
    \sw_312_module_data_out[0] }));
 scanchain scanchain_313 (.clk_in(sw_312_clk_out),
    .clk_out(sw_313_clk_out),
    .data_in(sw_312_data_out),
    .data_out(sw_313_data_out),
    .latch_enable_in(sw_312_latch_out),
    .latch_enable_out(sw_313_latch_out),
    .scan_select_in(sw_312_scan_out),
    .scan_select_out(sw_313_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_313_module_data_in[7] ,
    \sw_313_module_data_in[6] ,
    \sw_313_module_data_in[5] ,
    \sw_313_module_data_in[4] ,
    \sw_313_module_data_in[3] ,
    \sw_313_module_data_in[2] ,
    \sw_313_module_data_in[1] ,
    \sw_313_module_data_in[0] }),
    .module_data_out({\sw_313_module_data_out[7] ,
    \sw_313_module_data_out[6] ,
    \sw_313_module_data_out[5] ,
    \sw_313_module_data_out[4] ,
    \sw_313_module_data_out[3] ,
    \sw_313_module_data_out[2] ,
    \sw_313_module_data_out[1] ,
    \sw_313_module_data_out[0] }));
 scanchain scanchain_314 (.clk_in(sw_313_clk_out),
    .clk_out(sw_314_clk_out),
    .data_in(sw_313_data_out),
    .data_out(sw_314_data_out),
    .latch_enable_in(sw_313_latch_out),
    .latch_enable_out(sw_314_latch_out),
    .scan_select_in(sw_313_scan_out),
    .scan_select_out(sw_314_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_314_module_data_in[7] ,
    \sw_314_module_data_in[6] ,
    \sw_314_module_data_in[5] ,
    \sw_314_module_data_in[4] ,
    \sw_314_module_data_in[3] ,
    \sw_314_module_data_in[2] ,
    \sw_314_module_data_in[1] ,
    \sw_314_module_data_in[0] }),
    .module_data_out({\sw_314_module_data_out[7] ,
    \sw_314_module_data_out[6] ,
    \sw_314_module_data_out[5] ,
    \sw_314_module_data_out[4] ,
    \sw_314_module_data_out[3] ,
    \sw_314_module_data_out[2] ,
    \sw_314_module_data_out[1] ,
    \sw_314_module_data_out[0] }));
 scanchain scanchain_315 (.clk_in(sw_314_clk_out),
    .clk_out(sw_315_clk_out),
    .data_in(sw_314_data_out),
    .data_out(sw_315_data_out),
    .latch_enable_in(sw_314_latch_out),
    .latch_enable_out(sw_315_latch_out),
    .scan_select_in(sw_314_scan_out),
    .scan_select_out(sw_315_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_315_module_data_in[7] ,
    \sw_315_module_data_in[6] ,
    \sw_315_module_data_in[5] ,
    \sw_315_module_data_in[4] ,
    \sw_315_module_data_in[3] ,
    \sw_315_module_data_in[2] ,
    \sw_315_module_data_in[1] ,
    \sw_315_module_data_in[0] }),
    .module_data_out({\sw_315_module_data_out[7] ,
    \sw_315_module_data_out[6] ,
    \sw_315_module_data_out[5] ,
    \sw_315_module_data_out[4] ,
    \sw_315_module_data_out[3] ,
    \sw_315_module_data_out[2] ,
    \sw_315_module_data_out[1] ,
    \sw_315_module_data_out[0] }));
 scanchain scanchain_316 (.clk_in(sw_315_clk_out),
    .clk_out(sw_316_clk_out),
    .data_in(sw_315_data_out),
    .data_out(sw_316_data_out),
    .latch_enable_in(sw_315_latch_out),
    .latch_enable_out(sw_316_latch_out),
    .scan_select_in(sw_315_scan_out),
    .scan_select_out(sw_316_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_316_module_data_in[7] ,
    \sw_316_module_data_in[6] ,
    \sw_316_module_data_in[5] ,
    \sw_316_module_data_in[4] ,
    \sw_316_module_data_in[3] ,
    \sw_316_module_data_in[2] ,
    \sw_316_module_data_in[1] ,
    \sw_316_module_data_in[0] }),
    .module_data_out({\sw_316_module_data_out[7] ,
    \sw_316_module_data_out[6] ,
    \sw_316_module_data_out[5] ,
    \sw_316_module_data_out[4] ,
    \sw_316_module_data_out[3] ,
    \sw_316_module_data_out[2] ,
    \sw_316_module_data_out[1] ,
    \sw_316_module_data_out[0] }));
 scanchain scanchain_317 (.clk_in(sw_316_clk_out),
    .clk_out(sw_317_clk_out),
    .data_in(sw_316_data_out),
    .data_out(sw_317_data_out),
    .latch_enable_in(sw_316_latch_out),
    .latch_enable_out(sw_317_latch_out),
    .scan_select_in(sw_316_scan_out),
    .scan_select_out(sw_317_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_317_module_data_in[7] ,
    \sw_317_module_data_in[6] ,
    \sw_317_module_data_in[5] ,
    \sw_317_module_data_in[4] ,
    \sw_317_module_data_in[3] ,
    \sw_317_module_data_in[2] ,
    \sw_317_module_data_in[1] ,
    \sw_317_module_data_in[0] }),
    .module_data_out({\sw_317_module_data_out[7] ,
    \sw_317_module_data_out[6] ,
    \sw_317_module_data_out[5] ,
    \sw_317_module_data_out[4] ,
    \sw_317_module_data_out[3] ,
    \sw_317_module_data_out[2] ,
    \sw_317_module_data_out[1] ,
    \sw_317_module_data_out[0] }));
 scanchain scanchain_318 (.clk_in(sw_317_clk_out),
    .clk_out(sw_318_clk_out),
    .data_in(sw_317_data_out),
    .data_out(sw_318_data_out),
    .latch_enable_in(sw_317_latch_out),
    .latch_enable_out(sw_318_latch_out),
    .scan_select_in(sw_317_scan_out),
    .scan_select_out(sw_318_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_318_module_data_in[7] ,
    \sw_318_module_data_in[6] ,
    \sw_318_module_data_in[5] ,
    \sw_318_module_data_in[4] ,
    \sw_318_module_data_in[3] ,
    \sw_318_module_data_in[2] ,
    \sw_318_module_data_in[1] ,
    \sw_318_module_data_in[0] }),
    .module_data_out({\sw_318_module_data_out[7] ,
    \sw_318_module_data_out[6] ,
    \sw_318_module_data_out[5] ,
    \sw_318_module_data_out[4] ,
    \sw_318_module_data_out[3] ,
    \sw_318_module_data_out[2] ,
    \sw_318_module_data_out[1] ,
    \sw_318_module_data_out[0] }));
 scanchain scanchain_319 (.clk_in(sw_318_clk_out),
    .clk_out(sw_319_clk_out),
    .data_in(sw_318_data_out),
    .data_out(sw_319_data_out),
    .latch_enable_in(sw_318_latch_out),
    .latch_enable_out(sw_319_latch_out),
    .scan_select_in(sw_318_scan_out),
    .scan_select_out(sw_319_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_319_module_data_in[7] ,
    \sw_319_module_data_in[6] ,
    \sw_319_module_data_in[5] ,
    \sw_319_module_data_in[4] ,
    \sw_319_module_data_in[3] ,
    \sw_319_module_data_in[2] ,
    \sw_319_module_data_in[1] ,
    \sw_319_module_data_in[0] }),
    .module_data_out({\sw_319_module_data_out[7] ,
    \sw_319_module_data_out[6] ,
    \sw_319_module_data_out[5] ,
    \sw_319_module_data_out[4] ,
    \sw_319_module_data_out[3] ,
    \sw_319_module_data_out[2] ,
    \sw_319_module_data_out[1] ,
    \sw_319_module_data_out[0] }));
 scanchain scanchain_32 (.clk_in(sw_031_clk_out),
    .clk_out(sw_032_clk_out),
    .data_in(sw_031_data_out),
    .data_out(sw_032_data_out),
    .latch_enable_in(sw_031_latch_out),
    .latch_enable_out(sw_032_latch_out),
    .scan_select_in(sw_031_scan_out),
    .scan_select_out(sw_032_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_032_module_data_in[7] ,
    \sw_032_module_data_in[6] ,
    \sw_032_module_data_in[5] ,
    \sw_032_module_data_in[4] ,
    \sw_032_module_data_in[3] ,
    \sw_032_module_data_in[2] ,
    \sw_032_module_data_in[1] ,
    \sw_032_module_data_in[0] }),
    .module_data_out({\sw_032_module_data_out[7] ,
    \sw_032_module_data_out[6] ,
    \sw_032_module_data_out[5] ,
    \sw_032_module_data_out[4] ,
    \sw_032_module_data_out[3] ,
    \sw_032_module_data_out[2] ,
    \sw_032_module_data_out[1] ,
    \sw_032_module_data_out[0] }));
 scanchain scanchain_320 (.clk_in(sw_319_clk_out),
    .clk_out(sw_320_clk_out),
    .data_in(sw_319_data_out),
    .data_out(sw_320_data_out),
    .latch_enable_in(sw_319_latch_out),
    .latch_enable_out(sw_320_latch_out),
    .scan_select_in(sw_319_scan_out),
    .scan_select_out(sw_320_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_320_module_data_in[7] ,
    \sw_320_module_data_in[6] ,
    \sw_320_module_data_in[5] ,
    \sw_320_module_data_in[4] ,
    \sw_320_module_data_in[3] ,
    \sw_320_module_data_in[2] ,
    \sw_320_module_data_in[1] ,
    \sw_320_module_data_in[0] }),
    .module_data_out({\sw_320_module_data_out[7] ,
    \sw_320_module_data_out[6] ,
    \sw_320_module_data_out[5] ,
    \sw_320_module_data_out[4] ,
    \sw_320_module_data_out[3] ,
    \sw_320_module_data_out[2] ,
    \sw_320_module_data_out[1] ,
    \sw_320_module_data_out[0] }));
 scanchain scanchain_321 (.clk_in(sw_320_clk_out),
    .clk_out(sw_321_clk_out),
    .data_in(sw_320_data_out),
    .data_out(sw_321_data_out),
    .latch_enable_in(sw_320_latch_out),
    .latch_enable_out(sw_321_latch_out),
    .scan_select_in(sw_320_scan_out),
    .scan_select_out(sw_321_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_321_module_data_in[7] ,
    \sw_321_module_data_in[6] ,
    \sw_321_module_data_in[5] ,
    \sw_321_module_data_in[4] ,
    \sw_321_module_data_in[3] ,
    \sw_321_module_data_in[2] ,
    \sw_321_module_data_in[1] ,
    \sw_321_module_data_in[0] }),
    .module_data_out({\sw_321_module_data_out[7] ,
    \sw_321_module_data_out[6] ,
    \sw_321_module_data_out[5] ,
    \sw_321_module_data_out[4] ,
    \sw_321_module_data_out[3] ,
    \sw_321_module_data_out[2] ,
    \sw_321_module_data_out[1] ,
    \sw_321_module_data_out[0] }));
 scanchain scanchain_322 (.clk_in(sw_321_clk_out),
    .clk_out(sw_322_clk_out),
    .data_in(sw_321_data_out),
    .data_out(sw_322_data_out),
    .latch_enable_in(sw_321_latch_out),
    .latch_enable_out(sw_322_latch_out),
    .scan_select_in(sw_321_scan_out),
    .scan_select_out(sw_322_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_322_module_data_in[7] ,
    \sw_322_module_data_in[6] ,
    \sw_322_module_data_in[5] ,
    \sw_322_module_data_in[4] ,
    \sw_322_module_data_in[3] ,
    \sw_322_module_data_in[2] ,
    \sw_322_module_data_in[1] ,
    \sw_322_module_data_in[0] }),
    .module_data_out({\sw_322_module_data_out[7] ,
    \sw_322_module_data_out[6] ,
    \sw_322_module_data_out[5] ,
    \sw_322_module_data_out[4] ,
    \sw_322_module_data_out[3] ,
    \sw_322_module_data_out[2] ,
    \sw_322_module_data_out[1] ,
    \sw_322_module_data_out[0] }));
 scanchain scanchain_323 (.clk_in(sw_322_clk_out),
    .clk_out(sw_323_clk_out),
    .data_in(sw_322_data_out),
    .data_out(sw_323_data_out),
    .latch_enable_in(sw_322_latch_out),
    .latch_enable_out(sw_323_latch_out),
    .scan_select_in(sw_322_scan_out),
    .scan_select_out(sw_323_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_323_module_data_in[7] ,
    \sw_323_module_data_in[6] ,
    \sw_323_module_data_in[5] ,
    \sw_323_module_data_in[4] ,
    \sw_323_module_data_in[3] ,
    \sw_323_module_data_in[2] ,
    \sw_323_module_data_in[1] ,
    \sw_323_module_data_in[0] }),
    .module_data_out({\sw_323_module_data_out[7] ,
    \sw_323_module_data_out[6] ,
    \sw_323_module_data_out[5] ,
    \sw_323_module_data_out[4] ,
    \sw_323_module_data_out[3] ,
    \sw_323_module_data_out[2] ,
    \sw_323_module_data_out[1] ,
    \sw_323_module_data_out[0] }));
 scanchain scanchain_324 (.clk_in(sw_323_clk_out),
    .clk_out(sw_324_clk_out),
    .data_in(sw_323_data_out),
    .data_out(sw_324_data_out),
    .latch_enable_in(sw_323_latch_out),
    .latch_enable_out(sw_324_latch_out),
    .scan_select_in(sw_323_scan_out),
    .scan_select_out(sw_324_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_324_module_data_in[7] ,
    \sw_324_module_data_in[6] ,
    \sw_324_module_data_in[5] ,
    \sw_324_module_data_in[4] ,
    \sw_324_module_data_in[3] ,
    \sw_324_module_data_in[2] ,
    \sw_324_module_data_in[1] ,
    \sw_324_module_data_in[0] }),
    .module_data_out({\sw_324_module_data_out[7] ,
    \sw_324_module_data_out[6] ,
    \sw_324_module_data_out[5] ,
    \sw_324_module_data_out[4] ,
    \sw_324_module_data_out[3] ,
    \sw_324_module_data_out[2] ,
    \sw_324_module_data_out[1] ,
    \sw_324_module_data_out[0] }));
 scanchain scanchain_325 (.clk_in(sw_324_clk_out),
    .clk_out(sw_325_clk_out),
    .data_in(sw_324_data_out),
    .data_out(sw_325_data_out),
    .latch_enable_in(sw_324_latch_out),
    .latch_enable_out(sw_325_latch_out),
    .scan_select_in(sw_324_scan_out),
    .scan_select_out(sw_325_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_325_module_data_in[7] ,
    \sw_325_module_data_in[6] ,
    \sw_325_module_data_in[5] ,
    \sw_325_module_data_in[4] ,
    \sw_325_module_data_in[3] ,
    \sw_325_module_data_in[2] ,
    \sw_325_module_data_in[1] ,
    \sw_325_module_data_in[0] }),
    .module_data_out({\sw_325_module_data_out[7] ,
    \sw_325_module_data_out[6] ,
    \sw_325_module_data_out[5] ,
    \sw_325_module_data_out[4] ,
    \sw_325_module_data_out[3] ,
    \sw_325_module_data_out[2] ,
    \sw_325_module_data_out[1] ,
    \sw_325_module_data_out[0] }));
 scanchain scanchain_326 (.clk_in(sw_325_clk_out),
    .clk_out(sw_326_clk_out),
    .data_in(sw_325_data_out),
    .data_out(sw_326_data_out),
    .latch_enable_in(sw_325_latch_out),
    .latch_enable_out(sw_326_latch_out),
    .scan_select_in(sw_325_scan_out),
    .scan_select_out(sw_326_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_326_module_data_in[7] ,
    \sw_326_module_data_in[6] ,
    \sw_326_module_data_in[5] ,
    \sw_326_module_data_in[4] ,
    \sw_326_module_data_in[3] ,
    \sw_326_module_data_in[2] ,
    \sw_326_module_data_in[1] ,
    \sw_326_module_data_in[0] }),
    .module_data_out({\sw_326_module_data_out[7] ,
    \sw_326_module_data_out[6] ,
    \sw_326_module_data_out[5] ,
    \sw_326_module_data_out[4] ,
    \sw_326_module_data_out[3] ,
    \sw_326_module_data_out[2] ,
    \sw_326_module_data_out[1] ,
    \sw_326_module_data_out[0] }));
 scanchain scanchain_327 (.clk_in(sw_326_clk_out),
    .clk_out(sw_327_clk_out),
    .data_in(sw_326_data_out),
    .data_out(sw_327_data_out),
    .latch_enable_in(sw_326_latch_out),
    .latch_enable_out(sw_327_latch_out),
    .scan_select_in(sw_326_scan_out),
    .scan_select_out(sw_327_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_327_module_data_in[7] ,
    \sw_327_module_data_in[6] ,
    \sw_327_module_data_in[5] ,
    \sw_327_module_data_in[4] ,
    \sw_327_module_data_in[3] ,
    \sw_327_module_data_in[2] ,
    \sw_327_module_data_in[1] ,
    \sw_327_module_data_in[0] }),
    .module_data_out({\sw_327_module_data_out[7] ,
    \sw_327_module_data_out[6] ,
    \sw_327_module_data_out[5] ,
    \sw_327_module_data_out[4] ,
    \sw_327_module_data_out[3] ,
    \sw_327_module_data_out[2] ,
    \sw_327_module_data_out[1] ,
    \sw_327_module_data_out[0] }));
 scanchain scanchain_328 (.clk_in(sw_327_clk_out),
    .clk_out(sw_328_clk_out),
    .data_in(sw_327_data_out),
    .data_out(sw_328_data_out),
    .latch_enable_in(sw_327_latch_out),
    .latch_enable_out(sw_328_latch_out),
    .scan_select_in(sw_327_scan_out),
    .scan_select_out(sw_328_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_328_module_data_in[7] ,
    \sw_328_module_data_in[6] ,
    \sw_328_module_data_in[5] ,
    \sw_328_module_data_in[4] ,
    \sw_328_module_data_in[3] ,
    \sw_328_module_data_in[2] ,
    \sw_328_module_data_in[1] ,
    \sw_328_module_data_in[0] }),
    .module_data_out({\sw_328_module_data_out[7] ,
    \sw_328_module_data_out[6] ,
    \sw_328_module_data_out[5] ,
    \sw_328_module_data_out[4] ,
    \sw_328_module_data_out[3] ,
    \sw_328_module_data_out[2] ,
    \sw_328_module_data_out[1] ,
    \sw_328_module_data_out[0] }));
 scanchain scanchain_329 (.clk_in(sw_328_clk_out),
    .clk_out(sw_329_clk_out),
    .data_in(sw_328_data_out),
    .data_out(sw_329_data_out),
    .latch_enable_in(sw_328_latch_out),
    .latch_enable_out(sw_329_latch_out),
    .scan_select_in(sw_328_scan_out),
    .scan_select_out(sw_329_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_329_module_data_in[7] ,
    \sw_329_module_data_in[6] ,
    \sw_329_module_data_in[5] ,
    \sw_329_module_data_in[4] ,
    \sw_329_module_data_in[3] ,
    \sw_329_module_data_in[2] ,
    \sw_329_module_data_in[1] ,
    \sw_329_module_data_in[0] }),
    .module_data_out({\sw_329_module_data_out[7] ,
    \sw_329_module_data_out[6] ,
    \sw_329_module_data_out[5] ,
    \sw_329_module_data_out[4] ,
    \sw_329_module_data_out[3] ,
    \sw_329_module_data_out[2] ,
    \sw_329_module_data_out[1] ,
    \sw_329_module_data_out[0] }));
 scanchain scanchain_33 (.clk_in(sw_032_clk_out),
    .clk_out(sw_033_clk_out),
    .data_in(sw_032_data_out),
    .data_out(sw_033_data_out),
    .latch_enable_in(sw_032_latch_out),
    .latch_enable_out(sw_033_latch_out),
    .scan_select_in(sw_032_scan_out),
    .scan_select_out(sw_033_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_033_module_data_in[7] ,
    \sw_033_module_data_in[6] ,
    \sw_033_module_data_in[5] ,
    \sw_033_module_data_in[4] ,
    \sw_033_module_data_in[3] ,
    \sw_033_module_data_in[2] ,
    \sw_033_module_data_in[1] ,
    \sw_033_module_data_in[0] }),
    .module_data_out({\sw_033_module_data_out[7] ,
    \sw_033_module_data_out[6] ,
    \sw_033_module_data_out[5] ,
    \sw_033_module_data_out[4] ,
    \sw_033_module_data_out[3] ,
    \sw_033_module_data_out[2] ,
    \sw_033_module_data_out[1] ,
    \sw_033_module_data_out[0] }));
 scanchain scanchain_330 (.clk_in(sw_329_clk_out),
    .clk_out(sw_330_clk_out),
    .data_in(sw_329_data_out),
    .data_out(sw_330_data_out),
    .latch_enable_in(sw_329_latch_out),
    .latch_enable_out(sw_330_latch_out),
    .scan_select_in(sw_329_scan_out),
    .scan_select_out(sw_330_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_330_module_data_in[7] ,
    \sw_330_module_data_in[6] ,
    \sw_330_module_data_in[5] ,
    \sw_330_module_data_in[4] ,
    \sw_330_module_data_in[3] ,
    \sw_330_module_data_in[2] ,
    \sw_330_module_data_in[1] ,
    \sw_330_module_data_in[0] }),
    .module_data_out({\sw_330_module_data_out[7] ,
    \sw_330_module_data_out[6] ,
    \sw_330_module_data_out[5] ,
    \sw_330_module_data_out[4] ,
    \sw_330_module_data_out[3] ,
    \sw_330_module_data_out[2] ,
    \sw_330_module_data_out[1] ,
    \sw_330_module_data_out[0] }));
 scanchain scanchain_331 (.clk_in(sw_330_clk_out),
    .clk_out(sw_331_clk_out),
    .data_in(sw_330_data_out),
    .data_out(sw_331_data_out),
    .latch_enable_in(sw_330_latch_out),
    .latch_enable_out(sw_331_latch_out),
    .scan_select_in(sw_330_scan_out),
    .scan_select_out(sw_331_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_331_module_data_in[7] ,
    \sw_331_module_data_in[6] ,
    \sw_331_module_data_in[5] ,
    \sw_331_module_data_in[4] ,
    \sw_331_module_data_in[3] ,
    \sw_331_module_data_in[2] ,
    \sw_331_module_data_in[1] ,
    \sw_331_module_data_in[0] }),
    .module_data_out({\sw_331_module_data_out[7] ,
    \sw_331_module_data_out[6] ,
    \sw_331_module_data_out[5] ,
    \sw_331_module_data_out[4] ,
    \sw_331_module_data_out[3] ,
    \sw_331_module_data_out[2] ,
    \sw_331_module_data_out[1] ,
    \sw_331_module_data_out[0] }));
 scanchain scanchain_332 (.clk_in(sw_331_clk_out),
    .clk_out(sw_332_clk_out),
    .data_in(sw_331_data_out),
    .data_out(sw_332_data_out),
    .latch_enable_in(sw_331_latch_out),
    .latch_enable_out(sw_332_latch_out),
    .scan_select_in(sw_331_scan_out),
    .scan_select_out(sw_332_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_332_module_data_in[7] ,
    \sw_332_module_data_in[6] ,
    \sw_332_module_data_in[5] ,
    \sw_332_module_data_in[4] ,
    \sw_332_module_data_in[3] ,
    \sw_332_module_data_in[2] ,
    \sw_332_module_data_in[1] ,
    \sw_332_module_data_in[0] }),
    .module_data_out({\sw_332_module_data_out[7] ,
    \sw_332_module_data_out[6] ,
    \sw_332_module_data_out[5] ,
    \sw_332_module_data_out[4] ,
    \sw_332_module_data_out[3] ,
    \sw_332_module_data_out[2] ,
    \sw_332_module_data_out[1] ,
    \sw_332_module_data_out[0] }));
 scanchain scanchain_333 (.clk_in(sw_332_clk_out),
    .clk_out(sw_333_clk_out),
    .data_in(sw_332_data_out),
    .data_out(sw_333_data_out),
    .latch_enable_in(sw_332_latch_out),
    .latch_enable_out(sw_333_latch_out),
    .scan_select_in(sw_332_scan_out),
    .scan_select_out(sw_333_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_333_module_data_in[7] ,
    \sw_333_module_data_in[6] ,
    \sw_333_module_data_in[5] ,
    \sw_333_module_data_in[4] ,
    \sw_333_module_data_in[3] ,
    \sw_333_module_data_in[2] ,
    \sw_333_module_data_in[1] ,
    \sw_333_module_data_in[0] }),
    .module_data_out({\sw_333_module_data_out[7] ,
    \sw_333_module_data_out[6] ,
    \sw_333_module_data_out[5] ,
    \sw_333_module_data_out[4] ,
    \sw_333_module_data_out[3] ,
    \sw_333_module_data_out[2] ,
    \sw_333_module_data_out[1] ,
    \sw_333_module_data_out[0] }));
 scanchain scanchain_334 (.clk_in(sw_333_clk_out),
    .clk_out(sw_334_clk_out),
    .data_in(sw_333_data_out),
    .data_out(sw_334_data_out),
    .latch_enable_in(sw_333_latch_out),
    .latch_enable_out(sw_334_latch_out),
    .scan_select_in(sw_333_scan_out),
    .scan_select_out(sw_334_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_334_module_data_in[7] ,
    \sw_334_module_data_in[6] ,
    \sw_334_module_data_in[5] ,
    \sw_334_module_data_in[4] ,
    \sw_334_module_data_in[3] ,
    \sw_334_module_data_in[2] ,
    \sw_334_module_data_in[1] ,
    \sw_334_module_data_in[0] }),
    .module_data_out({\sw_334_module_data_out[7] ,
    \sw_334_module_data_out[6] ,
    \sw_334_module_data_out[5] ,
    \sw_334_module_data_out[4] ,
    \sw_334_module_data_out[3] ,
    \sw_334_module_data_out[2] ,
    \sw_334_module_data_out[1] ,
    \sw_334_module_data_out[0] }));
 scanchain scanchain_335 (.clk_in(sw_334_clk_out),
    .clk_out(sw_335_clk_out),
    .data_in(sw_334_data_out),
    .data_out(sw_335_data_out),
    .latch_enable_in(sw_334_latch_out),
    .latch_enable_out(sw_335_latch_out),
    .scan_select_in(sw_334_scan_out),
    .scan_select_out(sw_335_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_335_module_data_in[7] ,
    \sw_335_module_data_in[6] ,
    \sw_335_module_data_in[5] ,
    \sw_335_module_data_in[4] ,
    \sw_335_module_data_in[3] ,
    \sw_335_module_data_in[2] ,
    \sw_335_module_data_in[1] ,
    \sw_335_module_data_in[0] }),
    .module_data_out({\sw_335_module_data_out[7] ,
    \sw_335_module_data_out[6] ,
    \sw_335_module_data_out[5] ,
    \sw_335_module_data_out[4] ,
    \sw_335_module_data_out[3] ,
    \sw_335_module_data_out[2] ,
    \sw_335_module_data_out[1] ,
    \sw_335_module_data_out[0] }));
 scanchain scanchain_336 (.clk_in(sw_335_clk_out),
    .clk_out(sw_336_clk_out),
    .data_in(sw_335_data_out),
    .data_out(sw_336_data_out),
    .latch_enable_in(sw_335_latch_out),
    .latch_enable_out(sw_336_latch_out),
    .scan_select_in(sw_335_scan_out),
    .scan_select_out(sw_336_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_336_module_data_in[7] ,
    \sw_336_module_data_in[6] ,
    \sw_336_module_data_in[5] ,
    \sw_336_module_data_in[4] ,
    \sw_336_module_data_in[3] ,
    \sw_336_module_data_in[2] ,
    \sw_336_module_data_in[1] ,
    \sw_336_module_data_in[0] }),
    .module_data_out({\sw_336_module_data_out[7] ,
    \sw_336_module_data_out[6] ,
    \sw_336_module_data_out[5] ,
    \sw_336_module_data_out[4] ,
    \sw_336_module_data_out[3] ,
    \sw_336_module_data_out[2] ,
    \sw_336_module_data_out[1] ,
    \sw_336_module_data_out[0] }));
 scanchain scanchain_337 (.clk_in(sw_336_clk_out),
    .clk_out(sw_337_clk_out),
    .data_in(sw_336_data_out),
    .data_out(sw_337_data_out),
    .latch_enable_in(sw_336_latch_out),
    .latch_enable_out(sw_337_latch_out),
    .scan_select_in(sw_336_scan_out),
    .scan_select_out(sw_337_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_337_module_data_in[7] ,
    \sw_337_module_data_in[6] ,
    \sw_337_module_data_in[5] ,
    \sw_337_module_data_in[4] ,
    \sw_337_module_data_in[3] ,
    \sw_337_module_data_in[2] ,
    \sw_337_module_data_in[1] ,
    \sw_337_module_data_in[0] }),
    .module_data_out({\sw_337_module_data_out[7] ,
    \sw_337_module_data_out[6] ,
    \sw_337_module_data_out[5] ,
    \sw_337_module_data_out[4] ,
    \sw_337_module_data_out[3] ,
    \sw_337_module_data_out[2] ,
    \sw_337_module_data_out[1] ,
    \sw_337_module_data_out[0] }));
 scanchain scanchain_338 (.clk_in(sw_337_clk_out),
    .clk_out(sw_338_clk_out),
    .data_in(sw_337_data_out),
    .data_out(sw_338_data_out),
    .latch_enable_in(sw_337_latch_out),
    .latch_enable_out(sw_338_latch_out),
    .scan_select_in(sw_337_scan_out),
    .scan_select_out(sw_338_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_338_module_data_in[7] ,
    \sw_338_module_data_in[6] ,
    \sw_338_module_data_in[5] ,
    \sw_338_module_data_in[4] ,
    \sw_338_module_data_in[3] ,
    \sw_338_module_data_in[2] ,
    \sw_338_module_data_in[1] ,
    \sw_338_module_data_in[0] }),
    .module_data_out({\sw_338_module_data_out[7] ,
    \sw_338_module_data_out[6] ,
    \sw_338_module_data_out[5] ,
    \sw_338_module_data_out[4] ,
    \sw_338_module_data_out[3] ,
    \sw_338_module_data_out[2] ,
    \sw_338_module_data_out[1] ,
    \sw_338_module_data_out[0] }));
 scanchain scanchain_339 (.clk_in(sw_338_clk_out),
    .clk_out(sw_339_clk_out),
    .data_in(sw_338_data_out),
    .data_out(sw_339_data_out),
    .latch_enable_in(sw_338_latch_out),
    .latch_enable_out(sw_339_latch_out),
    .scan_select_in(sw_338_scan_out),
    .scan_select_out(sw_339_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_339_module_data_in[7] ,
    \sw_339_module_data_in[6] ,
    \sw_339_module_data_in[5] ,
    \sw_339_module_data_in[4] ,
    \sw_339_module_data_in[3] ,
    \sw_339_module_data_in[2] ,
    \sw_339_module_data_in[1] ,
    \sw_339_module_data_in[0] }),
    .module_data_out({\sw_339_module_data_out[7] ,
    \sw_339_module_data_out[6] ,
    \sw_339_module_data_out[5] ,
    \sw_339_module_data_out[4] ,
    \sw_339_module_data_out[3] ,
    \sw_339_module_data_out[2] ,
    \sw_339_module_data_out[1] ,
    \sw_339_module_data_out[0] }));
 scanchain scanchain_34 (.clk_in(sw_033_clk_out),
    .clk_out(sw_034_clk_out),
    .data_in(sw_033_data_out),
    .data_out(sw_034_data_out),
    .latch_enable_in(sw_033_latch_out),
    .latch_enable_out(sw_034_latch_out),
    .scan_select_in(sw_033_scan_out),
    .scan_select_out(sw_034_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_034_module_data_in[7] ,
    \sw_034_module_data_in[6] ,
    \sw_034_module_data_in[5] ,
    \sw_034_module_data_in[4] ,
    \sw_034_module_data_in[3] ,
    \sw_034_module_data_in[2] ,
    \sw_034_module_data_in[1] ,
    \sw_034_module_data_in[0] }),
    .module_data_out({\sw_034_module_data_out[7] ,
    \sw_034_module_data_out[6] ,
    \sw_034_module_data_out[5] ,
    \sw_034_module_data_out[4] ,
    \sw_034_module_data_out[3] ,
    \sw_034_module_data_out[2] ,
    \sw_034_module_data_out[1] ,
    \sw_034_module_data_out[0] }));
 scanchain scanchain_340 (.clk_in(sw_339_clk_out),
    .clk_out(sw_340_clk_out),
    .data_in(sw_339_data_out),
    .data_out(sw_340_data_out),
    .latch_enable_in(sw_339_latch_out),
    .latch_enable_out(sw_340_latch_out),
    .scan_select_in(sw_339_scan_out),
    .scan_select_out(sw_340_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_340_module_data_in[7] ,
    \sw_340_module_data_in[6] ,
    \sw_340_module_data_in[5] ,
    \sw_340_module_data_in[4] ,
    \sw_340_module_data_in[3] ,
    \sw_340_module_data_in[2] ,
    \sw_340_module_data_in[1] ,
    \sw_340_module_data_in[0] }),
    .module_data_out({\sw_340_module_data_out[7] ,
    \sw_340_module_data_out[6] ,
    \sw_340_module_data_out[5] ,
    \sw_340_module_data_out[4] ,
    \sw_340_module_data_out[3] ,
    \sw_340_module_data_out[2] ,
    \sw_340_module_data_out[1] ,
    \sw_340_module_data_out[0] }));
 scanchain scanchain_341 (.clk_in(sw_340_clk_out),
    .clk_out(sw_341_clk_out),
    .data_in(sw_340_data_out),
    .data_out(sw_341_data_out),
    .latch_enable_in(sw_340_latch_out),
    .latch_enable_out(sw_341_latch_out),
    .scan_select_in(sw_340_scan_out),
    .scan_select_out(sw_341_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_341_module_data_in[7] ,
    \sw_341_module_data_in[6] ,
    \sw_341_module_data_in[5] ,
    \sw_341_module_data_in[4] ,
    \sw_341_module_data_in[3] ,
    \sw_341_module_data_in[2] ,
    \sw_341_module_data_in[1] ,
    \sw_341_module_data_in[0] }),
    .module_data_out({\sw_341_module_data_out[7] ,
    \sw_341_module_data_out[6] ,
    \sw_341_module_data_out[5] ,
    \sw_341_module_data_out[4] ,
    \sw_341_module_data_out[3] ,
    \sw_341_module_data_out[2] ,
    \sw_341_module_data_out[1] ,
    \sw_341_module_data_out[0] }));
 scanchain scanchain_342 (.clk_in(sw_341_clk_out),
    .clk_out(sw_342_clk_out),
    .data_in(sw_341_data_out),
    .data_out(sw_342_data_out),
    .latch_enable_in(sw_341_latch_out),
    .latch_enable_out(sw_342_latch_out),
    .scan_select_in(sw_341_scan_out),
    .scan_select_out(sw_342_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_342_module_data_in[7] ,
    \sw_342_module_data_in[6] ,
    \sw_342_module_data_in[5] ,
    \sw_342_module_data_in[4] ,
    \sw_342_module_data_in[3] ,
    \sw_342_module_data_in[2] ,
    \sw_342_module_data_in[1] ,
    \sw_342_module_data_in[0] }),
    .module_data_out({\sw_342_module_data_out[7] ,
    \sw_342_module_data_out[6] ,
    \sw_342_module_data_out[5] ,
    \sw_342_module_data_out[4] ,
    \sw_342_module_data_out[3] ,
    \sw_342_module_data_out[2] ,
    \sw_342_module_data_out[1] ,
    \sw_342_module_data_out[0] }));
 scanchain scanchain_343 (.clk_in(sw_342_clk_out),
    .clk_out(sw_343_clk_out),
    .data_in(sw_342_data_out),
    .data_out(sw_343_data_out),
    .latch_enable_in(sw_342_latch_out),
    .latch_enable_out(sw_343_latch_out),
    .scan_select_in(sw_342_scan_out),
    .scan_select_out(sw_343_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_343_module_data_in[7] ,
    \sw_343_module_data_in[6] ,
    \sw_343_module_data_in[5] ,
    \sw_343_module_data_in[4] ,
    \sw_343_module_data_in[3] ,
    \sw_343_module_data_in[2] ,
    \sw_343_module_data_in[1] ,
    \sw_343_module_data_in[0] }),
    .module_data_out({\sw_343_module_data_out[7] ,
    \sw_343_module_data_out[6] ,
    \sw_343_module_data_out[5] ,
    \sw_343_module_data_out[4] ,
    \sw_343_module_data_out[3] ,
    \sw_343_module_data_out[2] ,
    \sw_343_module_data_out[1] ,
    \sw_343_module_data_out[0] }));
 scanchain scanchain_344 (.clk_in(sw_343_clk_out),
    .clk_out(sw_344_clk_out),
    .data_in(sw_343_data_out),
    .data_out(sw_344_data_out),
    .latch_enable_in(sw_343_latch_out),
    .latch_enable_out(sw_344_latch_out),
    .scan_select_in(sw_343_scan_out),
    .scan_select_out(sw_344_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_344_module_data_in[7] ,
    \sw_344_module_data_in[6] ,
    \sw_344_module_data_in[5] ,
    \sw_344_module_data_in[4] ,
    \sw_344_module_data_in[3] ,
    \sw_344_module_data_in[2] ,
    \sw_344_module_data_in[1] ,
    \sw_344_module_data_in[0] }),
    .module_data_out({\sw_344_module_data_out[7] ,
    \sw_344_module_data_out[6] ,
    \sw_344_module_data_out[5] ,
    \sw_344_module_data_out[4] ,
    \sw_344_module_data_out[3] ,
    \sw_344_module_data_out[2] ,
    \sw_344_module_data_out[1] ,
    \sw_344_module_data_out[0] }));
 scanchain scanchain_345 (.clk_in(sw_344_clk_out),
    .clk_out(sw_345_clk_out),
    .data_in(sw_344_data_out),
    .data_out(sw_345_data_out),
    .latch_enable_in(sw_344_latch_out),
    .latch_enable_out(sw_345_latch_out),
    .scan_select_in(sw_344_scan_out),
    .scan_select_out(sw_345_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_345_module_data_in[7] ,
    \sw_345_module_data_in[6] ,
    \sw_345_module_data_in[5] ,
    \sw_345_module_data_in[4] ,
    \sw_345_module_data_in[3] ,
    \sw_345_module_data_in[2] ,
    \sw_345_module_data_in[1] ,
    \sw_345_module_data_in[0] }),
    .module_data_out({\sw_345_module_data_out[7] ,
    \sw_345_module_data_out[6] ,
    \sw_345_module_data_out[5] ,
    \sw_345_module_data_out[4] ,
    \sw_345_module_data_out[3] ,
    \sw_345_module_data_out[2] ,
    \sw_345_module_data_out[1] ,
    \sw_345_module_data_out[0] }));
 scanchain scanchain_346 (.clk_in(sw_345_clk_out),
    .clk_out(sw_346_clk_out),
    .data_in(sw_345_data_out),
    .data_out(sw_346_data_out),
    .latch_enable_in(sw_345_latch_out),
    .latch_enable_out(sw_346_latch_out),
    .scan_select_in(sw_345_scan_out),
    .scan_select_out(sw_346_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_346_module_data_in[7] ,
    \sw_346_module_data_in[6] ,
    \sw_346_module_data_in[5] ,
    \sw_346_module_data_in[4] ,
    \sw_346_module_data_in[3] ,
    \sw_346_module_data_in[2] ,
    \sw_346_module_data_in[1] ,
    \sw_346_module_data_in[0] }),
    .module_data_out({\sw_346_module_data_out[7] ,
    \sw_346_module_data_out[6] ,
    \sw_346_module_data_out[5] ,
    \sw_346_module_data_out[4] ,
    \sw_346_module_data_out[3] ,
    \sw_346_module_data_out[2] ,
    \sw_346_module_data_out[1] ,
    \sw_346_module_data_out[0] }));
 scanchain scanchain_347 (.clk_in(sw_346_clk_out),
    .clk_out(sw_347_clk_out),
    .data_in(sw_346_data_out),
    .data_out(sw_347_data_out),
    .latch_enable_in(sw_346_latch_out),
    .latch_enable_out(sw_347_latch_out),
    .scan_select_in(sw_346_scan_out),
    .scan_select_out(sw_347_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_347_module_data_in[7] ,
    \sw_347_module_data_in[6] ,
    \sw_347_module_data_in[5] ,
    \sw_347_module_data_in[4] ,
    \sw_347_module_data_in[3] ,
    \sw_347_module_data_in[2] ,
    \sw_347_module_data_in[1] ,
    \sw_347_module_data_in[0] }),
    .module_data_out({\sw_347_module_data_out[7] ,
    \sw_347_module_data_out[6] ,
    \sw_347_module_data_out[5] ,
    \sw_347_module_data_out[4] ,
    \sw_347_module_data_out[3] ,
    \sw_347_module_data_out[2] ,
    \sw_347_module_data_out[1] ,
    \sw_347_module_data_out[0] }));
 scanchain scanchain_348 (.clk_in(sw_347_clk_out),
    .clk_out(sw_348_clk_out),
    .data_in(sw_347_data_out),
    .data_out(sw_348_data_out),
    .latch_enable_in(sw_347_latch_out),
    .latch_enable_out(sw_348_latch_out),
    .scan_select_in(sw_347_scan_out),
    .scan_select_out(sw_348_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_348_module_data_in[7] ,
    \sw_348_module_data_in[6] ,
    \sw_348_module_data_in[5] ,
    \sw_348_module_data_in[4] ,
    \sw_348_module_data_in[3] ,
    \sw_348_module_data_in[2] ,
    \sw_348_module_data_in[1] ,
    \sw_348_module_data_in[0] }),
    .module_data_out({\sw_348_module_data_out[7] ,
    \sw_348_module_data_out[6] ,
    \sw_348_module_data_out[5] ,
    \sw_348_module_data_out[4] ,
    \sw_348_module_data_out[3] ,
    \sw_348_module_data_out[2] ,
    \sw_348_module_data_out[1] ,
    \sw_348_module_data_out[0] }));
 scanchain scanchain_349 (.clk_in(sw_348_clk_out),
    .clk_out(sw_349_clk_out),
    .data_in(sw_348_data_out),
    .data_out(sw_349_data_out),
    .latch_enable_in(sw_348_latch_out),
    .latch_enable_out(sw_349_latch_out),
    .scan_select_in(sw_348_scan_out),
    .scan_select_out(sw_349_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_349_module_data_in[7] ,
    \sw_349_module_data_in[6] ,
    \sw_349_module_data_in[5] ,
    \sw_349_module_data_in[4] ,
    \sw_349_module_data_in[3] ,
    \sw_349_module_data_in[2] ,
    \sw_349_module_data_in[1] ,
    \sw_349_module_data_in[0] }),
    .module_data_out({\sw_349_module_data_out[7] ,
    \sw_349_module_data_out[6] ,
    \sw_349_module_data_out[5] ,
    \sw_349_module_data_out[4] ,
    \sw_349_module_data_out[3] ,
    \sw_349_module_data_out[2] ,
    \sw_349_module_data_out[1] ,
    \sw_349_module_data_out[0] }));
 scanchain scanchain_35 (.clk_in(sw_034_clk_out),
    .clk_out(sw_035_clk_out),
    .data_in(sw_034_data_out),
    .data_out(sw_035_data_out),
    .latch_enable_in(sw_034_latch_out),
    .latch_enable_out(sw_035_latch_out),
    .scan_select_in(sw_034_scan_out),
    .scan_select_out(sw_035_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_035_module_data_in[7] ,
    \sw_035_module_data_in[6] ,
    \sw_035_module_data_in[5] ,
    \sw_035_module_data_in[4] ,
    \sw_035_module_data_in[3] ,
    \sw_035_module_data_in[2] ,
    \sw_035_module_data_in[1] ,
    \sw_035_module_data_in[0] }),
    .module_data_out({\sw_035_module_data_out[7] ,
    \sw_035_module_data_out[6] ,
    \sw_035_module_data_out[5] ,
    \sw_035_module_data_out[4] ,
    \sw_035_module_data_out[3] ,
    \sw_035_module_data_out[2] ,
    \sw_035_module_data_out[1] ,
    \sw_035_module_data_out[0] }));
 scanchain scanchain_350 (.clk_in(sw_349_clk_out),
    .clk_out(sw_350_clk_out),
    .data_in(sw_349_data_out),
    .data_out(sw_350_data_out),
    .latch_enable_in(sw_349_latch_out),
    .latch_enable_out(sw_350_latch_out),
    .scan_select_in(sw_349_scan_out),
    .scan_select_out(sw_350_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_350_module_data_in[7] ,
    \sw_350_module_data_in[6] ,
    \sw_350_module_data_in[5] ,
    \sw_350_module_data_in[4] ,
    \sw_350_module_data_in[3] ,
    \sw_350_module_data_in[2] ,
    \sw_350_module_data_in[1] ,
    \sw_350_module_data_in[0] }),
    .module_data_out({\sw_350_module_data_out[7] ,
    \sw_350_module_data_out[6] ,
    \sw_350_module_data_out[5] ,
    \sw_350_module_data_out[4] ,
    \sw_350_module_data_out[3] ,
    \sw_350_module_data_out[2] ,
    \sw_350_module_data_out[1] ,
    \sw_350_module_data_out[0] }));
 scanchain scanchain_351 (.clk_in(sw_350_clk_out),
    .clk_out(sw_351_clk_out),
    .data_in(sw_350_data_out),
    .data_out(sw_351_data_out),
    .latch_enable_in(sw_350_latch_out),
    .latch_enable_out(sw_351_latch_out),
    .scan_select_in(sw_350_scan_out),
    .scan_select_out(sw_351_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_351_module_data_in[7] ,
    \sw_351_module_data_in[6] ,
    \sw_351_module_data_in[5] ,
    \sw_351_module_data_in[4] ,
    \sw_351_module_data_in[3] ,
    \sw_351_module_data_in[2] ,
    \sw_351_module_data_in[1] ,
    \sw_351_module_data_in[0] }),
    .module_data_out({\sw_351_module_data_out[7] ,
    \sw_351_module_data_out[6] ,
    \sw_351_module_data_out[5] ,
    \sw_351_module_data_out[4] ,
    \sw_351_module_data_out[3] ,
    \sw_351_module_data_out[2] ,
    \sw_351_module_data_out[1] ,
    \sw_351_module_data_out[0] }));
 scanchain scanchain_352 (.clk_in(sw_351_clk_out),
    .clk_out(sw_352_clk_out),
    .data_in(sw_351_data_out),
    .data_out(sw_352_data_out),
    .latch_enable_in(sw_351_latch_out),
    .latch_enable_out(sw_352_latch_out),
    .scan_select_in(sw_351_scan_out),
    .scan_select_out(sw_352_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_352_module_data_in[7] ,
    \sw_352_module_data_in[6] ,
    \sw_352_module_data_in[5] ,
    \sw_352_module_data_in[4] ,
    \sw_352_module_data_in[3] ,
    \sw_352_module_data_in[2] ,
    \sw_352_module_data_in[1] ,
    \sw_352_module_data_in[0] }),
    .module_data_out({\sw_352_module_data_out[7] ,
    \sw_352_module_data_out[6] ,
    \sw_352_module_data_out[5] ,
    \sw_352_module_data_out[4] ,
    \sw_352_module_data_out[3] ,
    \sw_352_module_data_out[2] ,
    \sw_352_module_data_out[1] ,
    \sw_352_module_data_out[0] }));
 scanchain scanchain_353 (.clk_in(sw_352_clk_out),
    .clk_out(sw_353_clk_out),
    .data_in(sw_352_data_out),
    .data_out(sw_353_data_out),
    .latch_enable_in(sw_352_latch_out),
    .latch_enable_out(sw_353_latch_out),
    .scan_select_in(sw_352_scan_out),
    .scan_select_out(sw_353_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_353_module_data_in[7] ,
    \sw_353_module_data_in[6] ,
    \sw_353_module_data_in[5] ,
    \sw_353_module_data_in[4] ,
    \sw_353_module_data_in[3] ,
    \sw_353_module_data_in[2] ,
    \sw_353_module_data_in[1] ,
    \sw_353_module_data_in[0] }),
    .module_data_out({\sw_353_module_data_out[7] ,
    \sw_353_module_data_out[6] ,
    \sw_353_module_data_out[5] ,
    \sw_353_module_data_out[4] ,
    \sw_353_module_data_out[3] ,
    \sw_353_module_data_out[2] ,
    \sw_353_module_data_out[1] ,
    \sw_353_module_data_out[0] }));
 scanchain scanchain_354 (.clk_in(sw_353_clk_out),
    .clk_out(sw_354_clk_out),
    .data_in(sw_353_data_out),
    .data_out(sw_354_data_out),
    .latch_enable_in(sw_353_latch_out),
    .latch_enable_out(sw_354_latch_out),
    .scan_select_in(sw_353_scan_out),
    .scan_select_out(sw_354_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_354_module_data_in[7] ,
    \sw_354_module_data_in[6] ,
    \sw_354_module_data_in[5] ,
    \sw_354_module_data_in[4] ,
    \sw_354_module_data_in[3] ,
    \sw_354_module_data_in[2] ,
    \sw_354_module_data_in[1] ,
    \sw_354_module_data_in[0] }),
    .module_data_out({\sw_354_module_data_out[7] ,
    \sw_354_module_data_out[6] ,
    \sw_354_module_data_out[5] ,
    \sw_354_module_data_out[4] ,
    \sw_354_module_data_out[3] ,
    \sw_354_module_data_out[2] ,
    \sw_354_module_data_out[1] ,
    \sw_354_module_data_out[0] }));
 scanchain scanchain_355 (.clk_in(sw_354_clk_out),
    .clk_out(sw_355_clk_out),
    .data_in(sw_354_data_out),
    .data_out(sw_355_data_out),
    .latch_enable_in(sw_354_latch_out),
    .latch_enable_out(sw_355_latch_out),
    .scan_select_in(sw_354_scan_out),
    .scan_select_out(sw_355_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_355_module_data_in[7] ,
    \sw_355_module_data_in[6] ,
    \sw_355_module_data_in[5] ,
    \sw_355_module_data_in[4] ,
    \sw_355_module_data_in[3] ,
    \sw_355_module_data_in[2] ,
    \sw_355_module_data_in[1] ,
    \sw_355_module_data_in[0] }),
    .module_data_out({\sw_355_module_data_out[7] ,
    \sw_355_module_data_out[6] ,
    \sw_355_module_data_out[5] ,
    \sw_355_module_data_out[4] ,
    \sw_355_module_data_out[3] ,
    \sw_355_module_data_out[2] ,
    \sw_355_module_data_out[1] ,
    \sw_355_module_data_out[0] }));
 scanchain scanchain_356 (.clk_in(sw_355_clk_out),
    .clk_out(sw_356_clk_out),
    .data_in(sw_355_data_out),
    .data_out(sw_356_data_out),
    .latch_enable_in(sw_355_latch_out),
    .latch_enable_out(sw_356_latch_out),
    .scan_select_in(sw_355_scan_out),
    .scan_select_out(sw_356_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_356_module_data_in[7] ,
    \sw_356_module_data_in[6] ,
    \sw_356_module_data_in[5] ,
    \sw_356_module_data_in[4] ,
    \sw_356_module_data_in[3] ,
    \sw_356_module_data_in[2] ,
    \sw_356_module_data_in[1] ,
    \sw_356_module_data_in[0] }),
    .module_data_out({\sw_356_module_data_out[7] ,
    \sw_356_module_data_out[6] ,
    \sw_356_module_data_out[5] ,
    \sw_356_module_data_out[4] ,
    \sw_356_module_data_out[3] ,
    \sw_356_module_data_out[2] ,
    \sw_356_module_data_out[1] ,
    \sw_356_module_data_out[0] }));
 scanchain scanchain_357 (.clk_in(sw_356_clk_out),
    .clk_out(sw_357_clk_out),
    .data_in(sw_356_data_out),
    .data_out(sw_357_data_out),
    .latch_enable_in(sw_356_latch_out),
    .latch_enable_out(sw_357_latch_out),
    .scan_select_in(sw_356_scan_out),
    .scan_select_out(sw_357_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_357_module_data_in[7] ,
    \sw_357_module_data_in[6] ,
    \sw_357_module_data_in[5] ,
    \sw_357_module_data_in[4] ,
    \sw_357_module_data_in[3] ,
    \sw_357_module_data_in[2] ,
    \sw_357_module_data_in[1] ,
    \sw_357_module_data_in[0] }),
    .module_data_out({\sw_357_module_data_out[7] ,
    \sw_357_module_data_out[6] ,
    \sw_357_module_data_out[5] ,
    \sw_357_module_data_out[4] ,
    \sw_357_module_data_out[3] ,
    \sw_357_module_data_out[2] ,
    \sw_357_module_data_out[1] ,
    \sw_357_module_data_out[0] }));
 scanchain scanchain_358 (.clk_in(sw_357_clk_out),
    .clk_out(sw_358_clk_out),
    .data_in(sw_357_data_out),
    .data_out(sw_358_data_out),
    .latch_enable_in(sw_357_latch_out),
    .latch_enable_out(sw_358_latch_out),
    .scan_select_in(sw_357_scan_out),
    .scan_select_out(sw_358_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_358_module_data_in[7] ,
    \sw_358_module_data_in[6] ,
    \sw_358_module_data_in[5] ,
    \sw_358_module_data_in[4] ,
    \sw_358_module_data_in[3] ,
    \sw_358_module_data_in[2] ,
    \sw_358_module_data_in[1] ,
    \sw_358_module_data_in[0] }),
    .module_data_out({\sw_358_module_data_out[7] ,
    \sw_358_module_data_out[6] ,
    \sw_358_module_data_out[5] ,
    \sw_358_module_data_out[4] ,
    \sw_358_module_data_out[3] ,
    \sw_358_module_data_out[2] ,
    \sw_358_module_data_out[1] ,
    \sw_358_module_data_out[0] }));
 scanchain scanchain_359 (.clk_in(sw_358_clk_out),
    .clk_out(sw_359_clk_out),
    .data_in(sw_358_data_out),
    .data_out(sw_359_data_out),
    .latch_enable_in(sw_358_latch_out),
    .latch_enable_out(sw_359_latch_out),
    .scan_select_in(sw_358_scan_out),
    .scan_select_out(sw_359_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_359_module_data_in[7] ,
    \sw_359_module_data_in[6] ,
    \sw_359_module_data_in[5] ,
    \sw_359_module_data_in[4] ,
    \sw_359_module_data_in[3] ,
    \sw_359_module_data_in[2] ,
    \sw_359_module_data_in[1] ,
    \sw_359_module_data_in[0] }),
    .module_data_out({\sw_359_module_data_out[7] ,
    \sw_359_module_data_out[6] ,
    \sw_359_module_data_out[5] ,
    \sw_359_module_data_out[4] ,
    \sw_359_module_data_out[3] ,
    \sw_359_module_data_out[2] ,
    \sw_359_module_data_out[1] ,
    \sw_359_module_data_out[0] }));
 scanchain scanchain_36 (.clk_in(sw_035_clk_out),
    .clk_out(sw_036_clk_out),
    .data_in(sw_035_data_out),
    .data_out(sw_036_data_out),
    .latch_enable_in(sw_035_latch_out),
    .latch_enable_out(sw_036_latch_out),
    .scan_select_in(sw_035_scan_out),
    .scan_select_out(sw_036_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_036_module_data_in[7] ,
    \sw_036_module_data_in[6] ,
    \sw_036_module_data_in[5] ,
    \sw_036_module_data_in[4] ,
    \sw_036_module_data_in[3] ,
    \sw_036_module_data_in[2] ,
    \sw_036_module_data_in[1] ,
    \sw_036_module_data_in[0] }),
    .module_data_out({\sw_036_module_data_out[7] ,
    \sw_036_module_data_out[6] ,
    \sw_036_module_data_out[5] ,
    \sw_036_module_data_out[4] ,
    \sw_036_module_data_out[3] ,
    \sw_036_module_data_out[2] ,
    \sw_036_module_data_out[1] ,
    \sw_036_module_data_out[0] }));
 scanchain scanchain_360 (.clk_in(sw_359_clk_out),
    .clk_out(sw_360_clk_out),
    .data_in(sw_359_data_out),
    .data_out(sw_360_data_out),
    .latch_enable_in(sw_359_latch_out),
    .latch_enable_out(sw_360_latch_out),
    .scan_select_in(sw_359_scan_out),
    .scan_select_out(sw_360_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_360_module_data_in[7] ,
    \sw_360_module_data_in[6] ,
    \sw_360_module_data_in[5] ,
    \sw_360_module_data_in[4] ,
    \sw_360_module_data_in[3] ,
    \sw_360_module_data_in[2] ,
    \sw_360_module_data_in[1] ,
    \sw_360_module_data_in[0] }),
    .module_data_out({\sw_360_module_data_out[7] ,
    \sw_360_module_data_out[6] ,
    \sw_360_module_data_out[5] ,
    \sw_360_module_data_out[4] ,
    \sw_360_module_data_out[3] ,
    \sw_360_module_data_out[2] ,
    \sw_360_module_data_out[1] ,
    \sw_360_module_data_out[0] }));
 scanchain scanchain_361 (.clk_in(sw_360_clk_out),
    .clk_out(sw_361_clk_out),
    .data_in(sw_360_data_out),
    .data_out(sw_361_data_out),
    .latch_enable_in(sw_360_latch_out),
    .latch_enable_out(sw_361_latch_out),
    .scan_select_in(sw_360_scan_out),
    .scan_select_out(sw_361_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_361_module_data_in[7] ,
    \sw_361_module_data_in[6] ,
    \sw_361_module_data_in[5] ,
    \sw_361_module_data_in[4] ,
    \sw_361_module_data_in[3] ,
    \sw_361_module_data_in[2] ,
    \sw_361_module_data_in[1] ,
    \sw_361_module_data_in[0] }),
    .module_data_out({\sw_361_module_data_out[7] ,
    \sw_361_module_data_out[6] ,
    \sw_361_module_data_out[5] ,
    \sw_361_module_data_out[4] ,
    \sw_361_module_data_out[3] ,
    \sw_361_module_data_out[2] ,
    \sw_361_module_data_out[1] ,
    \sw_361_module_data_out[0] }));
 scanchain scanchain_362 (.clk_in(sw_361_clk_out),
    .clk_out(sw_362_clk_out),
    .data_in(sw_361_data_out),
    .data_out(sw_362_data_out),
    .latch_enable_in(sw_361_latch_out),
    .latch_enable_out(sw_362_latch_out),
    .scan_select_in(sw_361_scan_out),
    .scan_select_out(sw_362_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_362_module_data_in[7] ,
    \sw_362_module_data_in[6] ,
    \sw_362_module_data_in[5] ,
    \sw_362_module_data_in[4] ,
    \sw_362_module_data_in[3] ,
    \sw_362_module_data_in[2] ,
    \sw_362_module_data_in[1] ,
    \sw_362_module_data_in[0] }),
    .module_data_out({\sw_362_module_data_out[7] ,
    \sw_362_module_data_out[6] ,
    \sw_362_module_data_out[5] ,
    \sw_362_module_data_out[4] ,
    \sw_362_module_data_out[3] ,
    \sw_362_module_data_out[2] ,
    \sw_362_module_data_out[1] ,
    \sw_362_module_data_out[0] }));
 scanchain scanchain_363 (.clk_in(sw_362_clk_out),
    .clk_out(sw_363_clk_out),
    .data_in(sw_362_data_out),
    .data_out(sw_363_data_out),
    .latch_enable_in(sw_362_latch_out),
    .latch_enable_out(sw_363_latch_out),
    .scan_select_in(sw_362_scan_out),
    .scan_select_out(sw_363_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_363_module_data_in[7] ,
    \sw_363_module_data_in[6] ,
    \sw_363_module_data_in[5] ,
    \sw_363_module_data_in[4] ,
    \sw_363_module_data_in[3] ,
    \sw_363_module_data_in[2] ,
    \sw_363_module_data_in[1] ,
    \sw_363_module_data_in[0] }),
    .module_data_out({\sw_363_module_data_out[7] ,
    \sw_363_module_data_out[6] ,
    \sw_363_module_data_out[5] ,
    \sw_363_module_data_out[4] ,
    \sw_363_module_data_out[3] ,
    \sw_363_module_data_out[2] ,
    \sw_363_module_data_out[1] ,
    \sw_363_module_data_out[0] }));
 scanchain scanchain_364 (.clk_in(sw_363_clk_out),
    .clk_out(sw_364_clk_out),
    .data_in(sw_363_data_out),
    .data_out(sw_364_data_out),
    .latch_enable_in(sw_363_latch_out),
    .latch_enable_out(sw_364_latch_out),
    .scan_select_in(sw_363_scan_out),
    .scan_select_out(sw_364_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_364_module_data_in[7] ,
    \sw_364_module_data_in[6] ,
    \sw_364_module_data_in[5] ,
    \sw_364_module_data_in[4] ,
    \sw_364_module_data_in[3] ,
    \sw_364_module_data_in[2] ,
    \sw_364_module_data_in[1] ,
    \sw_364_module_data_in[0] }),
    .module_data_out({\sw_364_module_data_out[7] ,
    \sw_364_module_data_out[6] ,
    \sw_364_module_data_out[5] ,
    \sw_364_module_data_out[4] ,
    \sw_364_module_data_out[3] ,
    \sw_364_module_data_out[2] ,
    \sw_364_module_data_out[1] ,
    \sw_364_module_data_out[0] }));
 scanchain scanchain_365 (.clk_in(sw_364_clk_out),
    .clk_out(sw_365_clk_out),
    .data_in(sw_364_data_out),
    .data_out(sw_365_data_out),
    .latch_enable_in(sw_364_latch_out),
    .latch_enable_out(sw_365_latch_out),
    .scan_select_in(sw_364_scan_out),
    .scan_select_out(sw_365_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_365_module_data_in[7] ,
    \sw_365_module_data_in[6] ,
    \sw_365_module_data_in[5] ,
    \sw_365_module_data_in[4] ,
    \sw_365_module_data_in[3] ,
    \sw_365_module_data_in[2] ,
    \sw_365_module_data_in[1] ,
    \sw_365_module_data_in[0] }),
    .module_data_out({\sw_365_module_data_out[7] ,
    \sw_365_module_data_out[6] ,
    \sw_365_module_data_out[5] ,
    \sw_365_module_data_out[4] ,
    \sw_365_module_data_out[3] ,
    \sw_365_module_data_out[2] ,
    \sw_365_module_data_out[1] ,
    \sw_365_module_data_out[0] }));
 scanchain scanchain_366 (.clk_in(sw_365_clk_out),
    .clk_out(sw_366_clk_out),
    .data_in(sw_365_data_out),
    .data_out(sw_366_data_out),
    .latch_enable_in(sw_365_latch_out),
    .latch_enable_out(sw_366_latch_out),
    .scan_select_in(sw_365_scan_out),
    .scan_select_out(sw_366_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_366_module_data_in[7] ,
    \sw_366_module_data_in[6] ,
    \sw_366_module_data_in[5] ,
    \sw_366_module_data_in[4] ,
    \sw_366_module_data_in[3] ,
    \sw_366_module_data_in[2] ,
    \sw_366_module_data_in[1] ,
    \sw_366_module_data_in[0] }),
    .module_data_out({\sw_366_module_data_out[7] ,
    \sw_366_module_data_out[6] ,
    \sw_366_module_data_out[5] ,
    \sw_366_module_data_out[4] ,
    \sw_366_module_data_out[3] ,
    \sw_366_module_data_out[2] ,
    \sw_366_module_data_out[1] ,
    \sw_366_module_data_out[0] }));
 scanchain scanchain_367 (.clk_in(sw_366_clk_out),
    .clk_out(sw_367_clk_out),
    .data_in(sw_366_data_out),
    .data_out(sw_367_data_out),
    .latch_enable_in(sw_366_latch_out),
    .latch_enable_out(sw_367_latch_out),
    .scan_select_in(sw_366_scan_out),
    .scan_select_out(sw_367_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_367_module_data_in[7] ,
    \sw_367_module_data_in[6] ,
    \sw_367_module_data_in[5] ,
    \sw_367_module_data_in[4] ,
    \sw_367_module_data_in[3] ,
    \sw_367_module_data_in[2] ,
    \sw_367_module_data_in[1] ,
    \sw_367_module_data_in[0] }),
    .module_data_out({\sw_367_module_data_out[7] ,
    \sw_367_module_data_out[6] ,
    \sw_367_module_data_out[5] ,
    \sw_367_module_data_out[4] ,
    \sw_367_module_data_out[3] ,
    \sw_367_module_data_out[2] ,
    \sw_367_module_data_out[1] ,
    \sw_367_module_data_out[0] }));
 scanchain scanchain_368 (.clk_in(sw_367_clk_out),
    .clk_out(sw_368_clk_out),
    .data_in(sw_367_data_out),
    .data_out(sw_368_data_out),
    .latch_enable_in(sw_367_latch_out),
    .latch_enable_out(sw_368_latch_out),
    .scan_select_in(sw_367_scan_out),
    .scan_select_out(sw_368_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_368_module_data_in[7] ,
    \sw_368_module_data_in[6] ,
    \sw_368_module_data_in[5] ,
    \sw_368_module_data_in[4] ,
    \sw_368_module_data_in[3] ,
    \sw_368_module_data_in[2] ,
    \sw_368_module_data_in[1] ,
    \sw_368_module_data_in[0] }),
    .module_data_out({\sw_368_module_data_out[7] ,
    \sw_368_module_data_out[6] ,
    \sw_368_module_data_out[5] ,
    \sw_368_module_data_out[4] ,
    \sw_368_module_data_out[3] ,
    \sw_368_module_data_out[2] ,
    \sw_368_module_data_out[1] ,
    \sw_368_module_data_out[0] }));
 scanchain scanchain_369 (.clk_in(sw_368_clk_out),
    .clk_out(sw_369_clk_out),
    .data_in(sw_368_data_out),
    .data_out(sw_369_data_out),
    .latch_enable_in(sw_368_latch_out),
    .latch_enable_out(sw_369_latch_out),
    .scan_select_in(sw_368_scan_out),
    .scan_select_out(sw_369_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_369_module_data_in[7] ,
    \sw_369_module_data_in[6] ,
    \sw_369_module_data_in[5] ,
    \sw_369_module_data_in[4] ,
    \sw_369_module_data_in[3] ,
    \sw_369_module_data_in[2] ,
    \sw_369_module_data_in[1] ,
    \sw_369_module_data_in[0] }),
    .module_data_out({\sw_369_module_data_out[7] ,
    \sw_369_module_data_out[6] ,
    \sw_369_module_data_out[5] ,
    \sw_369_module_data_out[4] ,
    \sw_369_module_data_out[3] ,
    \sw_369_module_data_out[2] ,
    \sw_369_module_data_out[1] ,
    \sw_369_module_data_out[0] }));
 scanchain scanchain_37 (.clk_in(sw_036_clk_out),
    .clk_out(sw_037_clk_out),
    .data_in(sw_036_data_out),
    .data_out(sw_037_data_out),
    .latch_enable_in(sw_036_latch_out),
    .latch_enable_out(sw_037_latch_out),
    .scan_select_in(sw_036_scan_out),
    .scan_select_out(sw_037_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_037_module_data_in[7] ,
    \sw_037_module_data_in[6] ,
    \sw_037_module_data_in[5] ,
    \sw_037_module_data_in[4] ,
    \sw_037_module_data_in[3] ,
    \sw_037_module_data_in[2] ,
    \sw_037_module_data_in[1] ,
    \sw_037_module_data_in[0] }),
    .module_data_out({\sw_037_module_data_out[7] ,
    \sw_037_module_data_out[6] ,
    \sw_037_module_data_out[5] ,
    \sw_037_module_data_out[4] ,
    \sw_037_module_data_out[3] ,
    \sw_037_module_data_out[2] ,
    \sw_037_module_data_out[1] ,
    \sw_037_module_data_out[0] }));
 scanchain scanchain_370 (.clk_in(sw_369_clk_out),
    .clk_out(sw_370_clk_out),
    .data_in(sw_369_data_out),
    .data_out(sw_370_data_out),
    .latch_enable_in(sw_369_latch_out),
    .latch_enable_out(sw_370_latch_out),
    .scan_select_in(sw_369_scan_out),
    .scan_select_out(sw_370_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_370_module_data_in[7] ,
    \sw_370_module_data_in[6] ,
    \sw_370_module_data_in[5] ,
    \sw_370_module_data_in[4] ,
    \sw_370_module_data_in[3] ,
    \sw_370_module_data_in[2] ,
    \sw_370_module_data_in[1] ,
    \sw_370_module_data_in[0] }),
    .module_data_out({\sw_370_module_data_out[7] ,
    \sw_370_module_data_out[6] ,
    \sw_370_module_data_out[5] ,
    \sw_370_module_data_out[4] ,
    \sw_370_module_data_out[3] ,
    \sw_370_module_data_out[2] ,
    \sw_370_module_data_out[1] ,
    \sw_370_module_data_out[0] }));
 scanchain scanchain_371 (.clk_in(sw_370_clk_out),
    .clk_out(sw_371_clk_out),
    .data_in(sw_370_data_out),
    .data_out(sw_371_data_out),
    .latch_enable_in(sw_370_latch_out),
    .latch_enable_out(sw_371_latch_out),
    .scan_select_in(sw_370_scan_out),
    .scan_select_out(sw_371_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_371_module_data_in[7] ,
    \sw_371_module_data_in[6] ,
    \sw_371_module_data_in[5] ,
    \sw_371_module_data_in[4] ,
    \sw_371_module_data_in[3] ,
    \sw_371_module_data_in[2] ,
    \sw_371_module_data_in[1] ,
    \sw_371_module_data_in[0] }),
    .module_data_out({\sw_371_module_data_out[7] ,
    \sw_371_module_data_out[6] ,
    \sw_371_module_data_out[5] ,
    \sw_371_module_data_out[4] ,
    \sw_371_module_data_out[3] ,
    \sw_371_module_data_out[2] ,
    \sw_371_module_data_out[1] ,
    \sw_371_module_data_out[0] }));
 scanchain scanchain_372 (.clk_in(sw_371_clk_out),
    .clk_out(sw_372_clk_out),
    .data_in(sw_371_data_out),
    .data_out(sw_372_data_out),
    .latch_enable_in(sw_371_latch_out),
    .latch_enable_out(sw_372_latch_out),
    .scan_select_in(sw_371_scan_out),
    .scan_select_out(sw_372_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_372_module_data_in[7] ,
    \sw_372_module_data_in[6] ,
    \sw_372_module_data_in[5] ,
    \sw_372_module_data_in[4] ,
    \sw_372_module_data_in[3] ,
    \sw_372_module_data_in[2] ,
    \sw_372_module_data_in[1] ,
    \sw_372_module_data_in[0] }),
    .module_data_out({\sw_372_module_data_out[7] ,
    \sw_372_module_data_out[6] ,
    \sw_372_module_data_out[5] ,
    \sw_372_module_data_out[4] ,
    \sw_372_module_data_out[3] ,
    \sw_372_module_data_out[2] ,
    \sw_372_module_data_out[1] ,
    \sw_372_module_data_out[0] }));
 scanchain scanchain_373 (.clk_in(sw_372_clk_out),
    .clk_out(sw_373_clk_out),
    .data_in(sw_372_data_out),
    .data_out(sw_373_data_out),
    .latch_enable_in(sw_372_latch_out),
    .latch_enable_out(sw_373_latch_out),
    .scan_select_in(sw_372_scan_out),
    .scan_select_out(sw_373_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_373_module_data_in[7] ,
    \sw_373_module_data_in[6] ,
    \sw_373_module_data_in[5] ,
    \sw_373_module_data_in[4] ,
    \sw_373_module_data_in[3] ,
    \sw_373_module_data_in[2] ,
    \sw_373_module_data_in[1] ,
    \sw_373_module_data_in[0] }),
    .module_data_out({\sw_373_module_data_out[7] ,
    \sw_373_module_data_out[6] ,
    \sw_373_module_data_out[5] ,
    \sw_373_module_data_out[4] ,
    \sw_373_module_data_out[3] ,
    \sw_373_module_data_out[2] ,
    \sw_373_module_data_out[1] ,
    \sw_373_module_data_out[0] }));
 scanchain scanchain_374 (.clk_in(sw_373_clk_out),
    .clk_out(sw_374_clk_out),
    .data_in(sw_373_data_out),
    .data_out(sw_374_data_out),
    .latch_enable_in(sw_373_latch_out),
    .latch_enable_out(sw_374_latch_out),
    .scan_select_in(sw_373_scan_out),
    .scan_select_out(sw_374_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_374_module_data_in[7] ,
    \sw_374_module_data_in[6] ,
    \sw_374_module_data_in[5] ,
    \sw_374_module_data_in[4] ,
    \sw_374_module_data_in[3] ,
    \sw_374_module_data_in[2] ,
    \sw_374_module_data_in[1] ,
    \sw_374_module_data_in[0] }),
    .module_data_out({\sw_374_module_data_out[7] ,
    \sw_374_module_data_out[6] ,
    \sw_374_module_data_out[5] ,
    \sw_374_module_data_out[4] ,
    \sw_374_module_data_out[3] ,
    \sw_374_module_data_out[2] ,
    \sw_374_module_data_out[1] ,
    \sw_374_module_data_out[0] }));
 scanchain scanchain_375 (.clk_in(sw_374_clk_out),
    .clk_out(sw_375_clk_out),
    .data_in(sw_374_data_out),
    .data_out(sw_375_data_out),
    .latch_enable_in(sw_374_latch_out),
    .latch_enable_out(sw_375_latch_out),
    .scan_select_in(sw_374_scan_out),
    .scan_select_out(sw_375_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_375_module_data_in[7] ,
    \sw_375_module_data_in[6] ,
    \sw_375_module_data_in[5] ,
    \sw_375_module_data_in[4] ,
    \sw_375_module_data_in[3] ,
    \sw_375_module_data_in[2] ,
    \sw_375_module_data_in[1] ,
    \sw_375_module_data_in[0] }),
    .module_data_out({\sw_375_module_data_out[7] ,
    \sw_375_module_data_out[6] ,
    \sw_375_module_data_out[5] ,
    \sw_375_module_data_out[4] ,
    \sw_375_module_data_out[3] ,
    \sw_375_module_data_out[2] ,
    \sw_375_module_data_out[1] ,
    \sw_375_module_data_out[0] }));
 scanchain scanchain_376 (.clk_in(sw_375_clk_out),
    .clk_out(sw_376_clk_out),
    .data_in(sw_375_data_out),
    .data_out(sw_376_data_out),
    .latch_enable_in(sw_375_latch_out),
    .latch_enable_out(sw_376_latch_out),
    .scan_select_in(sw_375_scan_out),
    .scan_select_out(sw_376_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_376_module_data_in[7] ,
    \sw_376_module_data_in[6] ,
    \sw_376_module_data_in[5] ,
    \sw_376_module_data_in[4] ,
    \sw_376_module_data_in[3] ,
    \sw_376_module_data_in[2] ,
    \sw_376_module_data_in[1] ,
    \sw_376_module_data_in[0] }),
    .module_data_out({\sw_376_module_data_out[7] ,
    \sw_376_module_data_out[6] ,
    \sw_376_module_data_out[5] ,
    \sw_376_module_data_out[4] ,
    \sw_376_module_data_out[3] ,
    \sw_376_module_data_out[2] ,
    \sw_376_module_data_out[1] ,
    \sw_376_module_data_out[0] }));
 scanchain scanchain_377 (.clk_in(sw_376_clk_out),
    .clk_out(sw_377_clk_out),
    .data_in(sw_376_data_out),
    .data_out(sw_377_data_out),
    .latch_enable_in(sw_376_latch_out),
    .latch_enable_out(sw_377_latch_out),
    .scan_select_in(sw_376_scan_out),
    .scan_select_out(sw_377_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_377_module_data_in[7] ,
    \sw_377_module_data_in[6] ,
    \sw_377_module_data_in[5] ,
    \sw_377_module_data_in[4] ,
    \sw_377_module_data_in[3] ,
    \sw_377_module_data_in[2] ,
    \sw_377_module_data_in[1] ,
    \sw_377_module_data_in[0] }),
    .module_data_out({\sw_377_module_data_out[7] ,
    \sw_377_module_data_out[6] ,
    \sw_377_module_data_out[5] ,
    \sw_377_module_data_out[4] ,
    \sw_377_module_data_out[3] ,
    \sw_377_module_data_out[2] ,
    \sw_377_module_data_out[1] ,
    \sw_377_module_data_out[0] }));
 scanchain scanchain_378 (.clk_in(sw_377_clk_out),
    .clk_out(sw_378_clk_out),
    .data_in(sw_377_data_out),
    .data_out(sw_378_data_out),
    .latch_enable_in(sw_377_latch_out),
    .latch_enable_out(sw_378_latch_out),
    .scan_select_in(sw_377_scan_out),
    .scan_select_out(sw_378_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_378_module_data_in[7] ,
    \sw_378_module_data_in[6] ,
    \sw_378_module_data_in[5] ,
    \sw_378_module_data_in[4] ,
    \sw_378_module_data_in[3] ,
    \sw_378_module_data_in[2] ,
    \sw_378_module_data_in[1] ,
    \sw_378_module_data_in[0] }),
    .module_data_out({\sw_378_module_data_out[7] ,
    \sw_378_module_data_out[6] ,
    \sw_378_module_data_out[5] ,
    \sw_378_module_data_out[4] ,
    \sw_378_module_data_out[3] ,
    \sw_378_module_data_out[2] ,
    \sw_378_module_data_out[1] ,
    \sw_378_module_data_out[0] }));
 scanchain scanchain_379 (.clk_in(sw_378_clk_out),
    .clk_out(sw_379_clk_out),
    .data_in(sw_378_data_out),
    .data_out(sw_379_data_out),
    .latch_enable_in(sw_378_latch_out),
    .latch_enable_out(sw_379_latch_out),
    .scan_select_in(sw_378_scan_out),
    .scan_select_out(sw_379_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_379_module_data_in[7] ,
    \sw_379_module_data_in[6] ,
    \sw_379_module_data_in[5] ,
    \sw_379_module_data_in[4] ,
    \sw_379_module_data_in[3] ,
    \sw_379_module_data_in[2] ,
    \sw_379_module_data_in[1] ,
    \sw_379_module_data_in[0] }),
    .module_data_out({\sw_379_module_data_out[7] ,
    \sw_379_module_data_out[6] ,
    \sw_379_module_data_out[5] ,
    \sw_379_module_data_out[4] ,
    \sw_379_module_data_out[3] ,
    \sw_379_module_data_out[2] ,
    \sw_379_module_data_out[1] ,
    \sw_379_module_data_out[0] }));
 scanchain scanchain_38 (.clk_in(sw_037_clk_out),
    .clk_out(sw_038_clk_out),
    .data_in(sw_037_data_out),
    .data_out(sw_038_data_out),
    .latch_enable_in(sw_037_latch_out),
    .latch_enable_out(sw_038_latch_out),
    .scan_select_in(sw_037_scan_out),
    .scan_select_out(sw_038_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_038_module_data_in[7] ,
    \sw_038_module_data_in[6] ,
    \sw_038_module_data_in[5] ,
    \sw_038_module_data_in[4] ,
    \sw_038_module_data_in[3] ,
    \sw_038_module_data_in[2] ,
    \sw_038_module_data_in[1] ,
    \sw_038_module_data_in[0] }),
    .module_data_out({\sw_038_module_data_out[7] ,
    \sw_038_module_data_out[6] ,
    \sw_038_module_data_out[5] ,
    \sw_038_module_data_out[4] ,
    \sw_038_module_data_out[3] ,
    \sw_038_module_data_out[2] ,
    \sw_038_module_data_out[1] ,
    \sw_038_module_data_out[0] }));
 scanchain scanchain_380 (.clk_in(sw_379_clk_out),
    .clk_out(sw_380_clk_out),
    .data_in(sw_379_data_out),
    .data_out(sw_380_data_out),
    .latch_enable_in(sw_379_latch_out),
    .latch_enable_out(sw_380_latch_out),
    .scan_select_in(sw_379_scan_out),
    .scan_select_out(sw_380_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_380_module_data_in[7] ,
    \sw_380_module_data_in[6] ,
    \sw_380_module_data_in[5] ,
    \sw_380_module_data_in[4] ,
    \sw_380_module_data_in[3] ,
    \sw_380_module_data_in[2] ,
    \sw_380_module_data_in[1] ,
    \sw_380_module_data_in[0] }),
    .module_data_out({\sw_380_module_data_out[7] ,
    \sw_380_module_data_out[6] ,
    \sw_380_module_data_out[5] ,
    \sw_380_module_data_out[4] ,
    \sw_380_module_data_out[3] ,
    \sw_380_module_data_out[2] ,
    \sw_380_module_data_out[1] ,
    \sw_380_module_data_out[0] }));
 scanchain scanchain_381 (.clk_in(sw_380_clk_out),
    .clk_out(sw_381_clk_out),
    .data_in(sw_380_data_out),
    .data_out(sw_381_data_out),
    .latch_enable_in(sw_380_latch_out),
    .latch_enable_out(sw_381_latch_out),
    .scan_select_in(sw_380_scan_out),
    .scan_select_out(sw_381_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_381_module_data_in[7] ,
    \sw_381_module_data_in[6] ,
    \sw_381_module_data_in[5] ,
    \sw_381_module_data_in[4] ,
    \sw_381_module_data_in[3] ,
    \sw_381_module_data_in[2] ,
    \sw_381_module_data_in[1] ,
    \sw_381_module_data_in[0] }),
    .module_data_out({\sw_381_module_data_out[7] ,
    \sw_381_module_data_out[6] ,
    \sw_381_module_data_out[5] ,
    \sw_381_module_data_out[4] ,
    \sw_381_module_data_out[3] ,
    \sw_381_module_data_out[2] ,
    \sw_381_module_data_out[1] ,
    \sw_381_module_data_out[0] }));
 scanchain scanchain_382 (.clk_in(sw_381_clk_out),
    .clk_out(sw_382_clk_out),
    .data_in(sw_381_data_out),
    .data_out(sw_382_data_out),
    .latch_enable_in(sw_381_latch_out),
    .latch_enable_out(sw_382_latch_out),
    .scan_select_in(sw_381_scan_out),
    .scan_select_out(sw_382_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_382_module_data_in[7] ,
    \sw_382_module_data_in[6] ,
    \sw_382_module_data_in[5] ,
    \sw_382_module_data_in[4] ,
    \sw_382_module_data_in[3] ,
    \sw_382_module_data_in[2] ,
    \sw_382_module_data_in[1] ,
    \sw_382_module_data_in[0] }),
    .module_data_out({\sw_382_module_data_out[7] ,
    \sw_382_module_data_out[6] ,
    \sw_382_module_data_out[5] ,
    \sw_382_module_data_out[4] ,
    \sw_382_module_data_out[3] ,
    \sw_382_module_data_out[2] ,
    \sw_382_module_data_out[1] ,
    \sw_382_module_data_out[0] }));
 scanchain scanchain_383 (.clk_in(sw_382_clk_out),
    .clk_out(sw_383_clk_out),
    .data_in(sw_382_data_out),
    .data_out(sw_383_data_out),
    .latch_enable_in(sw_382_latch_out),
    .latch_enable_out(sw_383_latch_out),
    .scan_select_in(sw_382_scan_out),
    .scan_select_out(sw_383_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_383_module_data_in[7] ,
    \sw_383_module_data_in[6] ,
    \sw_383_module_data_in[5] ,
    \sw_383_module_data_in[4] ,
    \sw_383_module_data_in[3] ,
    \sw_383_module_data_in[2] ,
    \sw_383_module_data_in[1] ,
    \sw_383_module_data_in[0] }),
    .module_data_out({\sw_383_module_data_out[7] ,
    \sw_383_module_data_out[6] ,
    \sw_383_module_data_out[5] ,
    \sw_383_module_data_out[4] ,
    \sw_383_module_data_out[3] ,
    \sw_383_module_data_out[2] ,
    \sw_383_module_data_out[1] ,
    \sw_383_module_data_out[0] }));
 scanchain scanchain_384 (.clk_in(sw_383_clk_out),
    .clk_out(sw_384_clk_out),
    .data_in(sw_383_data_out),
    .data_out(sw_384_data_out),
    .latch_enable_in(sw_383_latch_out),
    .latch_enable_out(sw_384_latch_out),
    .scan_select_in(sw_383_scan_out),
    .scan_select_out(sw_384_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_384_module_data_in[7] ,
    \sw_384_module_data_in[6] ,
    \sw_384_module_data_in[5] ,
    \sw_384_module_data_in[4] ,
    \sw_384_module_data_in[3] ,
    \sw_384_module_data_in[2] ,
    \sw_384_module_data_in[1] ,
    \sw_384_module_data_in[0] }),
    .module_data_out({\sw_384_module_data_out[7] ,
    \sw_384_module_data_out[6] ,
    \sw_384_module_data_out[5] ,
    \sw_384_module_data_out[4] ,
    \sw_384_module_data_out[3] ,
    \sw_384_module_data_out[2] ,
    \sw_384_module_data_out[1] ,
    \sw_384_module_data_out[0] }));
 scanchain scanchain_385 (.clk_in(sw_384_clk_out),
    .clk_out(sw_385_clk_out),
    .data_in(sw_384_data_out),
    .data_out(sw_385_data_out),
    .latch_enable_in(sw_384_latch_out),
    .latch_enable_out(sw_385_latch_out),
    .scan_select_in(sw_384_scan_out),
    .scan_select_out(sw_385_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_385_module_data_in[7] ,
    \sw_385_module_data_in[6] ,
    \sw_385_module_data_in[5] ,
    \sw_385_module_data_in[4] ,
    \sw_385_module_data_in[3] ,
    \sw_385_module_data_in[2] ,
    \sw_385_module_data_in[1] ,
    \sw_385_module_data_in[0] }),
    .module_data_out({\sw_385_module_data_out[7] ,
    \sw_385_module_data_out[6] ,
    \sw_385_module_data_out[5] ,
    \sw_385_module_data_out[4] ,
    \sw_385_module_data_out[3] ,
    \sw_385_module_data_out[2] ,
    \sw_385_module_data_out[1] ,
    \sw_385_module_data_out[0] }));
 scanchain scanchain_386 (.clk_in(sw_385_clk_out),
    .clk_out(sw_386_clk_out),
    .data_in(sw_385_data_out),
    .data_out(sw_386_data_out),
    .latch_enable_in(sw_385_latch_out),
    .latch_enable_out(sw_386_latch_out),
    .scan_select_in(sw_385_scan_out),
    .scan_select_out(sw_386_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_386_module_data_in[7] ,
    \sw_386_module_data_in[6] ,
    \sw_386_module_data_in[5] ,
    \sw_386_module_data_in[4] ,
    \sw_386_module_data_in[3] ,
    \sw_386_module_data_in[2] ,
    \sw_386_module_data_in[1] ,
    \sw_386_module_data_in[0] }),
    .module_data_out({\sw_386_module_data_out[7] ,
    \sw_386_module_data_out[6] ,
    \sw_386_module_data_out[5] ,
    \sw_386_module_data_out[4] ,
    \sw_386_module_data_out[3] ,
    \sw_386_module_data_out[2] ,
    \sw_386_module_data_out[1] ,
    \sw_386_module_data_out[0] }));
 scanchain scanchain_387 (.clk_in(sw_386_clk_out),
    .clk_out(sw_387_clk_out),
    .data_in(sw_386_data_out),
    .data_out(sw_387_data_out),
    .latch_enable_in(sw_386_latch_out),
    .latch_enable_out(sw_387_latch_out),
    .scan_select_in(sw_386_scan_out),
    .scan_select_out(sw_387_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_387_module_data_in[7] ,
    \sw_387_module_data_in[6] ,
    \sw_387_module_data_in[5] ,
    \sw_387_module_data_in[4] ,
    \sw_387_module_data_in[3] ,
    \sw_387_module_data_in[2] ,
    \sw_387_module_data_in[1] ,
    \sw_387_module_data_in[0] }),
    .module_data_out({\sw_387_module_data_out[7] ,
    \sw_387_module_data_out[6] ,
    \sw_387_module_data_out[5] ,
    \sw_387_module_data_out[4] ,
    \sw_387_module_data_out[3] ,
    \sw_387_module_data_out[2] ,
    \sw_387_module_data_out[1] ,
    \sw_387_module_data_out[0] }));
 scanchain scanchain_388 (.clk_in(sw_387_clk_out),
    .clk_out(sw_388_clk_out),
    .data_in(sw_387_data_out),
    .data_out(sw_388_data_out),
    .latch_enable_in(sw_387_latch_out),
    .latch_enable_out(sw_388_latch_out),
    .scan_select_in(sw_387_scan_out),
    .scan_select_out(sw_388_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_388_module_data_in[7] ,
    \sw_388_module_data_in[6] ,
    \sw_388_module_data_in[5] ,
    \sw_388_module_data_in[4] ,
    \sw_388_module_data_in[3] ,
    \sw_388_module_data_in[2] ,
    \sw_388_module_data_in[1] ,
    \sw_388_module_data_in[0] }),
    .module_data_out({\sw_388_module_data_out[7] ,
    \sw_388_module_data_out[6] ,
    \sw_388_module_data_out[5] ,
    \sw_388_module_data_out[4] ,
    \sw_388_module_data_out[3] ,
    \sw_388_module_data_out[2] ,
    \sw_388_module_data_out[1] ,
    \sw_388_module_data_out[0] }));
 scanchain scanchain_389 (.clk_in(sw_388_clk_out),
    .clk_out(sw_389_clk_out),
    .data_in(sw_388_data_out),
    .data_out(sw_389_data_out),
    .latch_enable_in(sw_388_latch_out),
    .latch_enable_out(sw_389_latch_out),
    .scan_select_in(sw_388_scan_out),
    .scan_select_out(sw_389_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_389_module_data_in[7] ,
    \sw_389_module_data_in[6] ,
    \sw_389_module_data_in[5] ,
    \sw_389_module_data_in[4] ,
    \sw_389_module_data_in[3] ,
    \sw_389_module_data_in[2] ,
    \sw_389_module_data_in[1] ,
    \sw_389_module_data_in[0] }),
    .module_data_out({\sw_389_module_data_out[7] ,
    \sw_389_module_data_out[6] ,
    \sw_389_module_data_out[5] ,
    \sw_389_module_data_out[4] ,
    \sw_389_module_data_out[3] ,
    \sw_389_module_data_out[2] ,
    \sw_389_module_data_out[1] ,
    \sw_389_module_data_out[0] }));
 scanchain scanchain_39 (.clk_in(sw_038_clk_out),
    .clk_out(sw_039_clk_out),
    .data_in(sw_038_data_out),
    .data_out(sw_039_data_out),
    .latch_enable_in(sw_038_latch_out),
    .latch_enable_out(sw_039_latch_out),
    .scan_select_in(sw_038_scan_out),
    .scan_select_out(sw_039_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_039_module_data_in[7] ,
    \sw_039_module_data_in[6] ,
    \sw_039_module_data_in[5] ,
    \sw_039_module_data_in[4] ,
    \sw_039_module_data_in[3] ,
    \sw_039_module_data_in[2] ,
    \sw_039_module_data_in[1] ,
    \sw_039_module_data_in[0] }),
    .module_data_out({\sw_039_module_data_out[7] ,
    \sw_039_module_data_out[6] ,
    \sw_039_module_data_out[5] ,
    \sw_039_module_data_out[4] ,
    \sw_039_module_data_out[3] ,
    \sw_039_module_data_out[2] ,
    \sw_039_module_data_out[1] ,
    \sw_039_module_data_out[0] }));
 scanchain scanchain_390 (.clk_in(sw_389_clk_out),
    .clk_out(sw_390_clk_out),
    .data_in(sw_389_data_out),
    .data_out(sw_390_data_out),
    .latch_enable_in(sw_389_latch_out),
    .latch_enable_out(sw_390_latch_out),
    .scan_select_in(sw_389_scan_out),
    .scan_select_out(sw_390_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_390_module_data_in[7] ,
    \sw_390_module_data_in[6] ,
    \sw_390_module_data_in[5] ,
    \sw_390_module_data_in[4] ,
    \sw_390_module_data_in[3] ,
    \sw_390_module_data_in[2] ,
    \sw_390_module_data_in[1] ,
    \sw_390_module_data_in[0] }),
    .module_data_out({\sw_390_module_data_out[7] ,
    \sw_390_module_data_out[6] ,
    \sw_390_module_data_out[5] ,
    \sw_390_module_data_out[4] ,
    \sw_390_module_data_out[3] ,
    \sw_390_module_data_out[2] ,
    \sw_390_module_data_out[1] ,
    \sw_390_module_data_out[0] }));
 scanchain scanchain_391 (.clk_in(sw_390_clk_out),
    .clk_out(sw_391_clk_out),
    .data_in(sw_390_data_out),
    .data_out(sw_391_data_out),
    .latch_enable_in(sw_390_latch_out),
    .latch_enable_out(sw_391_latch_out),
    .scan_select_in(sw_390_scan_out),
    .scan_select_out(sw_391_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_391_module_data_in[7] ,
    \sw_391_module_data_in[6] ,
    \sw_391_module_data_in[5] ,
    \sw_391_module_data_in[4] ,
    \sw_391_module_data_in[3] ,
    \sw_391_module_data_in[2] ,
    \sw_391_module_data_in[1] ,
    \sw_391_module_data_in[0] }),
    .module_data_out({\sw_391_module_data_out[7] ,
    \sw_391_module_data_out[6] ,
    \sw_391_module_data_out[5] ,
    \sw_391_module_data_out[4] ,
    \sw_391_module_data_out[3] ,
    \sw_391_module_data_out[2] ,
    \sw_391_module_data_out[1] ,
    \sw_391_module_data_out[0] }));
 scanchain scanchain_392 (.clk_in(sw_391_clk_out),
    .clk_out(sw_392_clk_out),
    .data_in(sw_391_data_out),
    .data_out(sw_392_data_out),
    .latch_enable_in(sw_391_latch_out),
    .latch_enable_out(sw_392_latch_out),
    .scan_select_in(sw_391_scan_out),
    .scan_select_out(sw_392_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_392_module_data_in[7] ,
    \sw_392_module_data_in[6] ,
    \sw_392_module_data_in[5] ,
    \sw_392_module_data_in[4] ,
    \sw_392_module_data_in[3] ,
    \sw_392_module_data_in[2] ,
    \sw_392_module_data_in[1] ,
    \sw_392_module_data_in[0] }),
    .module_data_out({\sw_392_module_data_out[7] ,
    \sw_392_module_data_out[6] ,
    \sw_392_module_data_out[5] ,
    \sw_392_module_data_out[4] ,
    \sw_392_module_data_out[3] ,
    \sw_392_module_data_out[2] ,
    \sw_392_module_data_out[1] ,
    \sw_392_module_data_out[0] }));
 scanchain scanchain_393 (.clk_in(sw_392_clk_out),
    .clk_out(sw_393_clk_out),
    .data_in(sw_392_data_out),
    .data_out(sw_393_data_out),
    .latch_enable_in(sw_392_latch_out),
    .latch_enable_out(sw_393_latch_out),
    .scan_select_in(sw_392_scan_out),
    .scan_select_out(sw_393_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_393_module_data_in[7] ,
    \sw_393_module_data_in[6] ,
    \sw_393_module_data_in[5] ,
    \sw_393_module_data_in[4] ,
    \sw_393_module_data_in[3] ,
    \sw_393_module_data_in[2] ,
    \sw_393_module_data_in[1] ,
    \sw_393_module_data_in[0] }),
    .module_data_out({\sw_393_module_data_out[7] ,
    \sw_393_module_data_out[6] ,
    \sw_393_module_data_out[5] ,
    \sw_393_module_data_out[4] ,
    \sw_393_module_data_out[3] ,
    \sw_393_module_data_out[2] ,
    \sw_393_module_data_out[1] ,
    \sw_393_module_data_out[0] }));
 scanchain scanchain_394 (.clk_in(sw_393_clk_out),
    .clk_out(sw_394_clk_out),
    .data_in(sw_393_data_out),
    .data_out(sw_394_data_out),
    .latch_enable_in(sw_393_latch_out),
    .latch_enable_out(sw_394_latch_out),
    .scan_select_in(sw_393_scan_out),
    .scan_select_out(sw_394_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_394_module_data_in[7] ,
    \sw_394_module_data_in[6] ,
    \sw_394_module_data_in[5] ,
    \sw_394_module_data_in[4] ,
    \sw_394_module_data_in[3] ,
    \sw_394_module_data_in[2] ,
    \sw_394_module_data_in[1] ,
    \sw_394_module_data_in[0] }),
    .module_data_out({\sw_394_module_data_out[7] ,
    \sw_394_module_data_out[6] ,
    \sw_394_module_data_out[5] ,
    \sw_394_module_data_out[4] ,
    \sw_394_module_data_out[3] ,
    \sw_394_module_data_out[2] ,
    \sw_394_module_data_out[1] ,
    \sw_394_module_data_out[0] }));
 scanchain scanchain_395 (.clk_in(sw_394_clk_out),
    .clk_out(sw_395_clk_out),
    .data_in(sw_394_data_out),
    .data_out(sw_395_data_out),
    .latch_enable_in(sw_394_latch_out),
    .latch_enable_out(sw_395_latch_out),
    .scan_select_in(sw_394_scan_out),
    .scan_select_out(sw_395_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_395_module_data_in[7] ,
    \sw_395_module_data_in[6] ,
    \sw_395_module_data_in[5] ,
    \sw_395_module_data_in[4] ,
    \sw_395_module_data_in[3] ,
    \sw_395_module_data_in[2] ,
    \sw_395_module_data_in[1] ,
    \sw_395_module_data_in[0] }),
    .module_data_out({\sw_395_module_data_out[7] ,
    \sw_395_module_data_out[6] ,
    \sw_395_module_data_out[5] ,
    \sw_395_module_data_out[4] ,
    \sw_395_module_data_out[3] ,
    \sw_395_module_data_out[2] ,
    \sw_395_module_data_out[1] ,
    \sw_395_module_data_out[0] }));
 scanchain scanchain_396 (.clk_in(sw_395_clk_out),
    .clk_out(sw_396_clk_out),
    .data_in(sw_395_data_out),
    .data_out(sw_396_data_out),
    .latch_enable_in(sw_395_latch_out),
    .latch_enable_out(sw_396_latch_out),
    .scan_select_in(sw_395_scan_out),
    .scan_select_out(sw_396_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_396_module_data_in[7] ,
    \sw_396_module_data_in[6] ,
    \sw_396_module_data_in[5] ,
    \sw_396_module_data_in[4] ,
    \sw_396_module_data_in[3] ,
    \sw_396_module_data_in[2] ,
    \sw_396_module_data_in[1] ,
    \sw_396_module_data_in[0] }),
    .module_data_out({\sw_396_module_data_out[7] ,
    \sw_396_module_data_out[6] ,
    \sw_396_module_data_out[5] ,
    \sw_396_module_data_out[4] ,
    \sw_396_module_data_out[3] ,
    \sw_396_module_data_out[2] ,
    \sw_396_module_data_out[1] ,
    \sw_396_module_data_out[0] }));
 scanchain scanchain_397 (.clk_in(sw_396_clk_out),
    .clk_out(sw_397_clk_out),
    .data_in(sw_396_data_out),
    .data_out(sw_397_data_out),
    .latch_enable_in(sw_396_latch_out),
    .latch_enable_out(sw_397_latch_out),
    .scan_select_in(sw_396_scan_out),
    .scan_select_out(sw_397_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_397_module_data_in[7] ,
    \sw_397_module_data_in[6] ,
    \sw_397_module_data_in[5] ,
    \sw_397_module_data_in[4] ,
    \sw_397_module_data_in[3] ,
    \sw_397_module_data_in[2] ,
    \sw_397_module_data_in[1] ,
    \sw_397_module_data_in[0] }),
    .module_data_out({\sw_397_module_data_out[7] ,
    \sw_397_module_data_out[6] ,
    \sw_397_module_data_out[5] ,
    \sw_397_module_data_out[4] ,
    \sw_397_module_data_out[3] ,
    \sw_397_module_data_out[2] ,
    \sw_397_module_data_out[1] ,
    \sw_397_module_data_out[0] }));
 scanchain scanchain_398 (.clk_in(sw_397_clk_out),
    .clk_out(sw_398_clk_out),
    .data_in(sw_397_data_out),
    .data_out(sw_398_data_out),
    .latch_enable_in(sw_397_latch_out),
    .latch_enable_out(sw_398_latch_out),
    .scan_select_in(sw_397_scan_out),
    .scan_select_out(sw_398_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_398_module_data_in[7] ,
    \sw_398_module_data_in[6] ,
    \sw_398_module_data_in[5] ,
    \sw_398_module_data_in[4] ,
    \sw_398_module_data_in[3] ,
    \sw_398_module_data_in[2] ,
    \sw_398_module_data_in[1] ,
    \sw_398_module_data_in[0] }),
    .module_data_out({\sw_398_module_data_out[7] ,
    \sw_398_module_data_out[6] ,
    \sw_398_module_data_out[5] ,
    \sw_398_module_data_out[4] ,
    \sw_398_module_data_out[3] ,
    \sw_398_module_data_out[2] ,
    \sw_398_module_data_out[1] ,
    \sw_398_module_data_out[0] }));
 scanchain scanchain_399 (.clk_in(sw_398_clk_out),
    .clk_out(sw_399_clk_out),
    .data_in(sw_398_data_out),
    .data_out(sw_399_data_out),
    .latch_enable_in(sw_398_latch_out),
    .latch_enable_out(sw_399_latch_out),
    .scan_select_in(sw_398_scan_out),
    .scan_select_out(sw_399_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_399_module_data_in[7] ,
    \sw_399_module_data_in[6] ,
    \sw_399_module_data_in[5] ,
    \sw_399_module_data_in[4] ,
    \sw_399_module_data_in[3] ,
    \sw_399_module_data_in[2] ,
    \sw_399_module_data_in[1] ,
    \sw_399_module_data_in[0] }),
    .module_data_out({\sw_399_module_data_out[7] ,
    \sw_399_module_data_out[6] ,
    \sw_399_module_data_out[5] ,
    \sw_399_module_data_out[4] ,
    \sw_399_module_data_out[3] ,
    \sw_399_module_data_out[2] ,
    \sw_399_module_data_out[1] ,
    \sw_399_module_data_out[0] }));
 scanchain scanchain_4 (.clk_in(sw_003_clk_out),
    .clk_out(sw_004_clk_out),
    .data_in(sw_003_data_out),
    .data_out(sw_004_data_out),
    .latch_enable_in(sw_003_latch_out),
    .latch_enable_out(sw_004_latch_out),
    .scan_select_in(sw_003_scan_out),
    .scan_select_out(sw_004_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_004_module_data_in[7] ,
    \sw_004_module_data_in[6] ,
    \sw_004_module_data_in[5] ,
    \sw_004_module_data_in[4] ,
    \sw_004_module_data_in[3] ,
    \sw_004_module_data_in[2] ,
    \sw_004_module_data_in[1] ,
    \sw_004_module_data_in[0] }),
    .module_data_out({\sw_004_module_data_out[7] ,
    \sw_004_module_data_out[6] ,
    \sw_004_module_data_out[5] ,
    \sw_004_module_data_out[4] ,
    \sw_004_module_data_out[3] ,
    \sw_004_module_data_out[2] ,
    \sw_004_module_data_out[1] ,
    \sw_004_module_data_out[0] }));
 scanchain scanchain_40 (.clk_in(sw_039_clk_out),
    .clk_out(sw_040_clk_out),
    .data_in(sw_039_data_out),
    .data_out(sw_040_data_out),
    .latch_enable_in(sw_039_latch_out),
    .latch_enable_out(sw_040_latch_out),
    .scan_select_in(sw_039_scan_out),
    .scan_select_out(sw_040_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_040_module_data_in[7] ,
    \sw_040_module_data_in[6] ,
    \sw_040_module_data_in[5] ,
    \sw_040_module_data_in[4] ,
    \sw_040_module_data_in[3] ,
    \sw_040_module_data_in[2] ,
    \sw_040_module_data_in[1] ,
    \sw_040_module_data_in[0] }),
    .module_data_out({\sw_040_module_data_out[7] ,
    \sw_040_module_data_out[6] ,
    \sw_040_module_data_out[5] ,
    \sw_040_module_data_out[4] ,
    \sw_040_module_data_out[3] ,
    \sw_040_module_data_out[2] ,
    \sw_040_module_data_out[1] ,
    \sw_040_module_data_out[0] }));
 scanchain scanchain_400 (.clk_in(sw_399_clk_out),
    .clk_out(sw_400_clk_out),
    .data_in(sw_399_data_out),
    .data_out(sw_400_data_out),
    .latch_enable_in(sw_399_latch_out),
    .latch_enable_out(sw_400_latch_out),
    .scan_select_in(sw_399_scan_out),
    .scan_select_out(sw_400_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_400_module_data_in[7] ,
    \sw_400_module_data_in[6] ,
    \sw_400_module_data_in[5] ,
    \sw_400_module_data_in[4] ,
    \sw_400_module_data_in[3] ,
    \sw_400_module_data_in[2] ,
    \sw_400_module_data_in[1] ,
    \sw_400_module_data_in[0] }),
    .module_data_out({\sw_400_module_data_out[7] ,
    \sw_400_module_data_out[6] ,
    \sw_400_module_data_out[5] ,
    \sw_400_module_data_out[4] ,
    \sw_400_module_data_out[3] ,
    \sw_400_module_data_out[2] ,
    \sw_400_module_data_out[1] ,
    \sw_400_module_data_out[0] }));
 scanchain scanchain_401 (.clk_in(sw_400_clk_out),
    .clk_out(sw_401_clk_out),
    .data_in(sw_400_data_out),
    .data_out(sw_401_data_out),
    .latch_enable_in(sw_400_latch_out),
    .latch_enable_out(sw_401_latch_out),
    .scan_select_in(sw_400_scan_out),
    .scan_select_out(sw_401_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_401_module_data_in[7] ,
    \sw_401_module_data_in[6] ,
    \sw_401_module_data_in[5] ,
    \sw_401_module_data_in[4] ,
    \sw_401_module_data_in[3] ,
    \sw_401_module_data_in[2] ,
    \sw_401_module_data_in[1] ,
    \sw_401_module_data_in[0] }),
    .module_data_out({\sw_401_module_data_out[7] ,
    \sw_401_module_data_out[6] ,
    \sw_401_module_data_out[5] ,
    \sw_401_module_data_out[4] ,
    \sw_401_module_data_out[3] ,
    \sw_401_module_data_out[2] ,
    \sw_401_module_data_out[1] ,
    \sw_401_module_data_out[0] }));
 scanchain scanchain_402 (.clk_in(sw_401_clk_out),
    .clk_out(sw_402_clk_out),
    .data_in(sw_401_data_out),
    .data_out(sw_402_data_out),
    .latch_enable_in(sw_401_latch_out),
    .latch_enable_out(sw_402_latch_out),
    .scan_select_in(sw_401_scan_out),
    .scan_select_out(sw_402_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_402_module_data_in[7] ,
    \sw_402_module_data_in[6] ,
    \sw_402_module_data_in[5] ,
    \sw_402_module_data_in[4] ,
    \sw_402_module_data_in[3] ,
    \sw_402_module_data_in[2] ,
    \sw_402_module_data_in[1] ,
    \sw_402_module_data_in[0] }),
    .module_data_out({\sw_402_module_data_out[7] ,
    \sw_402_module_data_out[6] ,
    \sw_402_module_data_out[5] ,
    \sw_402_module_data_out[4] ,
    \sw_402_module_data_out[3] ,
    \sw_402_module_data_out[2] ,
    \sw_402_module_data_out[1] ,
    \sw_402_module_data_out[0] }));
 scanchain scanchain_403 (.clk_in(sw_402_clk_out),
    .clk_out(sw_403_clk_out),
    .data_in(sw_402_data_out),
    .data_out(sw_403_data_out),
    .latch_enable_in(sw_402_latch_out),
    .latch_enable_out(sw_403_latch_out),
    .scan_select_in(sw_402_scan_out),
    .scan_select_out(sw_403_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_403_module_data_in[7] ,
    \sw_403_module_data_in[6] ,
    \sw_403_module_data_in[5] ,
    \sw_403_module_data_in[4] ,
    \sw_403_module_data_in[3] ,
    \sw_403_module_data_in[2] ,
    \sw_403_module_data_in[1] ,
    \sw_403_module_data_in[0] }),
    .module_data_out({\sw_403_module_data_out[7] ,
    \sw_403_module_data_out[6] ,
    \sw_403_module_data_out[5] ,
    \sw_403_module_data_out[4] ,
    \sw_403_module_data_out[3] ,
    \sw_403_module_data_out[2] ,
    \sw_403_module_data_out[1] ,
    \sw_403_module_data_out[0] }));
 scanchain scanchain_404 (.clk_in(sw_403_clk_out),
    .clk_out(sw_404_clk_out),
    .data_in(sw_403_data_out),
    .data_out(sw_404_data_out),
    .latch_enable_in(sw_403_latch_out),
    .latch_enable_out(sw_404_latch_out),
    .scan_select_in(sw_403_scan_out),
    .scan_select_out(sw_404_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_404_module_data_in[7] ,
    \sw_404_module_data_in[6] ,
    \sw_404_module_data_in[5] ,
    \sw_404_module_data_in[4] ,
    \sw_404_module_data_in[3] ,
    \sw_404_module_data_in[2] ,
    \sw_404_module_data_in[1] ,
    \sw_404_module_data_in[0] }),
    .module_data_out({\sw_404_module_data_out[7] ,
    \sw_404_module_data_out[6] ,
    \sw_404_module_data_out[5] ,
    \sw_404_module_data_out[4] ,
    \sw_404_module_data_out[3] ,
    \sw_404_module_data_out[2] ,
    \sw_404_module_data_out[1] ,
    \sw_404_module_data_out[0] }));
 scanchain scanchain_405 (.clk_in(sw_404_clk_out),
    .clk_out(sw_405_clk_out),
    .data_in(sw_404_data_out),
    .data_out(sw_405_data_out),
    .latch_enable_in(sw_404_latch_out),
    .latch_enable_out(sw_405_latch_out),
    .scan_select_in(sw_404_scan_out),
    .scan_select_out(sw_405_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_405_module_data_in[7] ,
    \sw_405_module_data_in[6] ,
    \sw_405_module_data_in[5] ,
    \sw_405_module_data_in[4] ,
    \sw_405_module_data_in[3] ,
    \sw_405_module_data_in[2] ,
    \sw_405_module_data_in[1] ,
    \sw_405_module_data_in[0] }),
    .module_data_out({\sw_405_module_data_out[7] ,
    \sw_405_module_data_out[6] ,
    \sw_405_module_data_out[5] ,
    \sw_405_module_data_out[4] ,
    \sw_405_module_data_out[3] ,
    \sw_405_module_data_out[2] ,
    \sw_405_module_data_out[1] ,
    \sw_405_module_data_out[0] }));
 scanchain scanchain_406 (.clk_in(sw_405_clk_out),
    .clk_out(sw_406_clk_out),
    .data_in(sw_405_data_out),
    .data_out(sw_406_data_out),
    .latch_enable_in(sw_405_latch_out),
    .latch_enable_out(sw_406_latch_out),
    .scan_select_in(sw_405_scan_out),
    .scan_select_out(sw_406_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_406_module_data_in[7] ,
    \sw_406_module_data_in[6] ,
    \sw_406_module_data_in[5] ,
    \sw_406_module_data_in[4] ,
    \sw_406_module_data_in[3] ,
    \sw_406_module_data_in[2] ,
    \sw_406_module_data_in[1] ,
    \sw_406_module_data_in[0] }),
    .module_data_out({\sw_406_module_data_out[7] ,
    \sw_406_module_data_out[6] ,
    \sw_406_module_data_out[5] ,
    \sw_406_module_data_out[4] ,
    \sw_406_module_data_out[3] ,
    \sw_406_module_data_out[2] ,
    \sw_406_module_data_out[1] ,
    \sw_406_module_data_out[0] }));
 scanchain scanchain_407 (.clk_in(sw_406_clk_out),
    .clk_out(sw_407_clk_out),
    .data_in(sw_406_data_out),
    .data_out(sw_407_data_out),
    .latch_enable_in(sw_406_latch_out),
    .latch_enable_out(sw_407_latch_out),
    .scan_select_in(sw_406_scan_out),
    .scan_select_out(sw_407_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_407_module_data_in[7] ,
    \sw_407_module_data_in[6] ,
    \sw_407_module_data_in[5] ,
    \sw_407_module_data_in[4] ,
    \sw_407_module_data_in[3] ,
    \sw_407_module_data_in[2] ,
    \sw_407_module_data_in[1] ,
    \sw_407_module_data_in[0] }),
    .module_data_out({\sw_407_module_data_out[7] ,
    \sw_407_module_data_out[6] ,
    \sw_407_module_data_out[5] ,
    \sw_407_module_data_out[4] ,
    \sw_407_module_data_out[3] ,
    \sw_407_module_data_out[2] ,
    \sw_407_module_data_out[1] ,
    \sw_407_module_data_out[0] }));
 scanchain scanchain_408 (.clk_in(sw_407_clk_out),
    .clk_out(sw_408_clk_out),
    .data_in(sw_407_data_out),
    .data_out(sw_408_data_out),
    .latch_enable_in(sw_407_latch_out),
    .latch_enable_out(sw_408_latch_out),
    .scan_select_in(sw_407_scan_out),
    .scan_select_out(sw_408_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_408_module_data_in[7] ,
    \sw_408_module_data_in[6] ,
    \sw_408_module_data_in[5] ,
    \sw_408_module_data_in[4] ,
    \sw_408_module_data_in[3] ,
    \sw_408_module_data_in[2] ,
    \sw_408_module_data_in[1] ,
    \sw_408_module_data_in[0] }),
    .module_data_out({\sw_408_module_data_out[7] ,
    \sw_408_module_data_out[6] ,
    \sw_408_module_data_out[5] ,
    \sw_408_module_data_out[4] ,
    \sw_408_module_data_out[3] ,
    \sw_408_module_data_out[2] ,
    \sw_408_module_data_out[1] ,
    \sw_408_module_data_out[0] }));
 scanchain scanchain_409 (.clk_in(sw_408_clk_out),
    .clk_out(sw_409_clk_out),
    .data_in(sw_408_data_out),
    .data_out(sw_409_data_out),
    .latch_enable_in(sw_408_latch_out),
    .latch_enable_out(sw_409_latch_out),
    .scan_select_in(sw_408_scan_out),
    .scan_select_out(sw_409_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_409_module_data_in[7] ,
    \sw_409_module_data_in[6] ,
    \sw_409_module_data_in[5] ,
    \sw_409_module_data_in[4] ,
    \sw_409_module_data_in[3] ,
    \sw_409_module_data_in[2] ,
    \sw_409_module_data_in[1] ,
    \sw_409_module_data_in[0] }),
    .module_data_out({\sw_409_module_data_out[7] ,
    \sw_409_module_data_out[6] ,
    \sw_409_module_data_out[5] ,
    \sw_409_module_data_out[4] ,
    \sw_409_module_data_out[3] ,
    \sw_409_module_data_out[2] ,
    \sw_409_module_data_out[1] ,
    \sw_409_module_data_out[0] }));
 scanchain scanchain_41 (.clk_in(sw_040_clk_out),
    .clk_out(sw_041_clk_out),
    .data_in(sw_040_data_out),
    .data_out(sw_041_data_out),
    .latch_enable_in(sw_040_latch_out),
    .latch_enable_out(sw_041_latch_out),
    .scan_select_in(sw_040_scan_out),
    .scan_select_out(sw_041_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_041_module_data_in[7] ,
    \sw_041_module_data_in[6] ,
    \sw_041_module_data_in[5] ,
    \sw_041_module_data_in[4] ,
    \sw_041_module_data_in[3] ,
    \sw_041_module_data_in[2] ,
    \sw_041_module_data_in[1] ,
    \sw_041_module_data_in[0] }),
    .module_data_out({\sw_041_module_data_out[7] ,
    \sw_041_module_data_out[6] ,
    \sw_041_module_data_out[5] ,
    \sw_041_module_data_out[4] ,
    \sw_041_module_data_out[3] ,
    \sw_041_module_data_out[2] ,
    \sw_041_module_data_out[1] ,
    \sw_041_module_data_out[0] }));
 scanchain scanchain_410 (.clk_in(sw_409_clk_out),
    .clk_out(sw_410_clk_out),
    .data_in(sw_409_data_out),
    .data_out(sw_410_data_out),
    .latch_enable_in(sw_409_latch_out),
    .latch_enable_out(sw_410_latch_out),
    .scan_select_in(sw_409_scan_out),
    .scan_select_out(sw_410_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_410_module_data_in[7] ,
    \sw_410_module_data_in[6] ,
    \sw_410_module_data_in[5] ,
    \sw_410_module_data_in[4] ,
    \sw_410_module_data_in[3] ,
    \sw_410_module_data_in[2] ,
    \sw_410_module_data_in[1] ,
    \sw_410_module_data_in[0] }),
    .module_data_out({\sw_410_module_data_out[7] ,
    \sw_410_module_data_out[6] ,
    \sw_410_module_data_out[5] ,
    \sw_410_module_data_out[4] ,
    \sw_410_module_data_out[3] ,
    \sw_410_module_data_out[2] ,
    \sw_410_module_data_out[1] ,
    \sw_410_module_data_out[0] }));
 scanchain scanchain_411 (.clk_in(sw_410_clk_out),
    .clk_out(sw_411_clk_out),
    .data_in(sw_410_data_out),
    .data_out(sw_411_data_out),
    .latch_enable_in(sw_410_latch_out),
    .latch_enable_out(sw_411_latch_out),
    .scan_select_in(sw_410_scan_out),
    .scan_select_out(sw_411_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_411_module_data_in[7] ,
    \sw_411_module_data_in[6] ,
    \sw_411_module_data_in[5] ,
    \sw_411_module_data_in[4] ,
    \sw_411_module_data_in[3] ,
    \sw_411_module_data_in[2] ,
    \sw_411_module_data_in[1] ,
    \sw_411_module_data_in[0] }),
    .module_data_out({\sw_411_module_data_out[7] ,
    \sw_411_module_data_out[6] ,
    \sw_411_module_data_out[5] ,
    \sw_411_module_data_out[4] ,
    \sw_411_module_data_out[3] ,
    \sw_411_module_data_out[2] ,
    \sw_411_module_data_out[1] ,
    \sw_411_module_data_out[0] }));
 scanchain scanchain_412 (.clk_in(sw_411_clk_out),
    .clk_out(sw_412_clk_out),
    .data_in(sw_411_data_out),
    .data_out(sw_412_data_out),
    .latch_enable_in(sw_411_latch_out),
    .latch_enable_out(sw_412_latch_out),
    .scan_select_in(sw_411_scan_out),
    .scan_select_out(sw_412_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_412_module_data_in[7] ,
    \sw_412_module_data_in[6] ,
    \sw_412_module_data_in[5] ,
    \sw_412_module_data_in[4] ,
    \sw_412_module_data_in[3] ,
    \sw_412_module_data_in[2] ,
    \sw_412_module_data_in[1] ,
    \sw_412_module_data_in[0] }),
    .module_data_out({\sw_412_module_data_out[7] ,
    \sw_412_module_data_out[6] ,
    \sw_412_module_data_out[5] ,
    \sw_412_module_data_out[4] ,
    \sw_412_module_data_out[3] ,
    \sw_412_module_data_out[2] ,
    \sw_412_module_data_out[1] ,
    \sw_412_module_data_out[0] }));
 scanchain scanchain_413 (.clk_in(sw_412_clk_out),
    .clk_out(sw_413_clk_out),
    .data_in(sw_412_data_out),
    .data_out(sw_413_data_out),
    .latch_enable_in(sw_412_latch_out),
    .latch_enable_out(sw_413_latch_out),
    .scan_select_in(sw_412_scan_out),
    .scan_select_out(sw_413_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_413_module_data_in[7] ,
    \sw_413_module_data_in[6] ,
    \sw_413_module_data_in[5] ,
    \sw_413_module_data_in[4] ,
    \sw_413_module_data_in[3] ,
    \sw_413_module_data_in[2] ,
    \sw_413_module_data_in[1] ,
    \sw_413_module_data_in[0] }),
    .module_data_out({\sw_413_module_data_out[7] ,
    \sw_413_module_data_out[6] ,
    \sw_413_module_data_out[5] ,
    \sw_413_module_data_out[4] ,
    \sw_413_module_data_out[3] ,
    \sw_413_module_data_out[2] ,
    \sw_413_module_data_out[1] ,
    \sw_413_module_data_out[0] }));
 scanchain scanchain_414 (.clk_in(sw_413_clk_out),
    .clk_out(sw_414_clk_out),
    .data_in(sw_413_data_out),
    .data_out(sw_414_data_out),
    .latch_enable_in(sw_413_latch_out),
    .latch_enable_out(sw_414_latch_out),
    .scan_select_in(sw_413_scan_out),
    .scan_select_out(sw_414_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_414_module_data_in[7] ,
    \sw_414_module_data_in[6] ,
    \sw_414_module_data_in[5] ,
    \sw_414_module_data_in[4] ,
    \sw_414_module_data_in[3] ,
    \sw_414_module_data_in[2] ,
    \sw_414_module_data_in[1] ,
    \sw_414_module_data_in[0] }),
    .module_data_out({\sw_414_module_data_out[7] ,
    \sw_414_module_data_out[6] ,
    \sw_414_module_data_out[5] ,
    \sw_414_module_data_out[4] ,
    \sw_414_module_data_out[3] ,
    \sw_414_module_data_out[2] ,
    \sw_414_module_data_out[1] ,
    \sw_414_module_data_out[0] }));
 scanchain scanchain_415 (.clk_in(sw_414_clk_out),
    .clk_out(sw_415_clk_out),
    .data_in(sw_414_data_out),
    .data_out(sw_415_data_out),
    .latch_enable_in(sw_414_latch_out),
    .latch_enable_out(sw_415_latch_out),
    .scan_select_in(sw_414_scan_out),
    .scan_select_out(sw_415_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_415_module_data_in[7] ,
    \sw_415_module_data_in[6] ,
    \sw_415_module_data_in[5] ,
    \sw_415_module_data_in[4] ,
    \sw_415_module_data_in[3] ,
    \sw_415_module_data_in[2] ,
    \sw_415_module_data_in[1] ,
    \sw_415_module_data_in[0] }),
    .module_data_out({\sw_415_module_data_out[7] ,
    \sw_415_module_data_out[6] ,
    \sw_415_module_data_out[5] ,
    \sw_415_module_data_out[4] ,
    \sw_415_module_data_out[3] ,
    \sw_415_module_data_out[2] ,
    \sw_415_module_data_out[1] ,
    \sw_415_module_data_out[0] }));
 scanchain scanchain_416 (.clk_in(sw_415_clk_out),
    .clk_out(sw_416_clk_out),
    .data_in(sw_415_data_out),
    .data_out(sw_416_data_out),
    .latch_enable_in(sw_415_latch_out),
    .latch_enable_out(sw_416_latch_out),
    .scan_select_in(sw_415_scan_out),
    .scan_select_out(sw_416_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_416_module_data_in[7] ,
    \sw_416_module_data_in[6] ,
    \sw_416_module_data_in[5] ,
    \sw_416_module_data_in[4] ,
    \sw_416_module_data_in[3] ,
    \sw_416_module_data_in[2] ,
    \sw_416_module_data_in[1] ,
    \sw_416_module_data_in[0] }),
    .module_data_out({\sw_416_module_data_out[7] ,
    \sw_416_module_data_out[6] ,
    \sw_416_module_data_out[5] ,
    \sw_416_module_data_out[4] ,
    \sw_416_module_data_out[3] ,
    \sw_416_module_data_out[2] ,
    \sw_416_module_data_out[1] ,
    \sw_416_module_data_out[0] }));
 scanchain scanchain_417 (.clk_in(sw_416_clk_out),
    .clk_out(sw_417_clk_out),
    .data_in(sw_416_data_out),
    .data_out(sw_417_data_out),
    .latch_enable_in(sw_416_latch_out),
    .latch_enable_out(sw_417_latch_out),
    .scan_select_in(sw_416_scan_out),
    .scan_select_out(sw_417_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_417_module_data_in[7] ,
    \sw_417_module_data_in[6] ,
    \sw_417_module_data_in[5] ,
    \sw_417_module_data_in[4] ,
    \sw_417_module_data_in[3] ,
    \sw_417_module_data_in[2] ,
    \sw_417_module_data_in[1] ,
    \sw_417_module_data_in[0] }),
    .module_data_out({\sw_417_module_data_out[7] ,
    \sw_417_module_data_out[6] ,
    \sw_417_module_data_out[5] ,
    \sw_417_module_data_out[4] ,
    \sw_417_module_data_out[3] ,
    \sw_417_module_data_out[2] ,
    \sw_417_module_data_out[1] ,
    \sw_417_module_data_out[0] }));
 scanchain scanchain_418 (.clk_in(sw_417_clk_out),
    .clk_out(sw_418_clk_out),
    .data_in(sw_417_data_out),
    .data_out(sw_418_data_out),
    .latch_enable_in(sw_417_latch_out),
    .latch_enable_out(sw_418_latch_out),
    .scan_select_in(sw_417_scan_out),
    .scan_select_out(sw_418_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_418_module_data_in[7] ,
    \sw_418_module_data_in[6] ,
    \sw_418_module_data_in[5] ,
    \sw_418_module_data_in[4] ,
    \sw_418_module_data_in[3] ,
    \sw_418_module_data_in[2] ,
    \sw_418_module_data_in[1] ,
    \sw_418_module_data_in[0] }),
    .module_data_out({\sw_418_module_data_out[7] ,
    \sw_418_module_data_out[6] ,
    \sw_418_module_data_out[5] ,
    \sw_418_module_data_out[4] ,
    \sw_418_module_data_out[3] ,
    \sw_418_module_data_out[2] ,
    \sw_418_module_data_out[1] ,
    \sw_418_module_data_out[0] }));
 scanchain scanchain_419 (.clk_in(sw_418_clk_out),
    .clk_out(sw_419_clk_out),
    .data_in(sw_418_data_out),
    .data_out(sw_419_data_out),
    .latch_enable_in(sw_418_latch_out),
    .latch_enable_out(sw_419_latch_out),
    .scan_select_in(sw_418_scan_out),
    .scan_select_out(sw_419_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_419_module_data_in[7] ,
    \sw_419_module_data_in[6] ,
    \sw_419_module_data_in[5] ,
    \sw_419_module_data_in[4] ,
    \sw_419_module_data_in[3] ,
    \sw_419_module_data_in[2] ,
    \sw_419_module_data_in[1] ,
    \sw_419_module_data_in[0] }),
    .module_data_out({\sw_419_module_data_out[7] ,
    \sw_419_module_data_out[6] ,
    \sw_419_module_data_out[5] ,
    \sw_419_module_data_out[4] ,
    \sw_419_module_data_out[3] ,
    \sw_419_module_data_out[2] ,
    \sw_419_module_data_out[1] ,
    \sw_419_module_data_out[0] }));
 scanchain scanchain_42 (.clk_in(sw_041_clk_out),
    .clk_out(sw_042_clk_out),
    .data_in(sw_041_data_out),
    .data_out(sw_042_data_out),
    .latch_enable_in(sw_041_latch_out),
    .latch_enable_out(sw_042_latch_out),
    .scan_select_in(sw_041_scan_out),
    .scan_select_out(sw_042_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_042_module_data_in[7] ,
    \sw_042_module_data_in[6] ,
    \sw_042_module_data_in[5] ,
    \sw_042_module_data_in[4] ,
    \sw_042_module_data_in[3] ,
    \sw_042_module_data_in[2] ,
    \sw_042_module_data_in[1] ,
    \sw_042_module_data_in[0] }),
    .module_data_out({\sw_042_module_data_out[7] ,
    \sw_042_module_data_out[6] ,
    \sw_042_module_data_out[5] ,
    \sw_042_module_data_out[4] ,
    \sw_042_module_data_out[3] ,
    \sw_042_module_data_out[2] ,
    \sw_042_module_data_out[1] ,
    \sw_042_module_data_out[0] }));
 scanchain scanchain_420 (.clk_in(sw_419_clk_out),
    .clk_out(sw_420_clk_out),
    .data_in(sw_419_data_out),
    .data_out(sw_420_data_out),
    .latch_enable_in(sw_419_latch_out),
    .latch_enable_out(sw_420_latch_out),
    .scan_select_in(sw_419_scan_out),
    .scan_select_out(sw_420_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_420_module_data_in[7] ,
    \sw_420_module_data_in[6] ,
    \sw_420_module_data_in[5] ,
    \sw_420_module_data_in[4] ,
    \sw_420_module_data_in[3] ,
    \sw_420_module_data_in[2] ,
    \sw_420_module_data_in[1] ,
    \sw_420_module_data_in[0] }),
    .module_data_out({\sw_420_module_data_out[7] ,
    \sw_420_module_data_out[6] ,
    \sw_420_module_data_out[5] ,
    \sw_420_module_data_out[4] ,
    \sw_420_module_data_out[3] ,
    \sw_420_module_data_out[2] ,
    \sw_420_module_data_out[1] ,
    \sw_420_module_data_out[0] }));
 scanchain scanchain_421 (.clk_in(sw_420_clk_out),
    .clk_out(sw_421_clk_out),
    .data_in(sw_420_data_out),
    .data_out(sw_421_data_out),
    .latch_enable_in(sw_420_latch_out),
    .latch_enable_out(sw_421_latch_out),
    .scan_select_in(sw_420_scan_out),
    .scan_select_out(sw_421_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_421_module_data_in[7] ,
    \sw_421_module_data_in[6] ,
    \sw_421_module_data_in[5] ,
    \sw_421_module_data_in[4] ,
    \sw_421_module_data_in[3] ,
    \sw_421_module_data_in[2] ,
    \sw_421_module_data_in[1] ,
    \sw_421_module_data_in[0] }),
    .module_data_out({\sw_421_module_data_out[7] ,
    \sw_421_module_data_out[6] ,
    \sw_421_module_data_out[5] ,
    \sw_421_module_data_out[4] ,
    \sw_421_module_data_out[3] ,
    \sw_421_module_data_out[2] ,
    \sw_421_module_data_out[1] ,
    \sw_421_module_data_out[0] }));
 scanchain scanchain_422 (.clk_in(sw_421_clk_out),
    .clk_out(sw_422_clk_out),
    .data_in(sw_421_data_out),
    .data_out(sw_422_data_out),
    .latch_enable_in(sw_421_latch_out),
    .latch_enable_out(sw_422_latch_out),
    .scan_select_in(sw_421_scan_out),
    .scan_select_out(sw_422_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_422_module_data_in[7] ,
    \sw_422_module_data_in[6] ,
    \sw_422_module_data_in[5] ,
    \sw_422_module_data_in[4] ,
    \sw_422_module_data_in[3] ,
    \sw_422_module_data_in[2] ,
    \sw_422_module_data_in[1] ,
    \sw_422_module_data_in[0] }),
    .module_data_out({\sw_422_module_data_out[7] ,
    \sw_422_module_data_out[6] ,
    \sw_422_module_data_out[5] ,
    \sw_422_module_data_out[4] ,
    \sw_422_module_data_out[3] ,
    \sw_422_module_data_out[2] ,
    \sw_422_module_data_out[1] ,
    \sw_422_module_data_out[0] }));
 scanchain scanchain_423 (.clk_in(sw_422_clk_out),
    .clk_out(sw_423_clk_out),
    .data_in(sw_422_data_out),
    .data_out(sw_423_data_out),
    .latch_enable_in(sw_422_latch_out),
    .latch_enable_out(sw_423_latch_out),
    .scan_select_in(sw_422_scan_out),
    .scan_select_out(sw_423_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_423_module_data_in[7] ,
    \sw_423_module_data_in[6] ,
    \sw_423_module_data_in[5] ,
    \sw_423_module_data_in[4] ,
    \sw_423_module_data_in[3] ,
    \sw_423_module_data_in[2] ,
    \sw_423_module_data_in[1] ,
    \sw_423_module_data_in[0] }),
    .module_data_out({\sw_423_module_data_out[7] ,
    \sw_423_module_data_out[6] ,
    \sw_423_module_data_out[5] ,
    \sw_423_module_data_out[4] ,
    \sw_423_module_data_out[3] ,
    \sw_423_module_data_out[2] ,
    \sw_423_module_data_out[1] ,
    \sw_423_module_data_out[0] }));
 scanchain scanchain_424 (.clk_in(sw_423_clk_out),
    .clk_out(sw_424_clk_out),
    .data_in(sw_423_data_out),
    .data_out(sw_424_data_out),
    .latch_enable_in(sw_423_latch_out),
    .latch_enable_out(sw_424_latch_out),
    .scan_select_in(sw_423_scan_out),
    .scan_select_out(sw_424_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_424_module_data_in[7] ,
    \sw_424_module_data_in[6] ,
    \sw_424_module_data_in[5] ,
    \sw_424_module_data_in[4] ,
    \sw_424_module_data_in[3] ,
    \sw_424_module_data_in[2] ,
    \sw_424_module_data_in[1] ,
    \sw_424_module_data_in[0] }),
    .module_data_out({\sw_424_module_data_out[7] ,
    \sw_424_module_data_out[6] ,
    \sw_424_module_data_out[5] ,
    \sw_424_module_data_out[4] ,
    \sw_424_module_data_out[3] ,
    \sw_424_module_data_out[2] ,
    \sw_424_module_data_out[1] ,
    \sw_424_module_data_out[0] }));
 scanchain scanchain_425 (.clk_in(sw_424_clk_out),
    .clk_out(sw_425_clk_out),
    .data_in(sw_424_data_out),
    .data_out(sw_425_data_out),
    .latch_enable_in(sw_424_latch_out),
    .latch_enable_out(sw_425_latch_out),
    .scan_select_in(sw_424_scan_out),
    .scan_select_out(sw_425_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_425_module_data_in[7] ,
    \sw_425_module_data_in[6] ,
    \sw_425_module_data_in[5] ,
    \sw_425_module_data_in[4] ,
    \sw_425_module_data_in[3] ,
    \sw_425_module_data_in[2] ,
    \sw_425_module_data_in[1] ,
    \sw_425_module_data_in[0] }),
    .module_data_out({\sw_425_module_data_out[7] ,
    \sw_425_module_data_out[6] ,
    \sw_425_module_data_out[5] ,
    \sw_425_module_data_out[4] ,
    \sw_425_module_data_out[3] ,
    \sw_425_module_data_out[2] ,
    \sw_425_module_data_out[1] ,
    \sw_425_module_data_out[0] }));
 scanchain scanchain_426 (.clk_in(sw_425_clk_out),
    .clk_out(sw_426_clk_out),
    .data_in(sw_425_data_out),
    .data_out(sw_426_data_out),
    .latch_enable_in(sw_425_latch_out),
    .latch_enable_out(sw_426_latch_out),
    .scan_select_in(sw_425_scan_out),
    .scan_select_out(sw_426_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_426_module_data_in[7] ,
    \sw_426_module_data_in[6] ,
    \sw_426_module_data_in[5] ,
    \sw_426_module_data_in[4] ,
    \sw_426_module_data_in[3] ,
    \sw_426_module_data_in[2] ,
    \sw_426_module_data_in[1] ,
    \sw_426_module_data_in[0] }),
    .module_data_out({\sw_426_module_data_out[7] ,
    \sw_426_module_data_out[6] ,
    \sw_426_module_data_out[5] ,
    \sw_426_module_data_out[4] ,
    \sw_426_module_data_out[3] ,
    \sw_426_module_data_out[2] ,
    \sw_426_module_data_out[1] ,
    \sw_426_module_data_out[0] }));
 scanchain scanchain_427 (.clk_in(sw_426_clk_out),
    .clk_out(sw_427_clk_out),
    .data_in(sw_426_data_out),
    .data_out(sw_427_data_out),
    .latch_enable_in(sw_426_latch_out),
    .latch_enable_out(sw_427_latch_out),
    .scan_select_in(sw_426_scan_out),
    .scan_select_out(sw_427_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_427_module_data_in[7] ,
    \sw_427_module_data_in[6] ,
    \sw_427_module_data_in[5] ,
    \sw_427_module_data_in[4] ,
    \sw_427_module_data_in[3] ,
    \sw_427_module_data_in[2] ,
    \sw_427_module_data_in[1] ,
    \sw_427_module_data_in[0] }),
    .module_data_out({\sw_427_module_data_out[7] ,
    \sw_427_module_data_out[6] ,
    \sw_427_module_data_out[5] ,
    \sw_427_module_data_out[4] ,
    \sw_427_module_data_out[3] ,
    \sw_427_module_data_out[2] ,
    \sw_427_module_data_out[1] ,
    \sw_427_module_data_out[0] }));
 scanchain scanchain_428 (.clk_in(sw_427_clk_out),
    .clk_out(sw_428_clk_out),
    .data_in(sw_427_data_out),
    .data_out(sw_428_data_out),
    .latch_enable_in(sw_427_latch_out),
    .latch_enable_out(sw_428_latch_out),
    .scan_select_in(sw_427_scan_out),
    .scan_select_out(sw_428_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_428_module_data_in[7] ,
    \sw_428_module_data_in[6] ,
    \sw_428_module_data_in[5] ,
    \sw_428_module_data_in[4] ,
    \sw_428_module_data_in[3] ,
    \sw_428_module_data_in[2] ,
    \sw_428_module_data_in[1] ,
    \sw_428_module_data_in[0] }),
    .module_data_out({\sw_428_module_data_out[7] ,
    \sw_428_module_data_out[6] ,
    \sw_428_module_data_out[5] ,
    \sw_428_module_data_out[4] ,
    \sw_428_module_data_out[3] ,
    \sw_428_module_data_out[2] ,
    \sw_428_module_data_out[1] ,
    \sw_428_module_data_out[0] }));
 scanchain scanchain_429 (.clk_in(sw_428_clk_out),
    .clk_out(sw_429_clk_out),
    .data_in(sw_428_data_out),
    .data_out(sw_429_data_out),
    .latch_enable_in(sw_428_latch_out),
    .latch_enable_out(sw_429_latch_out),
    .scan_select_in(sw_428_scan_out),
    .scan_select_out(sw_429_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_429_module_data_in[7] ,
    \sw_429_module_data_in[6] ,
    \sw_429_module_data_in[5] ,
    \sw_429_module_data_in[4] ,
    \sw_429_module_data_in[3] ,
    \sw_429_module_data_in[2] ,
    \sw_429_module_data_in[1] ,
    \sw_429_module_data_in[0] }),
    .module_data_out({\sw_429_module_data_out[7] ,
    \sw_429_module_data_out[6] ,
    \sw_429_module_data_out[5] ,
    \sw_429_module_data_out[4] ,
    \sw_429_module_data_out[3] ,
    \sw_429_module_data_out[2] ,
    \sw_429_module_data_out[1] ,
    \sw_429_module_data_out[0] }));
 scanchain scanchain_43 (.clk_in(sw_042_clk_out),
    .clk_out(sw_043_clk_out),
    .data_in(sw_042_data_out),
    .data_out(sw_043_data_out),
    .latch_enable_in(sw_042_latch_out),
    .latch_enable_out(sw_043_latch_out),
    .scan_select_in(sw_042_scan_out),
    .scan_select_out(sw_043_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_043_module_data_in[7] ,
    \sw_043_module_data_in[6] ,
    \sw_043_module_data_in[5] ,
    \sw_043_module_data_in[4] ,
    \sw_043_module_data_in[3] ,
    \sw_043_module_data_in[2] ,
    \sw_043_module_data_in[1] ,
    \sw_043_module_data_in[0] }),
    .module_data_out({\sw_043_module_data_out[7] ,
    \sw_043_module_data_out[6] ,
    \sw_043_module_data_out[5] ,
    \sw_043_module_data_out[4] ,
    \sw_043_module_data_out[3] ,
    \sw_043_module_data_out[2] ,
    \sw_043_module_data_out[1] ,
    \sw_043_module_data_out[0] }));
 scanchain scanchain_430 (.clk_in(sw_429_clk_out),
    .clk_out(sw_430_clk_out),
    .data_in(sw_429_data_out),
    .data_out(sw_430_data_out),
    .latch_enable_in(sw_429_latch_out),
    .latch_enable_out(sw_430_latch_out),
    .scan_select_in(sw_429_scan_out),
    .scan_select_out(sw_430_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_430_module_data_in[7] ,
    \sw_430_module_data_in[6] ,
    \sw_430_module_data_in[5] ,
    \sw_430_module_data_in[4] ,
    \sw_430_module_data_in[3] ,
    \sw_430_module_data_in[2] ,
    \sw_430_module_data_in[1] ,
    \sw_430_module_data_in[0] }),
    .module_data_out({\sw_430_module_data_out[7] ,
    \sw_430_module_data_out[6] ,
    \sw_430_module_data_out[5] ,
    \sw_430_module_data_out[4] ,
    \sw_430_module_data_out[3] ,
    \sw_430_module_data_out[2] ,
    \sw_430_module_data_out[1] ,
    \sw_430_module_data_out[0] }));
 scanchain scanchain_431 (.clk_in(sw_430_clk_out),
    .clk_out(sw_431_clk_out),
    .data_in(sw_430_data_out),
    .data_out(sw_431_data_out),
    .latch_enable_in(sw_430_latch_out),
    .latch_enable_out(sw_431_latch_out),
    .scan_select_in(sw_430_scan_out),
    .scan_select_out(sw_431_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_431_module_data_in[7] ,
    \sw_431_module_data_in[6] ,
    \sw_431_module_data_in[5] ,
    \sw_431_module_data_in[4] ,
    \sw_431_module_data_in[3] ,
    \sw_431_module_data_in[2] ,
    \sw_431_module_data_in[1] ,
    \sw_431_module_data_in[0] }),
    .module_data_out({\sw_431_module_data_out[7] ,
    \sw_431_module_data_out[6] ,
    \sw_431_module_data_out[5] ,
    \sw_431_module_data_out[4] ,
    \sw_431_module_data_out[3] ,
    \sw_431_module_data_out[2] ,
    \sw_431_module_data_out[1] ,
    \sw_431_module_data_out[0] }));
 scanchain scanchain_432 (.clk_in(sw_431_clk_out),
    .clk_out(sw_432_clk_out),
    .data_in(sw_431_data_out),
    .data_out(sw_432_data_out),
    .latch_enable_in(sw_431_latch_out),
    .latch_enable_out(sw_432_latch_out),
    .scan_select_in(sw_431_scan_out),
    .scan_select_out(sw_432_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_432_module_data_in[7] ,
    \sw_432_module_data_in[6] ,
    \sw_432_module_data_in[5] ,
    \sw_432_module_data_in[4] ,
    \sw_432_module_data_in[3] ,
    \sw_432_module_data_in[2] ,
    \sw_432_module_data_in[1] ,
    \sw_432_module_data_in[0] }),
    .module_data_out({\sw_432_module_data_out[7] ,
    \sw_432_module_data_out[6] ,
    \sw_432_module_data_out[5] ,
    \sw_432_module_data_out[4] ,
    \sw_432_module_data_out[3] ,
    \sw_432_module_data_out[2] ,
    \sw_432_module_data_out[1] ,
    \sw_432_module_data_out[0] }));
 scanchain scanchain_433 (.clk_in(sw_432_clk_out),
    .clk_out(sw_433_clk_out),
    .data_in(sw_432_data_out),
    .data_out(sw_433_data_out),
    .latch_enable_in(sw_432_latch_out),
    .latch_enable_out(sw_433_latch_out),
    .scan_select_in(sw_432_scan_out),
    .scan_select_out(sw_433_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_433_module_data_in[7] ,
    \sw_433_module_data_in[6] ,
    \sw_433_module_data_in[5] ,
    \sw_433_module_data_in[4] ,
    \sw_433_module_data_in[3] ,
    \sw_433_module_data_in[2] ,
    \sw_433_module_data_in[1] ,
    \sw_433_module_data_in[0] }),
    .module_data_out({\sw_433_module_data_out[7] ,
    \sw_433_module_data_out[6] ,
    \sw_433_module_data_out[5] ,
    \sw_433_module_data_out[4] ,
    \sw_433_module_data_out[3] ,
    \sw_433_module_data_out[2] ,
    \sw_433_module_data_out[1] ,
    \sw_433_module_data_out[0] }));
 scanchain scanchain_434 (.clk_in(sw_433_clk_out),
    .clk_out(sw_434_clk_out),
    .data_in(sw_433_data_out),
    .data_out(sw_434_data_out),
    .latch_enable_in(sw_433_latch_out),
    .latch_enable_out(sw_434_latch_out),
    .scan_select_in(sw_433_scan_out),
    .scan_select_out(sw_434_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_434_module_data_in[7] ,
    \sw_434_module_data_in[6] ,
    \sw_434_module_data_in[5] ,
    \sw_434_module_data_in[4] ,
    \sw_434_module_data_in[3] ,
    \sw_434_module_data_in[2] ,
    \sw_434_module_data_in[1] ,
    \sw_434_module_data_in[0] }),
    .module_data_out({\sw_434_module_data_out[7] ,
    \sw_434_module_data_out[6] ,
    \sw_434_module_data_out[5] ,
    \sw_434_module_data_out[4] ,
    \sw_434_module_data_out[3] ,
    \sw_434_module_data_out[2] ,
    \sw_434_module_data_out[1] ,
    \sw_434_module_data_out[0] }));
 scanchain scanchain_435 (.clk_in(sw_434_clk_out),
    .clk_out(sw_435_clk_out),
    .data_in(sw_434_data_out),
    .data_out(sw_435_data_out),
    .latch_enable_in(sw_434_latch_out),
    .latch_enable_out(sw_435_latch_out),
    .scan_select_in(sw_434_scan_out),
    .scan_select_out(sw_435_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_435_module_data_in[7] ,
    \sw_435_module_data_in[6] ,
    \sw_435_module_data_in[5] ,
    \sw_435_module_data_in[4] ,
    \sw_435_module_data_in[3] ,
    \sw_435_module_data_in[2] ,
    \sw_435_module_data_in[1] ,
    \sw_435_module_data_in[0] }),
    .module_data_out({\sw_435_module_data_out[7] ,
    \sw_435_module_data_out[6] ,
    \sw_435_module_data_out[5] ,
    \sw_435_module_data_out[4] ,
    \sw_435_module_data_out[3] ,
    \sw_435_module_data_out[2] ,
    \sw_435_module_data_out[1] ,
    \sw_435_module_data_out[0] }));
 scanchain scanchain_436 (.clk_in(sw_435_clk_out),
    .clk_out(sw_436_clk_out),
    .data_in(sw_435_data_out),
    .data_out(sw_436_data_out),
    .latch_enable_in(sw_435_latch_out),
    .latch_enable_out(sw_436_latch_out),
    .scan_select_in(sw_435_scan_out),
    .scan_select_out(sw_436_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_436_module_data_in[7] ,
    \sw_436_module_data_in[6] ,
    \sw_436_module_data_in[5] ,
    \sw_436_module_data_in[4] ,
    \sw_436_module_data_in[3] ,
    \sw_436_module_data_in[2] ,
    \sw_436_module_data_in[1] ,
    \sw_436_module_data_in[0] }),
    .module_data_out({\sw_436_module_data_out[7] ,
    \sw_436_module_data_out[6] ,
    \sw_436_module_data_out[5] ,
    \sw_436_module_data_out[4] ,
    \sw_436_module_data_out[3] ,
    \sw_436_module_data_out[2] ,
    \sw_436_module_data_out[1] ,
    \sw_436_module_data_out[0] }));
 scanchain scanchain_437 (.clk_in(sw_436_clk_out),
    .clk_out(sw_437_clk_out),
    .data_in(sw_436_data_out),
    .data_out(sw_437_data_out),
    .latch_enable_in(sw_436_latch_out),
    .latch_enable_out(sw_437_latch_out),
    .scan_select_in(sw_436_scan_out),
    .scan_select_out(sw_437_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_437_module_data_in[7] ,
    \sw_437_module_data_in[6] ,
    \sw_437_module_data_in[5] ,
    \sw_437_module_data_in[4] ,
    \sw_437_module_data_in[3] ,
    \sw_437_module_data_in[2] ,
    \sw_437_module_data_in[1] ,
    \sw_437_module_data_in[0] }),
    .module_data_out({\sw_437_module_data_out[7] ,
    \sw_437_module_data_out[6] ,
    \sw_437_module_data_out[5] ,
    \sw_437_module_data_out[4] ,
    \sw_437_module_data_out[3] ,
    \sw_437_module_data_out[2] ,
    \sw_437_module_data_out[1] ,
    \sw_437_module_data_out[0] }));
 scanchain scanchain_438 (.clk_in(sw_437_clk_out),
    .clk_out(sw_438_clk_out),
    .data_in(sw_437_data_out),
    .data_out(sw_438_data_out),
    .latch_enable_in(sw_437_latch_out),
    .latch_enable_out(sw_438_latch_out),
    .scan_select_in(sw_437_scan_out),
    .scan_select_out(sw_438_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_438_module_data_in[7] ,
    \sw_438_module_data_in[6] ,
    \sw_438_module_data_in[5] ,
    \sw_438_module_data_in[4] ,
    \sw_438_module_data_in[3] ,
    \sw_438_module_data_in[2] ,
    \sw_438_module_data_in[1] ,
    \sw_438_module_data_in[0] }),
    .module_data_out({\sw_438_module_data_out[7] ,
    \sw_438_module_data_out[6] ,
    \sw_438_module_data_out[5] ,
    \sw_438_module_data_out[4] ,
    \sw_438_module_data_out[3] ,
    \sw_438_module_data_out[2] ,
    \sw_438_module_data_out[1] ,
    \sw_438_module_data_out[0] }));
 scanchain scanchain_439 (.clk_in(sw_438_clk_out),
    .clk_out(sw_439_clk_out),
    .data_in(sw_438_data_out),
    .data_out(sw_439_data_out),
    .latch_enable_in(sw_438_latch_out),
    .latch_enable_out(sw_439_latch_out),
    .scan_select_in(sw_438_scan_out),
    .scan_select_out(sw_439_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_439_module_data_in[7] ,
    \sw_439_module_data_in[6] ,
    \sw_439_module_data_in[5] ,
    \sw_439_module_data_in[4] ,
    \sw_439_module_data_in[3] ,
    \sw_439_module_data_in[2] ,
    \sw_439_module_data_in[1] ,
    \sw_439_module_data_in[0] }),
    .module_data_out({\sw_439_module_data_out[7] ,
    \sw_439_module_data_out[6] ,
    \sw_439_module_data_out[5] ,
    \sw_439_module_data_out[4] ,
    \sw_439_module_data_out[3] ,
    \sw_439_module_data_out[2] ,
    \sw_439_module_data_out[1] ,
    \sw_439_module_data_out[0] }));
 scanchain scanchain_44 (.clk_in(sw_043_clk_out),
    .clk_out(sw_044_clk_out),
    .data_in(sw_043_data_out),
    .data_out(sw_044_data_out),
    .latch_enable_in(sw_043_latch_out),
    .latch_enable_out(sw_044_latch_out),
    .scan_select_in(sw_043_scan_out),
    .scan_select_out(sw_044_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_044_module_data_in[7] ,
    \sw_044_module_data_in[6] ,
    \sw_044_module_data_in[5] ,
    \sw_044_module_data_in[4] ,
    \sw_044_module_data_in[3] ,
    \sw_044_module_data_in[2] ,
    \sw_044_module_data_in[1] ,
    \sw_044_module_data_in[0] }),
    .module_data_out({\sw_044_module_data_out[7] ,
    \sw_044_module_data_out[6] ,
    \sw_044_module_data_out[5] ,
    \sw_044_module_data_out[4] ,
    \sw_044_module_data_out[3] ,
    \sw_044_module_data_out[2] ,
    \sw_044_module_data_out[1] ,
    \sw_044_module_data_out[0] }));
 scanchain scanchain_440 (.clk_in(sw_439_clk_out),
    .clk_out(sw_440_clk_out),
    .data_in(sw_439_data_out),
    .data_out(sw_440_data_out),
    .latch_enable_in(sw_439_latch_out),
    .latch_enable_out(sw_440_latch_out),
    .scan_select_in(sw_439_scan_out),
    .scan_select_out(sw_440_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_440_module_data_in[7] ,
    \sw_440_module_data_in[6] ,
    \sw_440_module_data_in[5] ,
    \sw_440_module_data_in[4] ,
    \sw_440_module_data_in[3] ,
    \sw_440_module_data_in[2] ,
    \sw_440_module_data_in[1] ,
    \sw_440_module_data_in[0] }),
    .module_data_out({\sw_440_module_data_out[7] ,
    \sw_440_module_data_out[6] ,
    \sw_440_module_data_out[5] ,
    \sw_440_module_data_out[4] ,
    \sw_440_module_data_out[3] ,
    \sw_440_module_data_out[2] ,
    \sw_440_module_data_out[1] ,
    \sw_440_module_data_out[0] }));
 scanchain scanchain_441 (.clk_in(sw_440_clk_out),
    .clk_out(sw_441_clk_out),
    .data_in(sw_440_data_out),
    .data_out(sw_441_data_out),
    .latch_enable_in(sw_440_latch_out),
    .latch_enable_out(sw_441_latch_out),
    .scan_select_in(sw_440_scan_out),
    .scan_select_out(sw_441_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_441_module_data_in[7] ,
    \sw_441_module_data_in[6] ,
    \sw_441_module_data_in[5] ,
    \sw_441_module_data_in[4] ,
    \sw_441_module_data_in[3] ,
    \sw_441_module_data_in[2] ,
    \sw_441_module_data_in[1] ,
    \sw_441_module_data_in[0] }),
    .module_data_out({\sw_441_module_data_out[7] ,
    \sw_441_module_data_out[6] ,
    \sw_441_module_data_out[5] ,
    \sw_441_module_data_out[4] ,
    \sw_441_module_data_out[3] ,
    \sw_441_module_data_out[2] ,
    \sw_441_module_data_out[1] ,
    \sw_441_module_data_out[0] }));
 scanchain scanchain_442 (.clk_in(sw_441_clk_out),
    .clk_out(sw_442_clk_out),
    .data_in(sw_441_data_out),
    .data_out(sw_442_data_out),
    .latch_enable_in(sw_441_latch_out),
    .latch_enable_out(sw_442_latch_out),
    .scan_select_in(sw_441_scan_out),
    .scan_select_out(sw_442_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_442_module_data_in[7] ,
    \sw_442_module_data_in[6] ,
    \sw_442_module_data_in[5] ,
    \sw_442_module_data_in[4] ,
    \sw_442_module_data_in[3] ,
    \sw_442_module_data_in[2] ,
    \sw_442_module_data_in[1] ,
    \sw_442_module_data_in[0] }),
    .module_data_out({\sw_442_module_data_out[7] ,
    \sw_442_module_data_out[6] ,
    \sw_442_module_data_out[5] ,
    \sw_442_module_data_out[4] ,
    \sw_442_module_data_out[3] ,
    \sw_442_module_data_out[2] ,
    \sw_442_module_data_out[1] ,
    \sw_442_module_data_out[0] }));
 scanchain scanchain_443 (.clk_in(sw_442_clk_out),
    .clk_out(sw_443_clk_out),
    .data_in(sw_442_data_out),
    .data_out(sw_443_data_out),
    .latch_enable_in(sw_442_latch_out),
    .latch_enable_out(sw_443_latch_out),
    .scan_select_in(sw_442_scan_out),
    .scan_select_out(sw_443_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_443_module_data_in[7] ,
    \sw_443_module_data_in[6] ,
    \sw_443_module_data_in[5] ,
    \sw_443_module_data_in[4] ,
    \sw_443_module_data_in[3] ,
    \sw_443_module_data_in[2] ,
    \sw_443_module_data_in[1] ,
    \sw_443_module_data_in[0] }),
    .module_data_out({\sw_443_module_data_out[7] ,
    \sw_443_module_data_out[6] ,
    \sw_443_module_data_out[5] ,
    \sw_443_module_data_out[4] ,
    \sw_443_module_data_out[3] ,
    \sw_443_module_data_out[2] ,
    \sw_443_module_data_out[1] ,
    \sw_443_module_data_out[0] }));
 scanchain scanchain_444 (.clk_in(sw_443_clk_out),
    .clk_out(sw_444_clk_out),
    .data_in(sw_443_data_out),
    .data_out(sw_444_data_out),
    .latch_enable_in(sw_443_latch_out),
    .latch_enable_out(sw_444_latch_out),
    .scan_select_in(sw_443_scan_out),
    .scan_select_out(sw_444_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_444_module_data_in[7] ,
    \sw_444_module_data_in[6] ,
    \sw_444_module_data_in[5] ,
    \sw_444_module_data_in[4] ,
    \sw_444_module_data_in[3] ,
    \sw_444_module_data_in[2] ,
    \sw_444_module_data_in[1] ,
    \sw_444_module_data_in[0] }),
    .module_data_out({\sw_444_module_data_out[7] ,
    \sw_444_module_data_out[6] ,
    \sw_444_module_data_out[5] ,
    \sw_444_module_data_out[4] ,
    \sw_444_module_data_out[3] ,
    \sw_444_module_data_out[2] ,
    \sw_444_module_data_out[1] ,
    \sw_444_module_data_out[0] }));
 scanchain scanchain_445 (.clk_in(sw_444_clk_out),
    .clk_out(sw_445_clk_out),
    .data_in(sw_444_data_out),
    .data_out(sw_445_data_out),
    .latch_enable_in(sw_444_latch_out),
    .latch_enable_out(sw_445_latch_out),
    .scan_select_in(sw_444_scan_out),
    .scan_select_out(sw_445_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_445_module_data_in[7] ,
    \sw_445_module_data_in[6] ,
    \sw_445_module_data_in[5] ,
    \sw_445_module_data_in[4] ,
    \sw_445_module_data_in[3] ,
    \sw_445_module_data_in[2] ,
    \sw_445_module_data_in[1] ,
    \sw_445_module_data_in[0] }),
    .module_data_out({\sw_445_module_data_out[7] ,
    \sw_445_module_data_out[6] ,
    \sw_445_module_data_out[5] ,
    \sw_445_module_data_out[4] ,
    \sw_445_module_data_out[3] ,
    \sw_445_module_data_out[2] ,
    \sw_445_module_data_out[1] ,
    \sw_445_module_data_out[0] }));
 scanchain scanchain_446 (.clk_in(sw_445_clk_out),
    .clk_out(sw_446_clk_out),
    .data_in(sw_445_data_out),
    .data_out(sw_446_data_out),
    .latch_enable_in(sw_445_latch_out),
    .latch_enable_out(sw_446_latch_out),
    .scan_select_in(sw_445_scan_out),
    .scan_select_out(sw_446_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_446_module_data_in[7] ,
    \sw_446_module_data_in[6] ,
    \sw_446_module_data_in[5] ,
    \sw_446_module_data_in[4] ,
    \sw_446_module_data_in[3] ,
    \sw_446_module_data_in[2] ,
    \sw_446_module_data_in[1] ,
    \sw_446_module_data_in[0] }),
    .module_data_out({\sw_446_module_data_out[7] ,
    \sw_446_module_data_out[6] ,
    \sw_446_module_data_out[5] ,
    \sw_446_module_data_out[4] ,
    \sw_446_module_data_out[3] ,
    \sw_446_module_data_out[2] ,
    \sw_446_module_data_out[1] ,
    \sw_446_module_data_out[0] }));
 scanchain scanchain_447 (.clk_in(sw_446_clk_out),
    .clk_out(sw_447_clk_out),
    .data_in(sw_446_data_out),
    .data_out(sw_447_data_out),
    .latch_enable_in(sw_446_latch_out),
    .latch_enable_out(sw_447_latch_out),
    .scan_select_in(sw_446_scan_out),
    .scan_select_out(sw_447_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_447_module_data_in[7] ,
    \sw_447_module_data_in[6] ,
    \sw_447_module_data_in[5] ,
    \sw_447_module_data_in[4] ,
    \sw_447_module_data_in[3] ,
    \sw_447_module_data_in[2] ,
    \sw_447_module_data_in[1] ,
    \sw_447_module_data_in[0] }),
    .module_data_out({\sw_447_module_data_out[7] ,
    \sw_447_module_data_out[6] ,
    \sw_447_module_data_out[5] ,
    \sw_447_module_data_out[4] ,
    \sw_447_module_data_out[3] ,
    \sw_447_module_data_out[2] ,
    \sw_447_module_data_out[1] ,
    \sw_447_module_data_out[0] }));
 scanchain scanchain_448 (.clk_in(sw_447_clk_out),
    .clk_out(sw_448_clk_out),
    .data_in(sw_447_data_out),
    .data_out(sw_448_data_out),
    .latch_enable_in(sw_447_latch_out),
    .latch_enable_out(sw_448_latch_out),
    .scan_select_in(sw_447_scan_out),
    .scan_select_out(sw_448_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_448_module_data_in[7] ,
    \sw_448_module_data_in[6] ,
    \sw_448_module_data_in[5] ,
    \sw_448_module_data_in[4] ,
    \sw_448_module_data_in[3] ,
    \sw_448_module_data_in[2] ,
    \sw_448_module_data_in[1] ,
    \sw_448_module_data_in[0] }),
    .module_data_out({\sw_448_module_data_out[7] ,
    \sw_448_module_data_out[6] ,
    \sw_448_module_data_out[5] ,
    \sw_448_module_data_out[4] ,
    \sw_448_module_data_out[3] ,
    \sw_448_module_data_out[2] ,
    \sw_448_module_data_out[1] ,
    \sw_448_module_data_out[0] }));
 scanchain scanchain_449 (.clk_in(sw_448_clk_out),
    .clk_out(sw_449_clk_out),
    .data_in(sw_448_data_out),
    .data_out(sw_449_data_out),
    .latch_enable_in(sw_448_latch_out),
    .latch_enable_out(sw_449_latch_out),
    .scan_select_in(sw_448_scan_out),
    .scan_select_out(sw_449_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_449_module_data_in[7] ,
    \sw_449_module_data_in[6] ,
    \sw_449_module_data_in[5] ,
    \sw_449_module_data_in[4] ,
    \sw_449_module_data_in[3] ,
    \sw_449_module_data_in[2] ,
    \sw_449_module_data_in[1] ,
    \sw_449_module_data_in[0] }),
    .module_data_out({\sw_449_module_data_out[7] ,
    \sw_449_module_data_out[6] ,
    \sw_449_module_data_out[5] ,
    \sw_449_module_data_out[4] ,
    \sw_449_module_data_out[3] ,
    \sw_449_module_data_out[2] ,
    \sw_449_module_data_out[1] ,
    \sw_449_module_data_out[0] }));
 scanchain scanchain_45 (.clk_in(sw_044_clk_out),
    .clk_out(sw_045_clk_out),
    .data_in(sw_044_data_out),
    .data_out(sw_045_data_out),
    .latch_enable_in(sw_044_latch_out),
    .latch_enable_out(sw_045_latch_out),
    .scan_select_in(sw_044_scan_out),
    .scan_select_out(sw_045_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_045_module_data_in[7] ,
    \sw_045_module_data_in[6] ,
    \sw_045_module_data_in[5] ,
    \sw_045_module_data_in[4] ,
    \sw_045_module_data_in[3] ,
    \sw_045_module_data_in[2] ,
    \sw_045_module_data_in[1] ,
    \sw_045_module_data_in[0] }),
    .module_data_out({\sw_045_module_data_out[7] ,
    \sw_045_module_data_out[6] ,
    \sw_045_module_data_out[5] ,
    \sw_045_module_data_out[4] ,
    \sw_045_module_data_out[3] ,
    \sw_045_module_data_out[2] ,
    \sw_045_module_data_out[1] ,
    \sw_045_module_data_out[0] }));
 scanchain scanchain_450 (.clk_in(sw_449_clk_out),
    .clk_out(sw_450_clk_out),
    .data_in(sw_449_data_out),
    .data_out(sw_450_data_out),
    .latch_enable_in(sw_449_latch_out),
    .latch_enable_out(sw_450_latch_out),
    .scan_select_in(sw_449_scan_out),
    .scan_select_out(sw_450_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_450_module_data_in[7] ,
    \sw_450_module_data_in[6] ,
    \sw_450_module_data_in[5] ,
    \sw_450_module_data_in[4] ,
    \sw_450_module_data_in[3] ,
    \sw_450_module_data_in[2] ,
    \sw_450_module_data_in[1] ,
    \sw_450_module_data_in[0] }),
    .module_data_out({\sw_450_module_data_out[7] ,
    \sw_450_module_data_out[6] ,
    \sw_450_module_data_out[5] ,
    \sw_450_module_data_out[4] ,
    \sw_450_module_data_out[3] ,
    \sw_450_module_data_out[2] ,
    \sw_450_module_data_out[1] ,
    \sw_450_module_data_out[0] }));
 scanchain scanchain_451 (.clk_in(sw_450_clk_out),
    .clk_out(sw_451_clk_out),
    .data_in(sw_450_data_out),
    .data_out(sw_451_data_out),
    .latch_enable_in(sw_450_latch_out),
    .latch_enable_out(sw_451_latch_out),
    .scan_select_in(sw_450_scan_out),
    .scan_select_out(sw_451_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_451_module_data_in[7] ,
    \sw_451_module_data_in[6] ,
    \sw_451_module_data_in[5] ,
    \sw_451_module_data_in[4] ,
    \sw_451_module_data_in[3] ,
    \sw_451_module_data_in[2] ,
    \sw_451_module_data_in[1] ,
    \sw_451_module_data_in[0] }),
    .module_data_out({\sw_451_module_data_out[7] ,
    \sw_451_module_data_out[6] ,
    \sw_451_module_data_out[5] ,
    \sw_451_module_data_out[4] ,
    \sw_451_module_data_out[3] ,
    \sw_451_module_data_out[2] ,
    \sw_451_module_data_out[1] ,
    \sw_451_module_data_out[0] }));
 scanchain scanchain_452 (.clk_in(sw_451_clk_out),
    .clk_out(sw_452_clk_out),
    .data_in(sw_451_data_out),
    .data_out(sw_452_data_out),
    .latch_enable_in(sw_451_latch_out),
    .latch_enable_out(sw_452_latch_out),
    .scan_select_in(sw_451_scan_out),
    .scan_select_out(sw_452_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_452_module_data_in[7] ,
    \sw_452_module_data_in[6] ,
    \sw_452_module_data_in[5] ,
    \sw_452_module_data_in[4] ,
    \sw_452_module_data_in[3] ,
    \sw_452_module_data_in[2] ,
    \sw_452_module_data_in[1] ,
    \sw_452_module_data_in[0] }),
    .module_data_out({\sw_452_module_data_out[7] ,
    \sw_452_module_data_out[6] ,
    \sw_452_module_data_out[5] ,
    \sw_452_module_data_out[4] ,
    \sw_452_module_data_out[3] ,
    \sw_452_module_data_out[2] ,
    \sw_452_module_data_out[1] ,
    \sw_452_module_data_out[0] }));
 scanchain scanchain_453 (.clk_in(sw_452_clk_out),
    .clk_out(sw_453_clk_out),
    .data_in(sw_452_data_out),
    .data_out(sw_453_data_out),
    .latch_enable_in(sw_452_latch_out),
    .latch_enable_out(sw_453_latch_out),
    .scan_select_in(sw_452_scan_out),
    .scan_select_out(sw_453_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_453_module_data_in[7] ,
    \sw_453_module_data_in[6] ,
    \sw_453_module_data_in[5] ,
    \sw_453_module_data_in[4] ,
    \sw_453_module_data_in[3] ,
    \sw_453_module_data_in[2] ,
    \sw_453_module_data_in[1] ,
    \sw_453_module_data_in[0] }),
    .module_data_out({\sw_453_module_data_out[7] ,
    \sw_453_module_data_out[6] ,
    \sw_453_module_data_out[5] ,
    \sw_453_module_data_out[4] ,
    \sw_453_module_data_out[3] ,
    \sw_453_module_data_out[2] ,
    \sw_453_module_data_out[1] ,
    \sw_453_module_data_out[0] }));
 scanchain scanchain_454 (.clk_in(sw_453_clk_out),
    .clk_out(sw_454_clk_out),
    .data_in(sw_453_data_out),
    .data_out(sw_454_data_out),
    .latch_enable_in(sw_453_latch_out),
    .latch_enable_out(sw_454_latch_out),
    .scan_select_in(sw_453_scan_out),
    .scan_select_out(sw_454_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_454_module_data_in[7] ,
    \sw_454_module_data_in[6] ,
    \sw_454_module_data_in[5] ,
    \sw_454_module_data_in[4] ,
    \sw_454_module_data_in[3] ,
    \sw_454_module_data_in[2] ,
    \sw_454_module_data_in[1] ,
    \sw_454_module_data_in[0] }),
    .module_data_out({\sw_454_module_data_out[7] ,
    \sw_454_module_data_out[6] ,
    \sw_454_module_data_out[5] ,
    \sw_454_module_data_out[4] ,
    \sw_454_module_data_out[3] ,
    \sw_454_module_data_out[2] ,
    \sw_454_module_data_out[1] ,
    \sw_454_module_data_out[0] }));
 scanchain scanchain_455 (.clk_in(sw_454_clk_out),
    .clk_out(sw_455_clk_out),
    .data_in(sw_454_data_out),
    .data_out(sw_455_data_out),
    .latch_enable_in(sw_454_latch_out),
    .latch_enable_out(sw_455_latch_out),
    .scan_select_in(sw_454_scan_out),
    .scan_select_out(sw_455_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_455_module_data_in[7] ,
    \sw_455_module_data_in[6] ,
    \sw_455_module_data_in[5] ,
    \sw_455_module_data_in[4] ,
    \sw_455_module_data_in[3] ,
    \sw_455_module_data_in[2] ,
    \sw_455_module_data_in[1] ,
    \sw_455_module_data_in[0] }),
    .module_data_out({\sw_455_module_data_out[7] ,
    \sw_455_module_data_out[6] ,
    \sw_455_module_data_out[5] ,
    \sw_455_module_data_out[4] ,
    \sw_455_module_data_out[3] ,
    \sw_455_module_data_out[2] ,
    \sw_455_module_data_out[1] ,
    \sw_455_module_data_out[0] }));
 scanchain scanchain_456 (.clk_in(sw_455_clk_out),
    .clk_out(sw_456_clk_out),
    .data_in(sw_455_data_out),
    .data_out(sw_456_data_out),
    .latch_enable_in(sw_455_latch_out),
    .latch_enable_out(sw_456_latch_out),
    .scan_select_in(sw_455_scan_out),
    .scan_select_out(sw_456_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_456_module_data_in[7] ,
    \sw_456_module_data_in[6] ,
    \sw_456_module_data_in[5] ,
    \sw_456_module_data_in[4] ,
    \sw_456_module_data_in[3] ,
    \sw_456_module_data_in[2] ,
    \sw_456_module_data_in[1] ,
    \sw_456_module_data_in[0] }),
    .module_data_out({\sw_456_module_data_out[7] ,
    \sw_456_module_data_out[6] ,
    \sw_456_module_data_out[5] ,
    \sw_456_module_data_out[4] ,
    \sw_456_module_data_out[3] ,
    \sw_456_module_data_out[2] ,
    \sw_456_module_data_out[1] ,
    \sw_456_module_data_out[0] }));
 scanchain scanchain_457 (.clk_in(sw_456_clk_out),
    .clk_out(sw_457_clk_out),
    .data_in(sw_456_data_out),
    .data_out(sw_457_data_out),
    .latch_enable_in(sw_456_latch_out),
    .latch_enable_out(sw_457_latch_out),
    .scan_select_in(sw_456_scan_out),
    .scan_select_out(sw_457_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_457_module_data_in[7] ,
    \sw_457_module_data_in[6] ,
    \sw_457_module_data_in[5] ,
    \sw_457_module_data_in[4] ,
    \sw_457_module_data_in[3] ,
    \sw_457_module_data_in[2] ,
    \sw_457_module_data_in[1] ,
    \sw_457_module_data_in[0] }),
    .module_data_out({\sw_457_module_data_out[7] ,
    \sw_457_module_data_out[6] ,
    \sw_457_module_data_out[5] ,
    \sw_457_module_data_out[4] ,
    \sw_457_module_data_out[3] ,
    \sw_457_module_data_out[2] ,
    \sw_457_module_data_out[1] ,
    \sw_457_module_data_out[0] }));
 scanchain scanchain_458 (.clk_in(sw_457_clk_out),
    .clk_out(sw_458_clk_out),
    .data_in(sw_457_data_out),
    .data_out(sw_458_data_out),
    .latch_enable_in(sw_457_latch_out),
    .latch_enable_out(sw_458_latch_out),
    .scan_select_in(sw_457_scan_out),
    .scan_select_out(sw_458_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_458_module_data_in[7] ,
    \sw_458_module_data_in[6] ,
    \sw_458_module_data_in[5] ,
    \sw_458_module_data_in[4] ,
    \sw_458_module_data_in[3] ,
    \sw_458_module_data_in[2] ,
    \sw_458_module_data_in[1] ,
    \sw_458_module_data_in[0] }),
    .module_data_out({\sw_458_module_data_out[7] ,
    \sw_458_module_data_out[6] ,
    \sw_458_module_data_out[5] ,
    \sw_458_module_data_out[4] ,
    \sw_458_module_data_out[3] ,
    \sw_458_module_data_out[2] ,
    \sw_458_module_data_out[1] ,
    \sw_458_module_data_out[0] }));
 scanchain scanchain_459 (.clk_in(sw_458_clk_out),
    .clk_out(sw_459_clk_out),
    .data_in(sw_458_data_out),
    .data_out(sw_459_data_out),
    .latch_enable_in(sw_458_latch_out),
    .latch_enable_out(sw_459_latch_out),
    .scan_select_in(sw_458_scan_out),
    .scan_select_out(sw_459_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_459_module_data_in[7] ,
    \sw_459_module_data_in[6] ,
    \sw_459_module_data_in[5] ,
    \sw_459_module_data_in[4] ,
    \sw_459_module_data_in[3] ,
    \sw_459_module_data_in[2] ,
    \sw_459_module_data_in[1] ,
    \sw_459_module_data_in[0] }),
    .module_data_out({\sw_459_module_data_out[7] ,
    \sw_459_module_data_out[6] ,
    \sw_459_module_data_out[5] ,
    \sw_459_module_data_out[4] ,
    \sw_459_module_data_out[3] ,
    \sw_459_module_data_out[2] ,
    \sw_459_module_data_out[1] ,
    \sw_459_module_data_out[0] }));
 scanchain scanchain_46 (.clk_in(sw_045_clk_out),
    .clk_out(sw_046_clk_out),
    .data_in(sw_045_data_out),
    .data_out(sw_046_data_out),
    .latch_enable_in(sw_045_latch_out),
    .latch_enable_out(sw_046_latch_out),
    .scan_select_in(sw_045_scan_out),
    .scan_select_out(sw_046_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_046_module_data_in[7] ,
    \sw_046_module_data_in[6] ,
    \sw_046_module_data_in[5] ,
    \sw_046_module_data_in[4] ,
    \sw_046_module_data_in[3] ,
    \sw_046_module_data_in[2] ,
    \sw_046_module_data_in[1] ,
    \sw_046_module_data_in[0] }),
    .module_data_out({\sw_046_module_data_out[7] ,
    \sw_046_module_data_out[6] ,
    \sw_046_module_data_out[5] ,
    \sw_046_module_data_out[4] ,
    \sw_046_module_data_out[3] ,
    \sw_046_module_data_out[2] ,
    \sw_046_module_data_out[1] ,
    \sw_046_module_data_out[0] }));
 scanchain scanchain_460 (.clk_in(sw_459_clk_out),
    .clk_out(sw_460_clk_out),
    .data_in(sw_459_data_out),
    .data_out(sw_460_data_out),
    .latch_enable_in(sw_459_latch_out),
    .latch_enable_out(sw_460_latch_out),
    .scan_select_in(sw_459_scan_out),
    .scan_select_out(sw_460_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_460_module_data_in[7] ,
    \sw_460_module_data_in[6] ,
    \sw_460_module_data_in[5] ,
    \sw_460_module_data_in[4] ,
    \sw_460_module_data_in[3] ,
    \sw_460_module_data_in[2] ,
    \sw_460_module_data_in[1] ,
    \sw_460_module_data_in[0] }),
    .module_data_out({\sw_460_module_data_out[7] ,
    \sw_460_module_data_out[6] ,
    \sw_460_module_data_out[5] ,
    \sw_460_module_data_out[4] ,
    \sw_460_module_data_out[3] ,
    \sw_460_module_data_out[2] ,
    \sw_460_module_data_out[1] ,
    \sw_460_module_data_out[0] }));
 scanchain scanchain_461 (.clk_in(sw_460_clk_out),
    .clk_out(sw_461_clk_out),
    .data_in(sw_460_data_out),
    .data_out(sw_461_data_out),
    .latch_enable_in(sw_460_latch_out),
    .latch_enable_out(sw_461_latch_out),
    .scan_select_in(sw_460_scan_out),
    .scan_select_out(sw_461_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_461_module_data_in[7] ,
    \sw_461_module_data_in[6] ,
    \sw_461_module_data_in[5] ,
    \sw_461_module_data_in[4] ,
    \sw_461_module_data_in[3] ,
    \sw_461_module_data_in[2] ,
    \sw_461_module_data_in[1] ,
    \sw_461_module_data_in[0] }),
    .module_data_out({\sw_461_module_data_out[7] ,
    \sw_461_module_data_out[6] ,
    \sw_461_module_data_out[5] ,
    \sw_461_module_data_out[4] ,
    \sw_461_module_data_out[3] ,
    \sw_461_module_data_out[2] ,
    \sw_461_module_data_out[1] ,
    \sw_461_module_data_out[0] }));
 scanchain scanchain_462 (.clk_in(sw_461_clk_out),
    .clk_out(sw_462_clk_out),
    .data_in(sw_461_data_out),
    .data_out(sw_462_data_out),
    .latch_enable_in(sw_461_latch_out),
    .latch_enable_out(sw_462_latch_out),
    .scan_select_in(sw_461_scan_out),
    .scan_select_out(sw_462_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_462_module_data_in[7] ,
    \sw_462_module_data_in[6] ,
    \sw_462_module_data_in[5] ,
    \sw_462_module_data_in[4] ,
    \sw_462_module_data_in[3] ,
    \sw_462_module_data_in[2] ,
    \sw_462_module_data_in[1] ,
    \sw_462_module_data_in[0] }),
    .module_data_out({\sw_462_module_data_out[7] ,
    \sw_462_module_data_out[6] ,
    \sw_462_module_data_out[5] ,
    \sw_462_module_data_out[4] ,
    \sw_462_module_data_out[3] ,
    \sw_462_module_data_out[2] ,
    \sw_462_module_data_out[1] ,
    \sw_462_module_data_out[0] }));
 scanchain scanchain_463 (.clk_in(sw_462_clk_out),
    .clk_out(sw_463_clk_out),
    .data_in(sw_462_data_out),
    .data_out(sw_463_data_out),
    .latch_enable_in(sw_462_latch_out),
    .latch_enable_out(sw_463_latch_out),
    .scan_select_in(sw_462_scan_out),
    .scan_select_out(sw_463_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_463_module_data_in[7] ,
    \sw_463_module_data_in[6] ,
    \sw_463_module_data_in[5] ,
    \sw_463_module_data_in[4] ,
    \sw_463_module_data_in[3] ,
    \sw_463_module_data_in[2] ,
    \sw_463_module_data_in[1] ,
    \sw_463_module_data_in[0] }),
    .module_data_out({\sw_463_module_data_out[7] ,
    \sw_463_module_data_out[6] ,
    \sw_463_module_data_out[5] ,
    \sw_463_module_data_out[4] ,
    \sw_463_module_data_out[3] ,
    \sw_463_module_data_out[2] ,
    \sw_463_module_data_out[1] ,
    \sw_463_module_data_out[0] }));
 scanchain scanchain_464 (.clk_in(sw_463_clk_out),
    .clk_out(sw_464_clk_out),
    .data_in(sw_463_data_out),
    .data_out(sw_464_data_out),
    .latch_enable_in(sw_463_latch_out),
    .latch_enable_out(sw_464_latch_out),
    .scan_select_in(sw_463_scan_out),
    .scan_select_out(sw_464_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_464_module_data_in[7] ,
    \sw_464_module_data_in[6] ,
    \sw_464_module_data_in[5] ,
    \sw_464_module_data_in[4] ,
    \sw_464_module_data_in[3] ,
    \sw_464_module_data_in[2] ,
    \sw_464_module_data_in[1] ,
    \sw_464_module_data_in[0] }),
    .module_data_out({\sw_464_module_data_out[7] ,
    \sw_464_module_data_out[6] ,
    \sw_464_module_data_out[5] ,
    \sw_464_module_data_out[4] ,
    \sw_464_module_data_out[3] ,
    \sw_464_module_data_out[2] ,
    \sw_464_module_data_out[1] ,
    \sw_464_module_data_out[0] }));
 scanchain scanchain_465 (.clk_in(sw_464_clk_out),
    .clk_out(sw_465_clk_out),
    .data_in(sw_464_data_out),
    .data_out(sw_465_data_out),
    .latch_enable_in(sw_464_latch_out),
    .latch_enable_out(sw_465_latch_out),
    .scan_select_in(sw_464_scan_out),
    .scan_select_out(sw_465_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_465_module_data_in[7] ,
    \sw_465_module_data_in[6] ,
    \sw_465_module_data_in[5] ,
    \sw_465_module_data_in[4] ,
    \sw_465_module_data_in[3] ,
    \sw_465_module_data_in[2] ,
    \sw_465_module_data_in[1] ,
    \sw_465_module_data_in[0] }),
    .module_data_out({\sw_465_module_data_out[7] ,
    \sw_465_module_data_out[6] ,
    \sw_465_module_data_out[5] ,
    \sw_465_module_data_out[4] ,
    \sw_465_module_data_out[3] ,
    \sw_465_module_data_out[2] ,
    \sw_465_module_data_out[1] ,
    \sw_465_module_data_out[0] }));
 scanchain scanchain_466 (.clk_in(sw_465_clk_out),
    .clk_out(sw_466_clk_out),
    .data_in(sw_465_data_out),
    .data_out(sw_466_data_out),
    .latch_enable_in(sw_465_latch_out),
    .latch_enable_out(sw_466_latch_out),
    .scan_select_in(sw_465_scan_out),
    .scan_select_out(sw_466_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_466_module_data_in[7] ,
    \sw_466_module_data_in[6] ,
    \sw_466_module_data_in[5] ,
    \sw_466_module_data_in[4] ,
    \sw_466_module_data_in[3] ,
    \sw_466_module_data_in[2] ,
    \sw_466_module_data_in[1] ,
    \sw_466_module_data_in[0] }),
    .module_data_out({\sw_466_module_data_out[7] ,
    \sw_466_module_data_out[6] ,
    \sw_466_module_data_out[5] ,
    \sw_466_module_data_out[4] ,
    \sw_466_module_data_out[3] ,
    \sw_466_module_data_out[2] ,
    \sw_466_module_data_out[1] ,
    \sw_466_module_data_out[0] }));
 scanchain scanchain_467 (.clk_in(sw_466_clk_out),
    .clk_out(sw_467_clk_out),
    .data_in(sw_466_data_out),
    .data_out(sw_467_data_out),
    .latch_enable_in(sw_466_latch_out),
    .latch_enable_out(sw_467_latch_out),
    .scan_select_in(sw_466_scan_out),
    .scan_select_out(sw_467_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_467_module_data_in[7] ,
    \sw_467_module_data_in[6] ,
    \sw_467_module_data_in[5] ,
    \sw_467_module_data_in[4] ,
    \sw_467_module_data_in[3] ,
    \sw_467_module_data_in[2] ,
    \sw_467_module_data_in[1] ,
    \sw_467_module_data_in[0] }),
    .module_data_out({\sw_467_module_data_out[7] ,
    \sw_467_module_data_out[6] ,
    \sw_467_module_data_out[5] ,
    \sw_467_module_data_out[4] ,
    \sw_467_module_data_out[3] ,
    \sw_467_module_data_out[2] ,
    \sw_467_module_data_out[1] ,
    \sw_467_module_data_out[0] }));
 scanchain scanchain_468 (.clk_in(sw_467_clk_out),
    .clk_out(sw_468_clk_out),
    .data_in(sw_467_data_out),
    .data_out(sw_468_data_out),
    .latch_enable_in(sw_467_latch_out),
    .latch_enable_out(sw_468_latch_out),
    .scan_select_in(sw_467_scan_out),
    .scan_select_out(sw_468_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_468_module_data_in[7] ,
    \sw_468_module_data_in[6] ,
    \sw_468_module_data_in[5] ,
    \sw_468_module_data_in[4] ,
    \sw_468_module_data_in[3] ,
    \sw_468_module_data_in[2] ,
    \sw_468_module_data_in[1] ,
    \sw_468_module_data_in[0] }),
    .module_data_out({\sw_468_module_data_out[7] ,
    \sw_468_module_data_out[6] ,
    \sw_468_module_data_out[5] ,
    \sw_468_module_data_out[4] ,
    \sw_468_module_data_out[3] ,
    \sw_468_module_data_out[2] ,
    \sw_468_module_data_out[1] ,
    \sw_468_module_data_out[0] }));
 scanchain scanchain_469 (.clk_in(sw_468_clk_out),
    .clk_out(sw_469_clk_out),
    .data_in(sw_468_data_out),
    .data_out(sw_469_data_out),
    .latch_enable_in(sw_468_latch_out),
    .latch_enable_out(sw_469_latch_out),
    .scan_select_in(sw_468_scan_out),
    .scan_select_out(sw_469_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_469_module_data_in[7] ,
    \sw_469_module_data_in[6] ,
    \sw_469_module_data_in[5] ,
    \sw_469_module_data_in[4] ,
    \sw_469_module_data_in[3] ,
    \sw_469_module_data_in[2] ,
    \sw_469_module_data_in[1] ,
    \sw_469_module_data_in[0] }),
    .module_data_out({\sw_469_module_data_out[7] ,
    \sw_469_module_data_out[6] ,
    \sw_469_module_data_out[5] ,
    \sw_469_module_data_out[4] ,
    \sw_469_module_data_out[3] ,
    \sw_469_module_data_out[2] ,
    \sw_469_module_data_out[1] ,
    \sw_469_module_data_out[0] }));
 scanchain scanchain_47 (.clk_in(sw_046_clk_out),
    .clk_out(sw_047_clk_out),
    .data_in(sw_046_data_out),
    .data_out(sw_047_data_out),
    .latch_enable_in(sw_046_latch_out),
    .latch_enable_out(sw_047_latch_out),
    .scan_select_in(sw_046_scan_out),
    .scan_select_out(sw_047_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_047_module_data_in[7] ,
    \sw_047_module_data_in[6] ,
    \sw_047_module_data_in[5] ,
    \sw_047_module_data_in[4] ,
    \sw_047_module_data_in[3] ,
    \sw_047_module_data_in[2] ,
    \sw_047_module_data_in[1] ,
    \sw_047_module_data_in[0] }),
    .module_data_out({\sw_047_module_data_out[7] ,
    \sw_047_module_data_out[6] ,
    \sw_047_module_data_out[5] ,
    \sw_047_module_data_out[4] ,
    \sw_047_module_data_out[3] ,
    \sw_047_module_data_out[2] ,
    \sw_047_module_data_out[1] ,
    \sw_047_module_data_out[0] }));
 scanchain scanchain_470 (.clk_in(sw_469_clk_out),
    .clk_out(sw_470_clk_out),
    .data_in(sw_469_data_out),
    .data_out(sw_470_data_out),
    .latch_enable_in(sw_469_latch_out),
    .latch_enable_out(sw_470_latch_out),
    .scan_select_in(sw_469_scan_out),
    .scan_select_out(sw_470_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_470_module_data_in[7] ,
    \sw_470_module_data_in[6] ,
    \sw_470_module_data_in[5] ,
    \sw_470_module_data_in[4] ,
    \sw_470_module_data_in[3] ,
    \sw_470_module_data_in[2] ,
    \sw_470_module_data_in[1] ,
    \sw_470_module_data_in[0] }),
    .module_data_out({\sw_470_module_data_out[7] ,
    \sw_470_module_data_out[6] ,
    \sw_470_module_data_out[5] ,
    \sw_470_module_data_out[4] ,
    \sw_470_module_data_out[3] ,
    \sw_470_module_data_out[2] ,
    \sw_470_module_data_out[1] ,
    \sw_470_module_data_out[0] }));
 scanchain scanchain_471 (.clk_in(sw_470_clk_out),
    .clk_out(sw_471_clk_out),
    .data_in(sw_470_data_out),
    .data_out(sw_471_data_out),
    .latch_enable_in(sw_470_latch_out),
    .latch_enable_out(sw_471_latch_out),
    .scan_select_in(sw_470_scan_out),
    .scan_select_out(sw_471_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_471_module_data_in[7] ,
    \sw_471_module_data_in[6] ,
    \sw_471_module_data_in[5] ,
    \sw_471_module_data_in[4] ,
    \sw_471_module_data_in[3] ,
    \sw_471_module_data_in[2] ,
    \sw_471_module_data_in[1] ,
    \sw_471_module_data_in[0] }),
    .module_data_out({\sw_471_module_data_out[7] ,
    \sw_471_module_data_out[6] ,
    \sw_471_module_data_out[5] ,
    \sw_471_module_data_out[4] ,
    \sw_471_module_data_out[3] ,
    \sw_471_module_data_out[2] ,
    \sw_471_module_data_out[1] ,
    \sw_471_module_data_out[0] }));
 scanchain scanchain_472 (.clk_in(sw_471_clk_out),
    .clk_out(sc_clk_in),
    .data_in(sw_471_data_out),
    .data_out(sc_data_in),
    .latch_enable_in(sw_471_latch_out),
    .latch_enable_out(sw_472_latch_out),
    .scan_select_in(sw_471_scan_out),
    .scan_select_out(sw_472_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_472_module_data_in[7] ,
    \sw_472_module_data_in[6] ,
    \sw_472_module_data_in[5] ,
    \sw_472_module_data_in[4] ,
    \sw_472_module_data_in[3] ,
    \sw_472_module_data_in[2] ,
    \sw_472_module_data_in[1] ,
    \sw_472_module_data_in[0] }),
    .module_data_out({\sw_472_module_data_out[7] ,
    \sw_472_module_data_out[6] ,
    \sw_472_module_data_out[5] ,
    \sw_472_module_data_out[4] ,
    \sw_472_module_data_out[3] ,
    \sw_472_module_data_out[2] ,
    \sw_472_module_data_out[1] ,
    \sw_472_module_data_out[0] }));
 scanchain scanchain_48 (.clk_in(sw_047_clk_out),
    .clk_out(sw_048_clk_out),
    .data_in(sw_047_data_out),
    .data_out(sw_048_data_out),
    .latch_enable_in(sw_047_latch_out),
    .latch_enable_out(sw_048_latch_out),
    .scan_select_in(sw_047_scan_out),
    .scan_select_out(sw_048_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_048_module_data_in[7] ,
    \sw_048_module_data_in[6] ,
    \sw_048_module_data_in[5] ,
    \sw_048_module_data_in[4] ,
    \sw_048_module_data_in[3] ,
    \sw_048_module_data_in[2] ,
    \sw_048_module_data_in[1] ,
    \sw_048_module_data_in[0] }),
    .module_data_out({\sw_048_module_data_out[7] ,
    \sw_048_module_data_out[6] ,
    \sw_048_module_data_out[5] ,
    \sw_048_module_data_out[4] ,
    \sw_048_module_data_out[3] ,
    \sw_048_module_data_out[2] ,
    \sw_048_module_data_out[1] ,
    \sw_048_module_data_out[0] }));
 scanchain scanchain_49 (.clk_in(sw_048_clk_out),
    .clk_out(sw_049_clk_out),
    .data_in(sw_048_data_out),
    .data_out(sw_049_data_out),
    .latch_enable_in(sw_048_latch_out),
    .latch_enable_out(sw_049_latch_out),
    .scan_select_in(sw_048_scan_out),
    .scan_select_out(sw_049_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_049_module_data_in[7] ,
    \sw_049_module_data_in[6] ,
    \sw_049_module_data_in[5] ,
    \sw_049_module_data_in[4] ,
    \sw_049_module_data_in[3] ,
    \sw_049_module_data_in[2] ,
    \sw_049_module_data_in[1] ,
    \sw_049_module_data_in[0] }),
    .module_data_out({\sw_049_module_data_out[7] ,
    \sw_049_module_data_out[6] ,
    \sw_049_module_data_out[5] ,
    \sw_049_module_data_out[4] ,
    \sw_049_module_data_out[3] ,
    \sw_049_module_data_out[2] ,
    \sw_049_module_data_out[1] ,
    \sw_049_module_data_out[0] }));
 scanchain scanchain_5 (.clk_in(sw_004_clk_out),
    .clk_out(sw_005_clk_out),
    .data_in(sw_004_data_out),
    .data_out(sw_005_data_out),
    .latch_enable_in(sw_004_latch_out),
    .latch_enable_out(sw_005_latch_out),
    .scan_select_in(sw_004_scan_out),
    .scan_select_out(sw_005_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_005_module_data_in[7] ,
    \sw_005_module_data_in[6] ,
    \sw_005_module_data_in[5] ,
    \sw_005_module_data_in[4] ,
    \sw_005_module_data_in[3] ,
    \sw_005_module_data_in[2] ,
    \sw_005_module_data_in[1] ,
    \sw_005_module_data_in[0] }),
    .module_data_out({\sw_005_module_data_out[7] ,
    \sw_005_module_data_out[6] ,
    \sw_005_module_data_out[5] ,
    \sw_005_module_data_out[4] ,
    \sw_005_module_data_out[3] ,
    \sw_005_module_data_out[2] ,
    \sw_005_module_data_out[1] ,
    \sw_005_module_data_out[0] }));
 scanchain scanchain_50 (.clk_in(sw_049_clk_out),
    .clk_out(sw_050_clk_out),
    .data_in(sw_049_data_out),
    .data_out(sw_050_data_out),
    .latch_enable_in(sw_049_latch_out),
    .latch_enable_out(sw_050_latch_out),
    .scan_select_in(sw_049_scan_out),
    .scan_select_out(sw_050_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_050_module_data_in[7] ,
    \sw_050_module_data_in[6] ,
    \sw_050_module_data_in[5] ,
    \sw_050_module_data_in[4] ,
    \sw_050_module_data_in[3] ,
    \sw_050_module_data_in[2] ,
    \sw_050_module_data_in[1] ,
    \sw_050_module_data_in[0] }),
    .module_data_out({\sw_050_module_data_out[7] ,
    \sw_050_module_data_out[6] ,
    \sw_050_module_data_out[5] ,
    \sw_050_module_data_out[4] ,
    \sw_050_module_data_out[3] ,
    \sw_050_module_data_out[2] ,
    \sw_050_module_data_out[1] ,
    \sw_050_module_data_out[0] }));
 scanchain scanchain_51 (.clk_in(sw_050_clk_out),
    .clk_out(sw_051_clk_out),
    .data_in(sw_050_data_out),
    .data_out(sw_051_data_out),
    .latch_enable_in(sw_050_latch_out),
    .latch_enable_out(sw_051_latch_out),
    .scan_select_in(sw_050_scan_out),
    .scan_select_out(sw_051_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_051_module_data_in[7] ,
    \sw_051_module_data_in[6] ,
    \sw_051_module_data_in[5] ,
    \sw_051_module_data_in[4] ,
    \sw_051_module_data_in[3] ,
    \sw_051_module_data_in[2] ,
    \sw_051_module_data_in[1] ,
    \sw_051_module_data_in[0] }),
    .module_data_out({\sw_051_module_data_out[7] ,
    \sw_051_module_data_out[6] ,
    \sw_051_module_data_out[5] ,
    \sw_051_module_data_out[4] ,
    \sw_051_module_data_out[3] ,
    \sw_051_module_data_out[2] ,
    \sw_051_module_data_out[1] ,
    \sw_051_module_data_out[0] }));
 scanchain scanchain_52 (.clk_in(sw_051_clk_out),
    .clk_out(sw_052_clk_out),
    .data_in(sw_051_data_out),
    .data_out(sw_052_data_out),
    .latch_enable_in(sw_051_latch_out),
    .latch_enable_out(sw_052_latch_out),
    .scan_select_in(sw_051_scan_out),
    .scan_select_out(sw_052_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_052_module_data_in[7] ,
    \sw_052_module_data_in[6] ,
    \sw_052_module_data_in[5] ,
    \sw_052_module_data_in[4] ,
    \sw_052_module_data_in[3] ,
    \sw_052_module_data_in[2] ,
    \sw_052_module_data_in[1] ,
    \sw_052_module_data_in[0] }),
    .module_data_out({\sw_052_module_data_out[7] ,
    \sw_052_module_data_out[6] ,
    \sw_052_module_data_out[5] ,
    \sw_052_module_data_out[4] ,
    \sw_052_module_data_out[3] ,
    \sw_052_module_data_out[2] ,
    \sw_052_module_data_out[1] ,
    \sw_052_module_data_out[0] }));
 scanchain scanchain_53 (.clk_in(sw_052_clk_out),
    .clk_out(sw_053_clk_out),
    .data_in(sw_052_data_out),
    .data_out(sw_053_data_out),
    .latch_enable_in(sw_052_latch_out),
    .latch_enable_out(sw_053_latch_out),
    .scan_select_in(sw_052_scan_out),
    .scan_select_out(sw_053_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_053_module_data_in[7] ,
    \sw_053_module_data_in[6] ,
    \sw_053_module_data_in[5] ,
    \sw_053_module_data_in[4] ,
    \sw_053_module_data_in[3] ,
    \sw_053_module_data_in[2] ,
    \sw_053_module_data_in[1] ,
    \sw_053_module_data_in[0] }),
    .module_data_out({\sw_053_module_data_out[7] ,
    \sw_053_module_data_out[6] ,
    \sw_053_module_data_out[5] ,
    \sw_053_module_data_out[4] ,
    \sw_053_module_data_out[3] ,
    \sw_053_module_data_out[2] ,
    \sw_053_module_data_out[1] ,
    \sw_053_module_data_out[0] }));
 scanchain scanchain_54 (.clk_in(sw_053_clk_out),
    .clk_out(sw_054_clk_out),
    .data_in(sw_053_data_out),
    .data_out(sw_054_data_out),
    .latch_enable_in(sw_053_latch_out),
    .latch_enable_out(sw_054_latch_out),
    .scan_select_in(sw_053_scan_out),
    .scan_select_out(sw_054_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_054_module_data_in[7] ,
    \sw_054_module_data_in[6] ,
    \sw_054_module_data_in[5] ,
    \sw_054_module_data_in[4] ,
    \sw_054_module_data_in[3] ,
    \sw_054_module_data_in[2] ,
    \sw_054_module_data_in[1] ,
    \sw_054_module_data_in[0] }),
    .module_data_out({\sw_054_module_data_out[7] ,
    \sw_054_module_data_out[6] ,
    \sw_054_module_data_out[5] ,
    \sw_054_module_data_out[4] ,
    \sw_054_module_data_out[3] ,
    \sw_054_module_data_out[2] ,
    \sw_054_module_data_out[1] ,
    \sw_054_module_data_out[0] }));
 scanchain scanchain_55 (.clk_in(sw_054_clk_out),
    .clk_out(sw_055_clk_out),
    .data_in(sw_054_data_out),
    .data_out(sw_055_data_out),
    .latch_enable_in(sw_054_latch_out),
    .latch_enable_out(sw_055_latch_out),
    .scan_select_in(sw_054_scan_out),
    .scan_select_out(sw_055_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_055_module_data_in[7] ,
    \sw_055_module_data_in[6] ,
    \sw_055_module_data_in[5] ,
    \sw_055_module_data_in[4] ,
    \sw_055_module_data_in[3] ,
    \sw_055_module_data_in[2] ,
    \sw_055_module_data_in[1] ,
    \sw_055_module_data_in[0] }),
    .module_data_out({\sw_055_module_data_out[7] ,
    \sw_055_module_data_out[6] ,
    \sw_055_module_data_out[5] ,
    \sw_055_module_data_out[4] ,
    \sw_055_module_data_out[3] ,
    \sw_055_module_data_out[2] ,
    \sw_055_module_data_out[1] ,
    \sw_055_module_data_out[0] }));
 scanchain scanchain_56 (.clk_in(sw_055_clk_out),
    .clk_out(sw_056_clk_out),
    .data_in(sw_055_data_out),
    .data_out(sw_056_data_out),
    .latch_enable_in(sw_055_latch_out),
    .latch_enable_out(sw_056_latch_out),
    .scan_select_in(sw_055_scan_out),
    .scan_select_out(sw_056_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_056_module_data_in[7] ,
    \sw_056_module_data_in[6] ,
    \sw_056_module_data_in[5] ,
    \sw_056_module_data_in[4] ,
    \sw_056_module_data_in[3] ,
    \sw_056_module_data_in[2] ,
    \sw_056_module_data_in[1] ,
    \sw_056_module_data_in[0] }),
    .module_data_out({\sw_056_module_data_out[7] ,
    \sw_056_module_data_out[6] ,
    \sw_056_module_data_out[5] ,
    \sw_056_module_data_out[4] ,
    \sw_056_module_data_out[3] ,
    \sw_056_module_data_out[2] ,
    \sw_056_module_data_out[1] ,
    \sw_056_module_data_out[0] }));
 scanchain scanchain_57 (.clk_in(sw_056_clk_out),
    .clk_out(sw_057_clk_out),
    .data_in(sw_056_data_out),
    .data_out(sw_057_data_out),
    .latch_enable_in(sw_056_latch_out),
    .latch_enable_out(sw_057_latch_out),
    .scan_select_in(sw_056_scan_out),
    .scan_select_out(sw_057_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_057_module_data_in[7] ,
    \sw_057_module_data_in[6] ,
    \sw_057_module_data_in[5] ,
    \sw_057_module_data_in[4] ,
    \sw_057_module_data_in[3] ,
    \sw_057_module_data_in[2] ,
    \sw_057_module_data_in[1] ,
    \sw_057_module_data_in[0] }),
    .module_data_out({\sw_057_module_data_out[7] ,
    \sw_057_module_data_out[6] ,
    \sw_057_module_data_out[5] ,
    \sw_057_module_data_out[4] ,
    \sw_057_module_data_out[3] ,
    \sw_057_module_data_out[2] ,
    \sw_057_module_data_out[1] ,
    \sw_057_module_data_out[0] }));
 scanchain scanchain_58 (.clk_in(sw_057_clk_out),
    .clk_out(sw_058_clk_out),
    .data_in(sw_057_data_out),
    .data_out(sw_058_data_out),
    .latch_enable_in(sw_057_latch_out),
    .latch_enable_out(sw_058_latch_out),
    .scan_select_in(sw_057_scan_out),
    .scan_select_out(sw_058_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_058_module_data_in[7] ,
    \sw_058_module_data_in[6] ,
    \sw_058_module_data_in[5] ,
    \sw_058_module_data_in[4] ,
    \sw_058_module_data_in[3] ,
    \sw_058_module_data_in[2] ,
    \sw_058_module_data_in[1] ,
    \sw_058_module_data_in[0] }),
    .module_data_out({\sw_058_module_data_out[7] ,
    \sw_058_module_data_out[6] ,
    \sw_058_module_data_out[5] ,
    \sw_058_module_data_out[4] ,
    \sw_058_module_data_out[3] ,
    \sw_058_module_data_out[2] ,
    \sw_058_module_data_out[1] ,
    \sw_058_module_data_out[0] }));
 scanchain scanchain_59 (.clk_in(sw_058_clk_out),
    .clk_out(sw_059_clk_out),
    .data_in(sw_058_data_out),
    .data_out(sw_059_data_out),
    .latch_enable_in(sw_058_latch_out),
    .latch_enable_out(sw_059_latch_out),
    .scan_select_in(sw_058_scan_out),
    .scan_select_out(sw_059_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_059_module_data_in[7] ,
    \sw_059_module_data_in[6] ,
    \sw_059_module_data_in[5] ,
    \sw_059_module_data_in[4] ,
    \sw_059_module_data_in[3] ,
    \sw_059_module_data_in[2] ,
    \sw_059_module_data_in[1] ,
    \sw_059_module_data_in[0] }),
    .module_data_out({\sw_059_module_data_out[7] ,
    \sw_059_module_data_out[6] ,
    \sw_059_module_data_out[5] ,
    \sw_059_module_data_out[4] ,
    \sw_059_module_data_out[3] ,
    \sw_059_module_data_out[2] ,
    \sw_059_module_data_out[1] ,
    \sw_059_module_data_out[0] }));
 scanchain scanchain_6 (.clk_in(sw_005_clk_out),
    .clk_out(sw_006_clk_out),
    .data_in(sw_005_data_out),
    .data_out(sw_006_data_out),
    .latch_enable_in(sw_005_latch_out),
    .latch_enable_out(sw_006_latch_out),
    .scan_select_in(sw_005_scan_out),
    .scan_select_out(sw_006_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_006_module_data_in[7] ,
    \sw_006_module_data_in[6] ,
    \sw_006_module_data_in[5] ,
    \sw_006_module_data_in[4] ,
    \sw_006_module_data_in[3] ,
    \sw_006_module_data_in[2] ,
    \sw_006_module_data_in[1] ,
    \sw_006_module_data_in[0] }),
    .module_data_out({\sw_006_module_data_out[7] ,
    \sw_006_module_data_out[6] ,
    \sw_006_module_data_out[5] ,
    \sw_006_module_data_out[4] ,
    \sw_006_module_data_out[3] ,
    \sw_006_module_data_out[2] ,
    \sw_006_module_data_out[1] ,
    \sw_006_module_data_out[0] }));
 scanchain scanchain_60 (.clk_in(sw_059_clk_out),
    .clk_out(sw_060_clk_out),
    .data_in(sw_059_data_out),
    .data_out(sw_060_data_out),
    .latch_enable_in(sw_059_latch_out),
    .latch_enable_out(sw_060_latch_out),
    .scan_select_in(sw_059_scan_out),
    .scan_select_out(sw_060_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_060_module_data_in[7] ,
    \sw_060_module_data_in[6] ,
    \sw_060_module_data_in[5] ,
    \sw_060_module_data_in[4] ,
    \sw_060_module_data_in[3] ,
    \sw_060_module_data_in[2] ,
    \sw_060_module_data_in[1] ,
    \sw_060_module_data_in[0] }),
    .module_data_out({\sw_060_module_data_out[7] ,
    \sw_060_module_data_out[6] ,
    \sw_060_module_data_out[5] ,
    \sw_060_module_data_out[4] ,
    \sw_060_module_data_out[3] ,
    \sw_060_module_data_out[2] ,
    \sw_060_module_data_out[1] ,
    \sw_060_module_data_out[0] }));
 scanchain scanchain_61 (.clk_in(sw_060_clk_out),
    .clk_out(sw_061_clk_out),
    .data_in(sw_060_data_out),
    .data_out(sw_061_data_out),
    .latch_enable_in(sw_060_latch_out),
    .latch_enable_out(sw_061_latch_out),
    .scan_select_in(sw_060_scan_out),
    .scan_select_out(sw_061_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_061_module_data_in[7] ,
    \sw_061_module_data_in[6] ,
    \sw_061_module_data_in[5] ,
    \sw_061_module_data_in[4] ,
    \sw_061_module_data_in[3] ,
    \sw_061_module_data_in[2] ,
    \sw_061_module_data_in[1] ,
    \sw_061_module_data_in[0] }),
    .module_data_out({\sw_061_module_data_out[7] ,
    \sw_061_module_data_out[6] ,
    \sw_061_module_data_out[5] ,
    \sw_061_module_data_out[4] ,
    \sw_061_module_data_out[3] ,
    \sw_061_module_data_out[2] ,
    \sw_061_module_data_out[1] ,
    \sw_061_module_data_out[0] }));
 scanchain scanchain_62 (.clk_in(sw_061_clk_out),
    .clk_out(sw_062_clk_out),
    .data_in(sw_061_data_out),
    .data_out(sw_062_data_out),
    .latch_enable_in(sw_061_latch_out),
    .latch_enable_out(sw_062_latch_out),
    .scan_select_in(sw_061_scan_out),
    .scan_select_out(sw_062_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_062_module_data_in[7] ,
    \sw_062_module_data_in[6] ,
    \sw_062_module_data_in[5] ,
    \sw_062_module_data_in[4] ,
    \sw_062_module_data_in[3] ,
    \sw_062_module_data_in[2] ,
    \sw_062_module_data_in[1] ,
    \sw_062_module_data_in[0] }),
    .module_data_out({\sw_062_module_data_out[7] ,
    \sw_062_module_data_out[6] ,
    \sw_062_module_data_out[5] ,
    \sw_062_module_data_out[4] ,
    \sw_062_module_data_out[3] ,
    \sw_062_module_data_out[2] ,
    \sw_062_module_data_out[1] ,
    \sw_062_module_data_out[0] }));
 scanchain scanchain_63 (.clk_in(sw_062_clk_out),
    .clk_out(sw_063_clk_out),
    .data_in(sw_062_data_out),
    .data_out(sw_063_data_out),
    .latch_enable_in(sw_062_latch_out),
    .latch_enable_out(sw_063_latch_out),
    .scan_select_in(sw_062_scan_out),
    .scan_select_out(sw_063_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_063_module_data_in[7] ,
    \sw_063_module_data_in[6] ,
    \sw_063_module_data_in[5] ,
    \sw_063_module_data_in[4] ,
    \sw_063_module_data_in[3] ,
    \sw_063_module_data_in[2] ,
    \sw_063_module_data_in[1] ,
    \sw_063_module_data_in[0] }),
    .module_data_out({\sw_063_module_data_out[7] ,
    \sw_063_module_data_out[6] ,
    \sw_063_module_data_out[5] ,
    \sw_063_module_data_out[4] ,
    \sw_063_module_data_out[3] ,
    \sw_063_module_data_out[2] ,
    \sw_063_module_data_out[1] ,
    \sw_063_module_data_out[0] }));
 scanchain scanchain_64 (.clk_in(sw_063_clk_out),
    .clk_out(sw_064_clk_out),
    .data_in(sw_063_data_out),
    .data_out(sw_064_data_out),
    .latch_enable_in(sw_063_latch_out),
    .latch_enable_out(sw_064_latch_out),
    .scan_select_in(sw_063_scan_out),
    .scan_select_out(sw_064_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_064_module_data_in[7] ,
    \sw_064_module_data_in[6] ,
    \sw_064_module_data_in[5] ,
    \sw_064_module_data_in[4] ,
    \sw_064_module_data_in[3] ,
    \sw_064_module_data_in[2] ,
    \sw_064_module_data_in[1] ,
    \sw_064_module_data_in[0] }),
    .module_data_out({\sw_064_module_data_out[7] ,
    \sw_064_module_data_out[6] ,
    \sw_064_module_data_out[5] ,
    \sw_064_module_data_out[4] ,
    \sw_064_module_data_out[3] ,
    \sw_064_module_data_out[2] ,
    \sw_064_module_data_out[1] ,
    \sw_064_module_data_out[0] }));
 scanchain scanchain_65 (.clk_in(sw_064_clk_out),
    .clk_out(sw_065_clk_out),
    .data_in(sw_064_data_out),
    .data_out(sw_065_data_out),
    .latch_enable_in(sw_064_latch_out),
    .latch_enable_out(sw_065_latch_out),
    .scan_select_in(sw_064_scan_out),
    .scan_select_out(sw_065_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_065_module_data_in[7] ,
    \sw_065_module_data_in[6] ,
    \sw_065_module_data_in[5] ,
    \sw_065_module_data_in[4] ,
    \sw_065_module_data_in[3] ,
    \sw_065_module_data_in[2] ,
    \sw_065_module_data_in[1] ,
    \sw_065_module_data_in[0] }),
    .module_data_out({\sw_065_module_data_out[7] ,
    \sw_065_module_data_out[6] ,
    \sw_065_module_data_out[5] ,
    \sw_065_module_data_out[4] ,
    \sw_065_module_data_out[3] ,
    \sw_065_module_data_out[2] ,
    \sw_065_module_data_out[1] ,
    \sw_065_module_data_out[0] }));
 scanchain scanchain_66 (.clk_in(sw_065_clk_out),
    .clk_out(sw_066_clk_out),
    .data_in(sw_065_data_out),
    .data_out(sw_066_data_out),
    .latch_enable_in(sw_065_latch_out),
    .latch_enable_out(sw_066_latch_out),
    .scan_select_in(sw_065_scan_out),
    .scan_select_out(sw_066_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_066_module_data_in[7] ,
    \sw_066_module_data_in[6] ,
    \sw_066_module_data_in[5] ,
    \sw_066_module_data_in[4] ,
    \sw_066_module_data_in[3] ,
    \sw_066_module_data_in[2] ,
    \sw_066_module_data_in[1] ,
    \sw_066_module_data_in[0] }),
    .module_data_out({\sw_066_module_data_out[7] ,
    \sw_066_module_data_out[6] ,
    \sw_066_module_data_out[5] ,
    \sw_066_module_data_out[4] ,
    \sw_066_module_data_out[3] ,
    \sw_066_module_data_out[2] ,
    \sw_066_module_data_out[1] ,
    \sw_066_module_data_out[0] }));
 scanchain scanchain_67 (.clk_in(sw_066_clk_out),
    .clk_out(sw_067_clk_out),
    .data_in(sw_066_data_out),
    .data_out(sw_067_data_out),
    .latch_enable_in(sw_066_latch_out),
    .latch_enable_out(sw_067_latch_out),
    .scan_select_in(sw_066_scan_out),
    .scan_select_out(sw_067_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_067_module_data_in[7] ,
    \sw_067_module_data_in[6] ,
    \sw_067_module_data_in[5] ,
    \sw_067_module_data_in[4] ,
    \sw_067_module_data_in[3] ,
    \sw_067_module_data_in[2] ,
    \sw_067_module_data_in[1] ,
    \sw_067_module_data_in[0] }),
    .module_data_out({\sw_067_module_data_out[7] ,
    \sw_067_module_data_out[6] ,
    \sw_067_module_data_out[5] ,
    \sw_067_module_data_out[4] ,
    \sw_067_module_data_out[3] ,
    \sw_067_module_data_out[2] ,
    \sw_067_module_data_out[1] ,
    \sw_067_module_data_out[0] }));
 scanchain scanchain_68 (.clk_in(sw_067_clk_out),
    .clk_out(sw_068_clk_out),
    .data_in(sw_067_data_out),
    .data_out(sw_068_data_out),
    .latch_enable_in(sw_067_latch_out),
    .latch_enable_out(sw_068_latch_out),
    .scan_select_in(sw_067_scan_out),
    .scan_select_out(sw_068_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_068_module_data_in[7] ,
    \sw_068_module_data_in[6] ,
    \sw_068_module_data_in[5] ,
    \sw_068_module_data_in[4] ,
    \sw_068_module_data_in[3] ,
    \sw_068_module_data_in[2] ,
    \sw_068_module_data_in[1] ,
    \sw_068_module_data_in[0] }),
    .module_data_out({\sw_068_module_data_out[7] ,
    \sw_068_module_data_out[6] ,
    \sw_068_module_data_out[5] ,
    \sw_068_module_data_out[4] ,
    \sw_068_module_data_out[3] ,
    \sw_068_module_data_out[2] ,
    \sw_068_module_data_out[1] ,
    \sw_068_module_data_out[0] }));
 scanchain scanchain_69 (.clk_in(sw_068_clk_out),
    .clk_out(sw_069_clk_out),
    .data_in(sw_068_data_out),
    .data_out(sw_069_data_out),
    .latch_enable_in(sw_068_latch_out),
    .latch_enable_out(sw_069_latch_out),
    .scan_select_in(sw_068_scan_out),
    .scan_select_out(sw_069_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_069_module_data_in[7] ,
    \sw_069_module_data_in[6] ,
    \sw_069_module_data_in[5] ,
    \sw_069_module_data_in[4] ,
    \sw_069_module_data_in[3] ,
    \sw_069_module_data_in[2] ,
    \sw_069_module_data_in[1] ,
    \sw_069_module_data_in[0] }),
    .module_data_out({\sw_069_module_data_out[7] ,
    \sw_069_module_data_out[6] ,
    \sw_069_module_data_out[5] ,
    \sw_069_module_data_out[4] ,
    \sw_069_module_data_out[3] ,
    \sw_069_module_data_out[2] ,
    \sw_069_module_data_out[1] ,
    \sw_069_module_data_out[0] }));
 scanchain scanchain_7 (.clk_in(sw_006_clk_out),
    .clk_out(sw_007_clk_out),
    .data_in(sw_006_data_out),
    .data_out(sw_007_data_out),
    .latch_enable_in(sw_006_latch_out),
    .latch_enable_out(sw_007_latch_out),
    .scan_select_in(sw_006_scan_out),
    .scan_select_out(sw_007_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_007_module_data_in[7] ,
    \sw_007_module_data_in[6] ,
    \sw_007_module_data_in[5] ,
    \sw_007_module_data_in[4] ,
    \sw_007_module_data_in[3] ,
    \sw_007_module_data_in[2] ,
    \sw_007_module_data_in[1] ,
    \sw_007_module_data_in[0] }),
    .module_data_out({\sw_007_module_data_out[7] ,
    \sw_007_module_data_out[6] ,
    \sw_007_module_data_out[5] ,
    \sw_007_module_data_out[4] ,
    \sw_007_module_data_out[3] ,
    \sw_007_module_data_out[2] ,
    \sw_007_module_data_out[1] ,
    \sw_007_module_data_out[0] }));
 scanchain scanchain_70 (.clk_in(sw_069_clk_out),
    .clk_out(sw_070_clk_out),
    .data_in(sw_069_data_out),
    .data_out(sw_070_data_out),
    .latch_enable_in(sw_069_latch_out),
    .latch_enable_out(sw_070_latch_out),
    .scan_select_in(sw_069_scan_out),
    .scan_select_out(sw_070_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_070_module_data_in[7] ,
    \sw_070_module_data_in[6] ,
    \sw_070_module_data_in[5] ,
    \sw_070_module_data_in[4] ,
    \sw_070_module_data_in[3] ,
    \sw_070_module_data_in[2] ,
    \sw_070_module_data_in[1] ,
    \sw_070_module_data_in[0] }),
    .module_data_out({\sw_070_module_data_out[7] ,
    \sw_070_module_data_out[6] ,
    \sw_070_module_data_out[5] ,
    \sw_070_module_data_out[4] ,
    \sw_070_module_data_out[3] ,
    \sw_070_module_data_out[2] ,
    \sw_070_module_data_out[1] ,
    \sw_070_module_data_out[0] }));
 scanchain scanchain_71 (.clk_in(sw_070_clk_out),
    .clk_out(sw_071_clk_out),
    .data_in(sw_070_data_out),
    .data_out(sw_071_data_out),
    .latch_enable_in(sw_070_latch_out),
    .latch_enable_out(sw_071_latch_out),
    .scan_select_in(sw_070_scan_out),
    .scan_select_out(sw_071_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_071_module_data_in[7] ,
    \sw_071_module_data_in[6] ,
    \sw_071_module_data_in[5] ,
    \sw_071_module_data_in[4] ,
    \sw_071_module_data_in[3] ,
    \sw_071_module_data_in[2] ,
    \sw_071_module_data_in[1] ,
    \sw_071_module_data_in[0] }),
    .module_data_out({\sw_071_module_data_out[7] ,
    \sw_071_module_data_out[6] ,
    \sw_071_module_data_out[5] ,
    \sw_071_module_data_out[4] ,
    \sw_071_module_data_out[3] ,
    \sw_071_module_data_out[2] ,
    \sw_071_module_data_out[1] ,
    \sw_071_module_data_out[0] }));
 scanchain scanchain_72 (.clk_in(sw_071_clk_out),
    .clk_out(sw_072_clk_out),
    .data_in(sw_071_data_out),
    .data_out(sw_072_data_out),
    .latch_enable_in(sw_071_latch_out),
    .latch_enable_out(sw_072_latch_out),
    .scan_select_in(sw_071_scan_out),
    .scan_select_out(sw_072_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_072_module_data_in[7] ,
    \sw_072_module_data_in[6] ,
    \sw_072_module_data_in[5] ,
    \sw_072_module_data_in[4] ,
    \sw_072_module_data_in[3] ,
    \sw_072_module_data_in[2] ,
    \sw_072_module_data_in[1] ,
    \sw_072_module_data_in[0] }),
    .module_data_out({\sw_072_module_data_out[7] ,
    \sw_072_module_data_out[6] ,
    \sw_072_module_data_out[5] ,
    \sw_072_module_data_out[4] ,
    \sw_072_module_data_out[3] ,
    \sw_072_module_data_out[2] ,
    \sw_072_module_data_out[1] ,
    \sw_072_module_data_out[0] }));
 scanchain scanchain_73 (.clk_in(sw_072_clk_out),
    .clk_out(sw_073_clk_out),
    .data_in(sw_072_data_out),
    .data_out(sw_073_data_out),
    .latch_enable_in(sw_072_latch_out),
    .latch_enable_out(sw_073_latch_out),
    .scan_select_in(sw_072_scan_out),
    .scan_select_out(sw_073_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_073_module_data_in[7] ,
    \sw_073_module_data_in[6] ,
    \sw_073_module_data_in[5] ,
    \sw_073_module_data_in[4] ,
    \sw_073_module_data_in[3] ,
    \sw_073_module_data_in[2] ,
    \sw_073_module_data_in[1] ,
    \sw_073_module_data_in[0] }),
    .module_data_out({\sw_073_module_data_out[7] ,
    \sw_073_module_data_out[6] ,
    \sw_073_module_data_out[5] ,
    \sw_073_module_data_out[4] ,
    \sw_073_module_data_out[3] ,
    \sw_073_module_data_out[2] ,
    \sw_073_module_data_out[1] ,
    \sw_073_module_data_out[0] }));
 scanchain scanchain_74 (.clk_in(sw_073_clk_out),
    .clk_out(sw_074_clk_out),
    .data_in(sw_073_data_out),
    .data_out(sw_074_data_out),
    .latch_enable_in(sw_073_latch_out),
    .latch_enable_out(sw_074_latch_out),
    .scan_select_in(sw_073_scan_out),
    .scan_select_out(sw_074_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_074_module_data_in[7] ,
    \sw_074_module_data_in[6] ,
    \sw_074_module_data_in[5] ,
    \sw_074_module_data_in[4] ,
    \sw_074_module_data_in[3] ,
    \sw_074_module_data_in[2] ,
    \sw_074_module_data_in[1] ,
    \sw_074_module_data_in[0] }),
    .module_data_out({\sw_074_module_data_out[7] ,
    \sw_074_module_data_out[6] ,
    \sw_074_module_data_out[5] ,
    \sw_074_module_data_out[4] ,
    \sw_074_module_data_out[3] ,
    \sw_074_module_data_out[2] ,
    \sw_074_module_data_out[1] ,
    \sw_074_module_data_out[0] }));
 scanchain scanchain_75 (.clk_in(sw_074_clk_out),
    .clk_out(sw_075_clk_out),
    .data_in(sw_074_data_out),
    .data_out(sw_075_data_out),
    .latch_enable_in(sw_074_latch_out),
    .latch_enable_out(sw_075_latch_out),
    .scan_select_in(sw_074_scan_out),
    .scan_select_out(sw_075_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_075_module_data_in[7] ,
    \sw_075_module_data_in[6] ,
    \sw_075_module_data_in[5] ,
    \sw_075_module_data_in[4] ,
    \sw_075_module_data_in[3] ,
    \sw_075_module_data_in[2] ,
    \sw_075_module_data_in[1] ,
    \sw_075_module_data_in[0] }),
    .module_data_out({\sw_075_module_data_out[7] ,
    \sw_075_module_data_out[6] ,
    \sw_075_module_data_out[5] ,
    \sw_075_module_data_out[4] ,
    \sw_075_module_data_out[3] ,
    \sw_075_module_data_out[2] ,
    \sw_075_module_data_out[1] ,
    \sw_075_module_data_out[0] }));
 scanchain scanchain_76 (.clk_in(sw_075_clk_out),
    .clk_out(sw_076_clk_out),
    .data_in(sw_075_data_out),
    .data_out(sw_076_data_out),
    .latch_enable_in(sw_075_latch_out),
    .latch_enable_out(sw_076_latch_out),
    .scan_select_in(sw_075_scan_out),
    .scan_select_out(sw_076_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_076_module_data_in[7] ,
    \sw_076_module_data_in[6] ,
    \sw_076_module_data_in[5] ,
    \sw_076_module_data_in[4] ,
    \sw_076_module_data_in[3] ,
    \sw_076_module_data_in[2] ,
    \sw_076_module_data_in[1] ,
    \sw_076_module_data_in[0] }),
    .module_data_out({\sw_076_module_data_out[7] ,
    \sw_076_module_data_out[6] ,
    \sw_076_module_data_out[5] ,
    \sw_076_module_data_out[4] ,
    \sw_076_module_data_out[3] ,
    \sw_076_module_data_out[2] ,
    \sw_076_module_data_out[1] ,
    \sw_076_module_data_out[0] }));
 scanchain scanchain_77 (.clk_in(sw_076_clk_out),
    .clk_out(sw_077_clk_out),
    .data_in(sw_076_data_out),
    .data_out(sw_077_data_out),
    .latch_enable_in(sw_076_latch_out),
    .latch_enable_out(sw_077_latch_out),
    .scan_select_in(sw_076_scan_out),
    .scan_select_out(sw_077_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_077_module_data_in[7] ,
    \sw_077_module_data_in[6] ,
    \sw_077_module_data_in[5] ,
    \sw_077_module_data_in[4] ,
    \sw_077_module_data_in[3] ,
    \sw_077_module_data_in[2] ,
    \sw_077_module_data_in[1] ,
    \sw_077_module_data_in[0] }),
    .module_data_out({\sw_077_module_data_out[7] ,
    \sw_077_module_data_out[6] ,
    \sw_077_module_data_out[5] ,
    \sw_077_module_data_out[4] ,
    \sw_077_module_data_out[3] ,
    \sw_077_module_data_out[2] ,
    \sw_077_module_data_out[1] ,
    \sw_077_module_data_out[0] }));
 scanchain scanchain_78 (.clk_in(sw_077_clk_out),
    .clk_out(sw_078_clk_out),
    .data_in(sw_077_data_out),
    .data_out(sw_078_data_out),
    .latch_enable_in(sw_077_latch_out),
    .latch_enable_out(sw_078_latch_out),
    .scan_select_in(sw_077_scan_out),
    .scan_select_out(sw_078_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_078_module_data_in[7] ,
    \sw_078_module_data_in[6] ,
    \sw_078_module_data_in[5] ,
    \sw_078_module_data_in[4] ,
    \sw_078_module_data_in[3] ,
    \sw_078_module_data_in[2] ,
    \sw_078_module_data_in[1] ,
    \sw_078_module_data_in[0] }),
    .module_data_out({\sw_078_module_data_out[7] ,
    \sw_078_module_data_out[6] ,
    \sw_078_module_data_out[5] ,
    \sw_078_module_data_out[4] ,
    \sw_078_module_data_out[3] ,
    \sw_078_module_data_out[2] ,
    \sw_078_module_data_out[1] ,
    \sw_078_module_data_out[0] }));
 scanchain scanchain_79 (.clk_in(sw_078_clk_out),
    .clk_out(sw_079_clk_out),
    .data_in(sw_078_data_out),
    .data_out(sw_079_data_out),
    .latch_enable_in(sw_078_latch_out),
    .latch_enable_out(sw_079_latch_out),
    .scan_select_in(sw_078_scan_out),
    .scan_select_out(sw_079_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_079_module_data_in[7] ,
    \sw_079_module_data_in[6] ,
    \sw_079_module_data_in[5] ,
    \sw_079_module_data_in[4] ,
    \sw_079_module_data_in[3] ,
    \sw_079_module_data_in[2] ,
    \sw_079_module_data_in[1] ,
    \sw_079_module_data_in[0] }),
    .module_data_out({\sw_079_module_data_out[7] ,
    \sw_079_module_data_out[6] ,
    \sw_079_module_data_out[5] ,
    \sw_079_module_data_out[4] ,
    \sw_079_module_data_out[3] ,
    \sw_079_module_data_out[2] ,
    \sw_079_module_data_out[1] ,
    \sw_079_module_data_out[0] }));
 scanchain scanchain_8 (.clk_in(sw_007_clk_out),
    .clk_out(sw_008_clk_out),
    .data_in(sw_007_data_out),
    .data_out(sw_008_data_out),
    .latch_enable_in(sw_007_latch_out),
    .latch_enable_out(sw_008_latch_out),
    .scan_select_in(sw_007_scan_out),
    .scan_select_out(sw_008_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_008_module_data_in[7] ,
    \sw_008_module_data_in[6] ,
    \sw_008_module_data_in[5] ,
    \sw_008_module_data_in[4] ,
    \sw_008_module_data_in[3] ,
    \sw_008_module_data_in[2] ,
    \sw_008_module_data_in[1] ,
    \sw_008_module_data_in[0] }),
    .module_data_out({\sw_008_module_data_out[7] ,
    \sw_008_module_data_out[6] ,
    \sw_008_module_data_out[5] ,
    \sw_008_module_data_out[4] ,
    \sw_008_module_data_out[3] ,
    \sw_008_module_data_out[2] ,
    \sw_008_module_data_out[1] ,
    \sw_008_module_data_out[0] }));
 scanchain scanchain_80 (.clk_in(sw_079_clk_out),
    .clk_out(sw_080_clk_out),
    .data_in(sw_079_data_out),
    .data_out(sw_080_data_out),
    .latch_enable_in(sw_079_latch_out),
    .latch_enable_out(sw_080_latch_out),
    .scan_select_in(sw_079_scan_out),
    .scan_select_out(sw_080_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_080_module_data_in[7] ,
    \sw_080_module_data_in[6] ,
    \sw_080_module_data_in[5] ,
    \sw_080_module_data_in[4] ,
    \sw_080_module_data_in[3] ,
    \sw_080_module_data_in[2] ,
    \sw_080_module_data_in[1] ,
    \sw_080_module_data_in[0] }),
    .module_data_out({\sw_080_module_data_out[7] ,
    \sw_080_module_data_out[6] ,
    \sw_080_module_data_out[5] ,
    \sw_080_module_data_out[4] ,
    \sw_080_module_data_out[3] ,
    \sw_080_module_data_out[2] ,
    \sw_080_module_data_out[1] ,
    \sw_080_module_data_out[0] }));
 scanchain scanchain_81 (.clk_in(sw_080_clk_out),
    .clk_out(sw_081_clk_out),
    .data_in(sw_080_data_out),
    .data_out(sw_081_data_out),
    .latch_enable_in(sw_080_latch_out),
    .latch_enable_out(sw_081_latch_out),
    .scan_select_in(sw_080_scan_out),
    .scan_select_out(sw_081_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_081_module_data_in[7] ,
    \sw_081_module_data_in[6] ,
    \sw_081_module_data_in[5] ,
    \sw_081_module_data_in[4] ,
    \sw_081_module_data_in[3] ,
    \sw_081_module_data_in[2] ,
    \sw_081_module_data_in[1] ,
    \sw_081_module_data_in[0] }),
    .module_data_out({\sw_081_module_data_out[7] ,
    \sw_081_module_data_out[6] ,
    \sw_081_module_data_out[5] ,
    \sw_081_module_data_out[4] ,
    \sw_081_module_data_out[3] ,
    \sw_081_module_data_out[2] ,
    \sw_081_module_data_out[1] ,
    \sw_081_module_data_out[0] }));
 scanchain scanchain_82 (.clk_in(sw_081_clk_out),
    .clk_out(sw_082_clk_out),
    .data_in(sw_081_data_out),
    .data_out(sw_082_data_out),
    .latch_enable_in(sw_081_latch_out),
    .latch_enable_out(sw_082_latch_out),
    .scan_select_in(sw_081_scan_out),
    .scan_select_out(sw_082_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_082_module_data_in[7] ,
    \sw_082_module_data_in[6] ,
    \sw_082_module_data_in[5] ,
    \sw_082_module_data_in[4] ,
    \sw_082_module_data_in[3] ,
    \sw_082_module_data_in[2] ,
    \sw_082_module_data_in[1] ,
    \sw_082_module_data_in[0] }),
    .module_data_out({\sw_082_module_data_out[7] ,
    \sw_082_module_data_out[6] ,
    \sw_082_module_data_out[5] ,
    \sw_082_module_data_out[4] ,
    \sw_082_module_data_out[3] ,
    \sw_082_module_data_out[2] ,
    \sw_082_module_data_out[1] ,
    \sw_082_module_data_out[0] }));
 scanchain scanchain_83 (.clk_in(sw_082_clk_out),
    .clk_out(sw_083_clk_out),
    .data_in(sw_082_data_out),
    .data_out(sw_083_data_out),
    .latch_enable_in(sw_082_latch_out),
    .latch_enable_out(sw_083_latch_out),
    .scan_select_in(sw_082_scan_out),
    .scan_select_out(sw_083_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_083_module_data_in[7] ,
    \sw_083_module_data_in[6] ,
    \sw_083_module_data_in[5] ,
    \sw_083_module_data_in[4] ,
    \sw_083_module_data_in[3] ,
    \sw_083_module_data_in[2] ,
    \sw_083_module_data_in[1] ,
    \sw_083_module_data_in[0] }),
    .module_data_out({\sw_083_module_data_out[7] ,
    \sw_083_module_data_out[6] ,
    \sw_083_module_data_out[5] ,
    \sw_083_module_data_out[4] ,
    \sw_083_module_data_out[3] ,
    \sw_083_module_data_out[2] ,
    \sw_083_module_data_out[1] ,
    \sw_083_module_data_out[0] }));
 scanchain scanchain_84 (.clk_in(sw_083_clk_out),
    .clk_out(sw_084_clk_out),
    .data_in(sw_083_data_out),
    .data_out(sw_084_data_out),
    .latch_enable_in(sw_083_latch_out),
    .latch_enable_out(sw_084_latch_out),
    .scan_select_in(sw_083_scan_out),
    .scan_select_out(sw_084_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_084_module_data_in[7] ,
    \sw_084_module_data_in[6] ,
    \sw_084_module_data_in[5] ,
    \sw_084_module_data_in[4] ,
    \sw_084_module_data_in[3] ,
    \sw_084_module_data_in[2] ,
    \sw_084_module_data_in[1] ,
    \sw_084_module_data_in[0] }),
    .module_data_out({\sw_084_module_data_out[7] ,
    \sw_084_module_data_out[6] ,
    \sw_084_module_data_out[5] ,
    \sw_084_module_data_out[4] ,
    \sw_084_module_data_out[3] ,
    \sw_084_module_data_out[2] ,
    \sw_084_module_data_out[1] ,
    \sw_084_module_data_out[0] }));
 scanchain scanchain_85 (.clk_in(sw_084_clk_out),
    .clk_out(sw_085_clk_out),
    .data_in(sw_084_data_out),
    .data_out(sw_085_data_out),
    .latch_enable_in(sw_084_latch_out),
    .latch_enable_out(sw_085_latch_out),
    .scan_select_in(sw_084_scan_out),
    .scan_select_out(sw_085_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_085_module_data_in[7] ,
    \sw_085_module_data_in[6] ,
    \sw_085_module_data_in[5] ,
    \sw_085_module_data_in[4] ,
    \sw_085_module_data_in[3] ,
    \sw_085_module_data_in[2] ,
    \sw_085_module_data_in[1] ,
    \sw_085_module_data_in[0] }),
    .module_data_out({\sw_085_module_data_out[7] ,
    \sw_085_module_data_out[6] ,
    \sw_085_module_data_out[5] ,
    \sw_085_module_data_out[4] ,
    \sw_085_module_data_out[3] ,
    \sw_085_module_data_out[2] ,
    \sw_085_module_data_out[1] ,
    \sw_085_module_data_out[0] }));
 scanchain scanchain_86 (.clk_in(sw_085_clk_out),
    .clk_out(sw_086_clk_out),
    .data_in(sw_085_data_out),
    .data_out(sw_086_data_out),
    .latch_enable_in(sw_085_latch_out),
    .latch_enable_out(sw_086_latch_out),
    .scan_select_in(sw_085_scan_out),
    .scan_select_out(sw_086_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_086_module_data_in[7] ,
    \sw_086_module_data_in[6] ,
    \sw_086_module_data_in[5] ,
    \sw_086_module_data_in[4] ,
    \sw_086_module_data_in[3] ,
    \sw_086_module_data_in[2] ,
    \sw_086_module_data_in[1] ,
    \sw_086_module_data_in[0] }),
    .module_data_out({\sw_086_module_data_out[7] ,
    \sw_086_module_data_out[6] ,
    \sw_086_module_data_out[5] ,
    \sw_086_module_data_out[4] ,
    \sw_086_module_data_out[3] ,
    \sw_086_module_data_out[2] ,
    \sw_086_module_data_out[1] ,
    \sw_086_module_data_out[0] }));
 scanchain scanchain_87 (.clk_in(sw_086_clk_out),
    .clk_out(sw_087_clk_out),
    .data_in(sw_086_data_out),
    .data_out(sw_087_data_out),
    .latch_enable_in(sw_086_latch_out),
    .latch_enable_out(sw_087_latch_out),
    .scan_select_in(sw_086_scan_out),
    .scan_select_out(sw_087_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_087_module_data_in[7] ,
    \sw_087_module_data_in[6] ,
    \sw_087_module_data_in[5] ,
    \sw_087_module_data_in[4] ,
    \sw_087_module_data_in[3] ,
    \sw_087_module_data_in[2] ,
    \sw_087_module_data_in[1] ,
    \sw_087_module_data_in[0] }),
    .module_data_out({\sw_087_module_data_out[7] ,
    \sw_087_module_data_out[6] ,
    \sw_087_module_data_out[5] ,
    \sw_087_module_data_out[4] ,
    \sw_087_module_data_out[3] ,
    \sw_087_module_data_out[2] ,
    \sw_087_module_data_out[1] ,
    \sw_087_module_data_out[0] }));
 scanchain scanchain_88 (.clk_in(sw_087_clk_out),
    .clk_out(sw_088_clk_out),
    .data_in(sw_087_data_out),
    .data_out(sw_088_data_out),
    .latch_enable_in(sw_087_latch_out),
    .latch_enable_out(sw_088_latch_out),
    .scan_select_in(sw_087_scan_out),
    .scan_select_out(sw_088_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_088_module_data_in[7] ,
    \sw_088_module_data_in[6] ,
    \sw_088_module_data_in[5] ,
    \sw_088_module_data_in[4] ,
    \sw_088_module_data_in[3] ,
    \sw_088_module_data_in[2] ,
    \sw_088_module_data_in[1] ,
    \sw_088_module_data_in[0] }),
    .module_data_out({\sw_088_module_data_out[7] ,
    \sw_088_module_data_out[6] ,
    \sw_088_module_data_out[5] ,
    \sw_088_module_data_out[4] ,
    \sw_088_module_data_out[3] ,
    \sw_088_module_data_out[2] ,
    \sw_088_module_data_out[1] ,
    \sw_088_module_data_out[0] }));
 scanchain scanchain_89 (.clk_in(sw_088_clk_out),
    .clk_out(sw_089_clk_out),
    .data_in(sw_088_data_out),
    .data_out(sw_089_data_out),
    .latch_enable_in(sw_088_latch_out),
    .latch_enable_out(sw_089_latch_out),
    .scan_select_in(sw_088_scan_out),
    .scan_select_out(sw_089_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_089_module_data_in[7] ,
    \sw_089_module_data_in[6] ,
    \sw_089_module_data_in[5] ,
    \sw_089_module_data_in[4] ,
    \sw_089_module_data_in[3] ,
    \sw_089_module_data_in[2] ,
    \sw_089_module_data_in[1] ,
    \sw_089_module_data_in[0] }),
    .module_data_out({\sw_089_module_data_out[7] ,
    \sw_089_module_data_out[6] ,
    \sw_089_module_data_out[5] ,
    \sw_089_module_data_out[4] ,
    \sw_089_module_data_out[3] ,
    \sw_089_module_data_out[2] ,
    \sw_089_module_data_out[1] ,
    \sw_089_module_data_out[0] }));
 scanchain scanchain_9 (.clk_in(sw_008_clk_out),
    .clk_out(sw_009_clk_out),
    .data_in(sw_008_data_out),
    .data_out(sw_009_data_out),
    .latch_enable_in(sw_008_latch_out),
    .latch_enable_out(sw_009_latch_out),
    .scan_select_in(sw_008_scan_out),
    .scan_select_out(sw_009_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_009_module_data_in[7] ,
    \sw_009_module_data_in[6] ,
    \sw_009_module_data_in[5] ,
    \sw_009_module_data_in[4] ,
    \sw_009_module_data_in[3] ,
    \sw_009_module_data_in[2] ,
    \sw_009_module_data_in[1] ,
    \sw_009_module_data_in[0] }),
    .module_data_out({\sw_009_module_data_out[7] ,
    \sw_009_module_data_out[6] ,
    \sw_009_module_data_out[5] ,
    \sw_009_module_data_out[4] ,
    \sw_009_module_data_out[3] ,
    \sw_009_module_data_out[2] ,
    \sw_009_module_data_out[1] ,
    \sw_009_module_data_out[0] }));
 scanchain scanchain_90 (.clk_in(sw_089_clk_out),
    .clk_out(sw_090_clk_out),
    .data_in(sw_089_data_out),
    .data_out(sw_090_data_out),
    .latch_enable_in(sw_089_latch_out),
    .latch_enable_out(sw_090_latch_out),
    .scan_select_in(sw_089_scan_out),
    .scan_select_out(sw_090_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_090_module_data_in[7] ,
    \sw_090_module_data_in[6] ,
    \sw_090_module_data_in[5] ,
    \sw_090_module_data_in[4] ,
    \sw_090_module_data_in[3] ,
    \sw_090_module_data_in[2] ,
    \sw_090_module_data_in[1] ,
    \sw_090_module_data_in[0] }),
    .module_data_out({\sw_090_module_data_out[7] ,
    \sw_090_module_data_out[6] ,
    \sw_090_module_data_out[5] ,
    \sw_090_module_data_out[4] ,
    \sw_090_module_data_out[3] ,
    \sw_090_module_data_out[2] ,
    \sw_090_module_data_out[1] ,
    \sw_090_module_data_out[0] }));
 scanchain scanchain_91 (.clk_in(sw_090_clk_out),
    .clk_out(sw_091_clk_out),
    .data_in(sw_090_data_out),
    .data_out(sw_091_data_out),
    .latch_enable_in(sw_090_latch_out),
    .latch_enable_out(sw_091_latch_out),
    .scan_select_in(sw_090_scan_out),
    .scan_select_out(sw_091_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_091_module_data_in[7] ,
    \sw_091_module_data_in[6] ,
    \sw_091_module_data_in[5] ,
    \sw_091_module_data_in[4] ,
    \sw_091_module_data_in[3] ,
    \sw_091_module_data_in[2] ,
    \sw_091_module_data_in[1] ,
    \sw_091_module_data_in[0] }),
    .module_data_out({\sw_091_module_data_out[7] ,
    \sw_091_module_data_out[6] ,
    \sw_091_module_data_out[5] ,
    \sw_091_module_data_out[4] ,
    \sw_091_module_data_out[3] ,
    \sw_091_module_data_out[2] ,
    \sw_091_module_data_out[1] ,
    \sw_091_module_data_out[0] }));
 scanchain scanchain_92 (.clk_in(sw_091_clk_out),
    .clk_out(sw_092_clk_out),
    .data_in(sw_091_data_out),
    .data_out(sw_092_data_out),
    .latch_enable_in(sw_091_latch_out),
    .latch_enable_out(sw_092_latch_out),
    .scan_select_in(sw_091_scan_out),
    .scan_select_out(sw_092_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_092_module_data_in[7] ,
    \sw_092_module_data_in[6] ,
    \sw_092_module_data_in[5] ,
    \sw_092_module_data_in[4] ,
    \sw_092_module_data_in[3] ,
    \sw_092_module_data_in[2] ,
    \sw_092_module_data_in[1] ,
    \sw_092_module_data_in[0] }),
    .module_data_out({\sw_092_module_data_out[7] ,
    \sw_092_module_data_out[6] ,
    \sw_092_module_data_out[5] ,
    \sw_092_module_data_out[4] ,
    \sw_092_module_data_out[3] ,
    \sw_092_module_data_out[2] ,
    \sw_092_module_data_out[1] ,
    \sw_092_module_data_out[0] }));
 scanchain scanchain_93 (.clk_in(sw_092_clk_out),
    .clk_out(sw_093_clk_out),
    .data_in(sw_092_data_out),
    .data_out(sw_093_data_out),
    .latch_enable_in(sw_092_latch_out),
    .latch_enable_out(sw_093_latch_out),
    .scan_select_in(sw_092_scan_out),
    .scan_select_out(sw_093_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_093_module_data_in[7] ,
    \sw_093_module_data_in[6] ,
    \sw_093_module_data_in[5] ,
    \sw_093_module_data_in[4] ,
    \sw_093_module_data_in[3] ,
    \sw_093_module_data_in[2] ,
    \sw_093_module_data_in[1] ,
    \sw_093_module_data_in[0] }),
    .module_data_out({\sw_093_module_data_out[7] ,
    \sw_093_module_data_out[6] ,
    \sw_093_module_data_out[5] ,
    \sw_093_module_data_out[4] ,
    \sw_093_module_data_out[3] ,
    \sw_093_module_data_out[2] ,
    \sw_093_module_data_out[1] ,
    \sw_093_module_data_out[0] }));
 scanchain scanchain_94 (.clk_in(sw_093_clk_out),
    .clk_out(sw_094_clk_out),
    .data_in(sw_093_data_out),
    .data_out(sw_094_data_out),
    .latch_enable_in(sw_093_latch_out),
    .latch_enable_out(sw_094_latch_out),
    .scan_select_in(sw_093_scan_out),
    .scan_select_out(sw_094_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_094_module_data_in[7] ,
    \sw_094_module_data_in[6] ,
    \sw_094_module_data_in[5] ,
    \sw_094_module_data_in[4] ,
    \sw_094_module_data_in[3] ,
    \sw_094_module_data_in[2] ,
    \sw_094_module_data_in[1] ,
    \sw_094_module_data_in[0] }),
    .module_data_out({\sw_094_module_data_out[7] ,
    \sw_094_module_data_out[6] ,
    \sw_094_module_data_out[5] ,
    \sw_094_module_data_out[4] ,
    \sw_094_module_data_out[3] ,
    \sw_094_module_data_out[2] ,
    \sw_094_module_data_out[1] ,
    \sw_094_module_data_out[0] }));
 scanchain scanchain_95 (.clk_in(sw_094_clk_out),
    .clk_out(sw_095_clk_out),
    .data_in(sw_094_data_out),
    .data_out(sw_095_data_out),
    .latch_enable_in(sw_094_latch_out),
    .latch_enable_out(sw_095_latch_out),
    .scan_select_in(sw_094_scan_out),
    .scan_select_out(sw_095_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_095_module_data_in[7] ,
    \sw_095_module_data_in[6] ,
    \sw_095_module_data_in[5] ,
    \sw_095_module_data_in[4] ,
    \sw_095_module_data_in[3] ,
    \sw_095_module_data_in[2] ,
    \sw_095_module_data_in[1] ,
    \sw_095_module_data_in[0] }),
    .module_data_out({\sw_095_module_data_out[7] ,
    \sw_095_module_data_out[6] ,
    \sw_095_module_data_out[5] ,
    \sw_095_module_data_out[4] ,
    \sw_095_module_data_out[3] ,
    \sw_095_module_data_out[2] ,
    \sw_095_module_data_out[1] ,
    \sw_095_module_data_out[0] }));
 scanchain scanchain_96 (.clk_in(sw_095_clk_out),
    .clk_out(sw_096_clk_out),
    .data_in(sw_095_data_out),
    .data_out(sw_096_data_out),
    .latch_enable_in(sw_095_latch_out),
    .latch_enable_out(sw_096_latch_out),
    .scan_select_in(sw_095_scan_out),
    .scan_select_out(sw_096_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_096_module_data_in[7] ,
    \sw_096_module_data_in[6] ,
    \sw_096_module_data_in[5] ,
    \sw_096_module_data_in[4] ,
    \sw_096_module_data_in[3] ,
    \sw_096_module_data_in[2] ,
    \sw_096_module_data_in[1] ,
    \sw_096_module_data_in[0] }),
    .module_data_out({\sw_096_module_data_out[7] ,
    \sw_096_module_data_out[6] ,
    \sw_096_module_data_out[5] ,
    \sw_096_module_data_out[4] ,
    \sw_096_module_data_out[3] ,
    \sw_096_module_data_out[2] ,
    \sw_096_module_data_out[1] ,
    \sw_096_module_data_out[0] }));
 scanchain scanchain_97 (.clk_in(sw_096_clk_out),
    .clk_out(sw_097_clk_out),
    .data_in(sw_096_data_out),
    .data_out(sw_097_data_out),
    .latch_enable_in(sw_096_latch_out),
    .latch_enable_out(sw_097_latch_out),
    .scan_select_in(sw_096_scan_out),
    .scan_select_out(sw_097_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_097_module_data_in[7] ,
    \sw_097_module_data_in[6] ,
    \sw_097_module_data_in[5] ,
    \sw_097_module_data_in[4] ,
    \sw_097_module_data_in[3] ,
    \sw_097_module_data_in[2] ,
    \sw_097_module_data_in[1] ,
    \sw_097_module_data_in[0] }),
    .module_data_out({\sw_097_module_data_out[7] ,
    \sw_097_module_data_out[6] ,
    \sw_097_module_data_out[5] ,
    \sw_097_module_data_out[4] ,
    \sw_097_module_data_out[3] ,
    \sw_097_module_data_out[2] ,
    \sw_097_module_data_out[1] ,
    \sw_097_module_data_out[0] }));
 scanchain scanchain_98 (.clk_in(sw_097_clk_out),
    .clk_out(sw_098_clk_out),
    .data_in(sw_097_data_out),
    .data_out(sw_098_data_out),
    .latch_enable_in(sw_097_latch_out),
    .latch_enable_out(sw_098_latch_out),
    .scan_select_in(sw_097_scan_out),
    .scan_select_out(sw_098_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_098_module_data_in[7] ,
    \sw_098_module_data_in[6] ,
    \sw_098_module_data_in[5] ,
    \sw_098_module_data_in[4] ,
    \sw_098_module_data_in[3] ,
    \sw_098_module_data_in[2] ,
    \sw_098_module_data_in[1] ,
    \sw_098_module_data_in[0] }),
    .module_data_out({\sw_098_module_data_out[7] ,
    \sw_098_module_data_out[6] ,
    \sw_098_module_data_out[5] ,
    \sw_098_module_data_out[4] ,
    \sw_098_module_data_out[3] ,
    \sw_098_module_data_out[2] ,
    \sw_098_module_data_out[1] ,
    \sw_098_module_data_out[0] }));
 scanchain scanchain_99 (.clk_in(sw_098_clk_out),
    .clk_out(sw_099_clk_out),
    .data_in(sw_098_data_out),
    .data_out(sw_099_data_out),
    .latch_enable_in(sw_098_latch_out),
    .latch_enable_out(sw_099_latch_out),
    .scan_select_in(sw_098_scan_out),
    .scan_select_out(sw_099_scan_out),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .module_data_in({\sw_099_module_data_in[7] ,
    \sw_099_module_data_in[6] ,
    \sw_099_module_data_in[5] ,
    \sw_099_module_data_in[4] ,
    \sw_099_module_data_in[3] ,
    \sw_099_module_data_in[2] ,
    \sw_099_module_data_in[1] ,
    \sw_099_module_data_in[0] }),
    .module_data_out({\sw_099_module_data_out[7] ,
    \sw_099_module_data_out[6] ,
    \sw_099_module_data_out[5] ,
    \sw_099_module_data_out[4] ,
    \sw_099_module_data_out[3] ,
    \sw_099_module_data_out[2] ,
    \sw_099_module_data_out[1] ,
    \sw_099_module_data_out[0] }));
 tholin_avalonsemi_5401 tholin_avalonsemi_5401_14 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_014_module_data_in[7] ,
    \sw_014_module_data_in[6] ,
    \sw_014_module_data_in[5] ,
    \sw_014_module_data_in[4] ,
    \sw_014_module_data_in[3] ,
    \sw_014_module_data_in[2] ,
    \sw_014_module_data_in[1] ,
    \sw_014_module_data_in[0] }),
    .io_out({\sw_014_module_data_out[7] ,
    \sw_014_module_data_out[6] ,
    \sw_014_module_data_out[5] ,
    \sw_014_module_data_out[4] ,
    \sw_014_module_data_out[3] ,
    \sw_014_module_data_out[2] ,
    \sw_014_module_data_out[1] ,
    \sw_014_module_data_out[0] }));
 tholin_avalonsemi_tbb1143 tholin_avalonsemi_tbb1143_24 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_024_module_data_in[7] ,
    \sw_024_module_data_in[6] ,
    \sw_024_module_data_in[5] ,
    \sw_024_module_data_in[4] ,
    \sw_024_module_data_in[3] ,
    \sw_024_module_data_in[2] ,
    \sw_024_module_data_in[1] ,
    \sw_024_module_data_in[0] }),
    .io_out({\sw_024_module_data_out[7] ,
    \sw_024_module_data_out[6] ,
    \sw_024_module_data_out[5] ,
    \sw_024_module_data_out[4] ,
    \sw_024_module_data_out[3] ,
    \sw_024_module_data_out[2] ,
    \sw_024_module_data_out[1] ,
    \sw_024_module_data_out[0] }));
 tiny_fft tiny_fft_15 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_015_module_data_in[7] ,
    \sw_015_module_data_in[6] ,
    \sw_015_module_data_in[5] ,
    \sw_015_module_data_in[4] ,
    \sw_015_module_data_in[3] ,
    \sw_015_module_data_in[2] ,
    \sw_015_module_data_in[1] ,
    \sw_015_module_data_in[0] }),
    .io_out({\sw_015_module_data_out[7] ,
    \sw_015_module_data_out[6] ,
    \sw_015_module_data_out[5] ,
    \sw_015_module_data_out[4] ,
    \sw_015_module_data_out[3] ,
    \sw_015_module_data_out[2] ,
    \sw_015_module_data_out[1] ,
    \sw_015_module_data_out[0] }));
 tomkeddie_top_tto tomkeddie_top_tto_2 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_002_module_data_in[7] ,
    \sw_002_module_data_in[6] ,
    \sw_002_module_data_in[5] ,
    \sw_002_module_data_in[4] ,
    \sw_002_module_data_in[3] ,
    \sw_002_module_data_in[2] ,
    \sw_002_module_data_in[1] ,
    \sw_002_module_data_in[0] }),
    .io_out({\sw_002_module_data_out[7] ,
    \sw_002_module_data_out[6] ,
    \sw_002_module_data_out[5] ,
    \sw_002_module_data_out[4] ,
    \sw_002_module_data_out[3] ,
    \sw_002_module_data_out[2] ,
    \sw_002_module_data_out[1] ,
    \sw_002_module_data_out[0] }));
 tomkeddie_top_tto_a tomkeddie_top_tto_a_25 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_025_module_data_in[7] ,
    \sw_025_module_data_in[6] ,
    \sw_025_module_data_in[5] ,
    \sw_025_module_data_in[4] ,
    \sw_025_module_data_in[3] ,
    \sw_025_module_data_in[2] ,
    \sw_025_module_data_in[1] ,
    \sw_025_module_data_in[0] }),
    .io_out({\sw_025_module_data_out[7] ,
    \sw_025_module_data_out[6] ,
    \sw_025_module_data_out[5] ,
    \sw_025_module_data_out[4] ,
    \sw_025_module_data_out[3] ,
    \sw_025_module_data_out[2] ,
    \sw_025_module_data_out[1] ,
    \sw_025_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_0 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_000_module_data_in[7] ,
    \sw_000_module_data_in[6] ,
    \sw_000_module_data_in[5] ,
    \sw_000_module_data_in[4] ,
    \sw_000_module_data_in[3] ,
    \sw_000_module_data_in[2] ,
    \sw_000_module_data_in[1] ,
    \sw_000_module_data_in[0] }),
    .io_out({\sw_000_module_data_out[7] ,
    \sw_000_module_data_out[6] ,
    \sw_000_module_data_out[5] ,
    \sw_000_module_data_out[4] ,
    \sw_000_module_data_out[3] ,
    \sw_000_module_data_out[2] ,
    \sw_000_module_data_out[1] ,
    \sw_000_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_100 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_100_module_data_in[7] ,
    \sw_100_module_data_in[6] ,
    \sw_100_module_data_in[5] ,
    \sw_100_module_data_in[4] ,
    \sw_100_module_data_in[3] ,
    \sw_100_module_data_in[2] ,
    \sw_100_module_data_in[1] ,
    \sw_100_module_data_in[0] }),
    .io_out({\sw_100_module_data_out[7] ,
    \sw_100_module_data_out[6] ,
    \sw_100_module_data_out[5] ,
    \sw_100_module_data_out[4] ,
    \sw_100_module_data_out[3] ,
    \sw_100_module_data_out[2] ,
    \sw_100_module_data_out[1] ,
    \sw_100_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_101 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_101_module_data_in[7] ,
    \sw_101_module_data_in[6] ,
    \sw_101_module_data_in[5] ,
    \sw_101_module_data_in[4] ,
    \sw_101_module_data_in[3] ,
    \sw_101_module_data_in[2] ,
    \sw_101_module_data_in[1] ,
    \sw_101_module_data_in[0] }),
    .io_out({\sw_101_module_data_out[7] ,
    \sw_101_module_data_out[6] ,
    \sw_101_module_data_out[5] ,
    \sw_101_module_data_out[4] ,
    \sw_101_module_data_out[3] ,
    \sw_101_module_data_out[2] ,
    \sw_101_module_data_out[1] ,
    \sw_101_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_102 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_102_module_data_in[7] ,
    \sw_102_module_data_in[6] ,
    \sw_102_module_data_in[5] ,
    \sw_102_module_data_in[4] ,
    \sw_102_module_data_in[3] ,
    \sw_102_module_data_in[2] ,
    \sw_102_module_data_in[1] ,
    \sw_102_module_data_in[0] }),
    .io_out({\sw_102_module_data_out[7] ,
    \sw_102_module_data_out[6] ,
    \sw_102_module_data_out[5] ,
    \sw_102_module_data_out[4] ,
    \sw_102_module_data_out[3] ,
    \sw_102_module_data_out[2] ,
    \sw_102_module_data_out[1] ,
    \sw_102_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_103 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_103_module_data_in[7] ,
    \sw_103_module_data_in[6] ,
    \sw_103_module_data_in[5] ,
    \sw_103_module_data_in[4] ,
    \sw_103_module_data_in[3] ,
    \sw_103_module_data_in[2] ,
    \sw_103_module_data_in[1] ,
    \sw_103_module_data_in[0] }),
    .io_out({\sw_103_module_data_out[7] ,
    \sw_103_module_data_out[6] ,
    \sw_103_module_data_out[5] ,
    \sw_103_module_data_out[4] ,
    \sw_103_module_data_out[3] ,
    \sw_103_module_data_out[2] ,
    \sw_103_module_data_out[1] ,
    \sw_103_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_104 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_104_module_data_in[7] ,
    \sw_104_module_data_in[6] ,
    \sw_104_module_data_in[5] ,
    \sw_104_module_data_in[4] ,
    \sw_104_module_data_in[3] ,
    \sw_104_module_data_in[2] ,
    \sw_104_module_data_in[1] ,
    \sw_104_module_data_in[0] }),
    .io_out({\sw_104_module_data_out[7] ,
    \sw_104_module_data_out[6] ,
    \sw_104_module_data_out[5] ,
    \sw_104_module_data_out[4] ,
    \sw_104_module_data_out[3] ,
    \sw_104_module_data_out[2] ,
    \sw_104_module_data_out[1] ,
    \sw_104_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_105 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_105_module_data_in[7] ,
    \sw_105_module_data_in[6] ,
    \sw_105_module_data_in[5] ,
    \sw_105_module_data_in[4] ,
    \sw_105_module_data_in[3] ,
    \sw_105_module_data_in[2] ,
    \sw_105_module_data_in[1] ,
    \sw_105_module_data_in[0] }),
    .io_out({\sw_105_module_data_out[7] ,
    \sw_105_module_data_out[6] ,
    \sw_105_module_data_out[5] ,
    \sw_105_module_data_out[4] ,
    \sw_105_module_data_out[3] ,
    \sw_105_module_data_out[2] ,
    \sw_105_module_data_out[1] ,
    \sw_105_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_106 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_106_module_data_in[7] ,
    \sw_106_module_data_in[6] ,
    \sw_106_module_data_in[5] ,
    \sw_106_module_data_in[4] ,
    \sw_106_module_data_in[3] ,
    \sw_106_module_data_in[2] ,
    \sw_106_module_data_in[1] ,
    \sw_106_module_data_in[0] }),
    .io_out({\sw_106_module_data_out[7] ,
    \sw_106_module_data_out[6] ,
    \sw_106_module_data_out[5] ,
    \sw_106_module_data_out[4] ,
    \sw_106_module_data_out[3] ,
    \sw_106_module_data_out[2] ,
    \sw_106_module_data_out[1] ,
    \sw_106_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_107 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_107_module_data_in[7] ,
    \sw_107_module_data_in[6] ,
    \sw_107_module_data_in[5] ,
    \sw_107_module_data_in[4] ,
    \sw_107_module_data_in[3] ,
    \sw_107_module_data_in[2] ,
    \sw_107_module_data_in[1] ,
    \sw_107_module_data_in[0] }),
    .io_out({\sw_107_module_data_out[7] ,
    \sw_107_module_data_out[6] ,
    \sw_107_module_data_out[5] ,
    \sw_107_module_data_out[4] ,
    \sw_107_module_data_out[3] ,
    \sw_107_module_data_out[2] ,
    \sw_107_module_data_out[1] ,
    \sw_107_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_108 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_108_module_data_in[7] ,
    \sw_108_module_data_in[6] ,
    \sw_108_module_data_in[5] ,
    \sw_108_module_data_in[4] ,
    \sw_108_module_data_in[3] ,
    \sw_108_module_data_in[2] ,
    \sw_108_module_data_in[1] ,
    \sw_108_module_data_in[0] }),
    .io_out({\sw_108_module_data_out[7] ,
    \sw_108_module_data_out[6] ,
    \sw_108_module_data_out[5] ,
    \sw_108_module_data_out[4] ,
    \sw_108_module_data_out[3] ,
    \sw_108_module_data_out[2] ,
    \sw_108_module_data_out[1] ,
    \sw_108_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_109 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_109_module_data_in[7] ,
    \sw_109_module_data_in[6] ,
    \sw_109_module_data_in[5] ,
    \sw_109_module_data_in[4] ,
    \sw_109_module_data_in[3] ,
    \sw_109_module_data_in[2] ,
    \sw_109_module_data_in[1] ,
    \sw_109_module_data_in[0] }),
    .io_out({\sw_109_module_data_out[7] ,
    \sw_109_module_data_out[6] ,
    \sw_109_module_data_out[5] ,
    \sw_109_module_data_out[4] ,
    \sw_109_module_data_out[3] ,
    \sw_109_module_data_out[2] ,
    \sw_109_module_data_out[1] ,
    \sw_109_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_110 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_110_module_data_in[7] ,
    \sw_110_module_data_in[6] ,
    \sw_110_module_data_in[5] ,
    \sw_110_module_data_in[4] ,
    \sw_110_module_data_in[3] ,
    \sw_110_module_data_in[2] ,
    \sw_110_module_data_in[1] ,
    \sw_110_module_data_in[0] }),
    .io_out({\sw_110_module_data_out[7] ,
    \sw_110_module_data_out[6] ,
    \sw_110_module_data_out[5] ,
    \sw_110_module_data_out[4] ,
    \sw_110_module_data_out[3] ,
    \sw_110_module_data_out[2] ,
    \sw_110_module_data_out[1] ,
    \sw_110_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_111 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_111_module_data_in[7] ,
    \sw_111_module_data_in[6] ,
    \sw_111_module_data_in[5] ,
    \sw_111_module_data_in[4] ,
    \sw_111_module_data_in[3] ,
    \sw_111_module_data_in[2] ,
    \sw_111_module_data_in[1] ,
    \sw_111_module_data_in[0] }),
    .io_out({\sw_111_module_data_out[7] ,
    \sw_111_module_data_out[6] ,
    \sw_111_module_data_out[5] ,
    \sw_111_module_data_out[4] ,
    \sw_111_module_data_out[3] ,
    \sw_111_module_data_out[2] ,
    \sw_111_module_data_out[1] ,
    \sw_111_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_112 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_112_module_data_in[7] ,
    \sw_112_module_data_in[6] ,
    \sw_112_module_data_in[5] ,
    \sw_112_module_data_in[4] ,
    \sw_112_module_data_in[3] ,
    \sw_112_module_data_in[2] ,
    \sw_112_module_data_in[1] ,
    \sw_112_module_data_in[0] }),
    .io_out({\sw_112_module_data_out[7] ,
    \sw_112_module_data_out[6] ,
    \sw_112_module_data_out[5] ,
    \sw_112_module_data_out[4] ,
    \sw_112_module_data_out[3] ,
    \sw_112_module_data_out[2] ,
    \sw_112_module_data_out[1] ,
    \sw_112_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_113 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_113_module_data_in[7] ,
    \sw_113_module_data_in[6] ,
    \sw_113_module_data_in[5] ,
    \sw_113_module_data_in[4] ,
    \sw_113_module_data_in[3] ,
    \sw_113_module_data_in[2] ,
    \sw_113_module_data_in[1] ,
    \sw_113_module_data_in[0] }),
    .io_out({\sw_113_module_data_out[7] ,
    \sw_113_module_data_out[6] ,
    \sw_113_module_data_out[5] ,
    \sw_113_module_data_out[4] ,
    \sw_113_module_data_out[3] ,
    \sw_113_module_data_out[2] ,
    \sw_113_module_data_out[1] ,
    \sw_113_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_114 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_114_module_data_in[7] ,
    \sw_114_module_data_in[6] ,
    \sw_114_module_data_in[5] ,
    \sw_114_module_data_in[4] ,
    \sw_114_module_data_in[3] ,
    \sw_114_module_data_in[2] ,
    \sw_114_module_data_in[1] ,
    \sw_114_module_data_in[0] }),
    .io_out({\sw_114_module_data_out[7] ,
    \sw_114_module_data_out[6] ,
    \sw_114_module_data_out[5] ,
    \sw_114_module_data_out[4] ,
    \sw_114_module_data_out[3] ,
    \sw_114_module_data_out[2] ,
    \sw_114_module_data_out[1] ,
    \sw_114_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_115 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_115_module_data_in[7] ,
    \sw_115_module_data_in[6] ,
    \sw_115_module_data_in[5] ,
    \sw_115_module_data_in[4] ,
    \sw_115_module_data_in[3] ,
    \sw_115_module_data_in[2] ,
    \sw_115_module_data_in[1] ,
    \sw_115_module_data_in[0] }),
    .io_out({\sw_115_module_data_out[7] ,
    \sw_115_module_data_out[6] ,
    \sw_115_module_data_out[5] ,
    \sw_115_module_data_out[4] ,
    \sw_115_module_data_out[3] ,
    \sw_115_module_data_out[2] ,
    \sw_115_module_data_out[1] ,
    \sw_115_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_116 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_116_module_data_in[7] ,
    \sw_116_module_data_in[6] ,
    \sw_116_module_data_in[5] ,
    \sw_116_module_data_in[4] ,
    \sw_116_module_data_in[3] ,
    \sw_116_module_data_in[2] ,
    \sw_116_module_data_in[1] ,
    \sw_116_module_data_in[0] }),
    .io_out({\sw_116_module_data_out[7] ,
    \sw_116_module_data_out[6] ,
    \sw_116_module_data_out[5] ,
    \sw_116_module_data_out[4] ,
    \sw_116_module_data_out[3] ,
    \sw_116_module_data_out[2] ,
    \sw_116_module_data_out[1] ,
    \sw_116_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_117 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_117_module_data_in[7] ,
    \sw_117_module_data_in[6] ,
    \sw_117_module_data_in[5] ,
    \sw_117_module_data_in[4] ,
    \sw_117_module_data_in[3] ,
    \sw_117_module_data_in[2] ,
    \sw_117_module_data_in[1] ,
    \sw_117_module_data_in[0] }),
    .io_out({\sw_117_module_data_out[7] ,
    \sw_117_module_data_out[6] ,
    \sw_117_module_data_out[5] ,
    \sw_117_module_data_out[4] ,
    \sw_117_module_data_out[3] ,
    \sw_117_module_data_out[2] ,
    \sw_117_module_data_out[1] ,
    \sw_117_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_118 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_118_module_data_in[7] ,
    \sw_118_module_data_in[6] ,
    \sw_118_module_data_in[5] ,
    \sw_118_module_data_in[4] ,
    \sw_118_module_data_in[3] ,
    \sw_118_module_data_in[2] ,
    \sw_118_module_data_in[1] ,
    \sw_118_module_data_in[0] }),
    .io_out({\sw_118_module_data_out[7] ,
    \sw_118_module_data_out[6] ,
    \sw_118_module_data_out[5] ,
    \sw_118_module_data_out[4] ,
    \sw_118_module_data_out[3] ,
    \sw_118_module_data_out[2] ,
    \sw_118_module_data_out[1] ,
    \sw_118_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_119 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_119_module_data_in[7] ,
    \sw_119_module_data_in[6] ,
    \sw_119_module_data_in[5] ,
    \sw_119_module_data_in[4] ,
    \sw_119_module_data_in[3] ,
    \sw_119_module_data_in[2] ,
    \sw_119_module_data_in[1] ,
    \sw_119_module_data_in[0] }),
    .io_out({\sw_119_module_data_out[7] ,
    \sw_119_module_data_out[6] ,
    \sw_119_module_data_out[5] ,
    \sw_119_module_data_out[4] ,
    \sw_119_module_data_out[3] ,
    \sw_119_module_data_out[2] ,
    \sw_119_module_data_out[1] ,
    \sw_119_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_120 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_120_module_data_in[7] ,
    \sw_120_module_data_in[6] ,
    \sw_120_module_data_in[5] ,
    \sw_120_module_data_in[4] ,
    \sw_120_module_data_in[3] ,
    \sw_120_module_data_in[2] ,
    \sw_120_module_data_in[1] ,
    \sw_120_module_data_in[0] }),
    .io_out({\sw_120_module_data_out[7] ,
    \sw_120_module_data_out[6] ,
    \sw_120_module_data_out[5] ,
    \sw_120_module_data_out[4] ,
    \sw_120_module_data_out[3] ,
    \sw_120_module_data_out[2] ,
    \sw_120_module_data_out[1] ,
    \sw_120_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_121 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_121_module_data_in[7] ,
    \sw_121_module_data_in[6] ,
    \sw_121_module_data_in[5] ,
    \sw_121_module_data_in[4] ,
    \sw_121_module_data_in[3] ,
    \sw_121_module_data_in[2] ,
    \sw_121_module_data_in[1] ,
    \sw_121_module_data_in[0] }),
    .io_out({\sw_121_module_data_out[7] ,
    \sw_121_module_data_out[6] ,
    \sw_121_module_data_out[5] ,
    \sw_121_module_data_out[4] ,
    \sw_121_module_data_out[3] ,
    \sw_121_module_data_out[2] ,
    \sw_121_module_data_out[1] ,
    \sw_121_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_122 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_122_module_data_in[7] ,
    \sw_122_module_data_in[6] ,
    \sw_122_module_data_in[5] ,
    \sw_122_module_data_in[4] ,
    \sw_122_module_data_in[3] ,
    \sw_122_module_data_in[2] ,
    \sw_122_module_data_in[1] ,
    \sw_122_module_data_in[0] }),
    .io_out({\sw_122_module_data_out[7] ,
    \sw_122_module_data_out[6] ,
    \sw_122_module_data_out[5] ,
    \sw_122_module_data_out[4] ,
    \sw_122_module_data_out[3] ,
    \sw_122_module_data_out[2] ,
    \sw_122_module_data_out[1] ,
    \sw_122_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_123 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_123_module_data_in[7] ,
    \sw_123_module_data_in[6] ,
    \sw_123_module_data_in[5] ,
    \sw_123_module_data_in[4] ,
    \sw_123_module_data_in[3] ,
    \sw_123_module_data_in[2] ,
    \sw_123_module_data_in[1] ,
    \sw_123_module_data_in[0] }),
    .io_out({\sw_123_module_data_out[7] ,
    \sw_123_module_data_out[6] ,
    \sw_123_module_data_out[5] ,
    \sw_123_module_data_out[4] ,
    \sw_123_module_data_out[3] ,
    \sw_123_module_data_out[2] ,
    \sw_123_module_data_out[1] ,
    \sw_123_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_124 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_124_module_data_in[7] ,
    \sw_124_module_data_in[6] ,
    \sw_124_module_data_in[5] ,
    \sw_124_module_data_in[4] ,
    \sw_124_module_data_in[3] ,
    \sw_124_module_data_in[2] ,
    \sw_124_module_data_in[1] ,
    \sw_124_module_data_in[0] }),
    .io_out({\sw_124_module_data_out[7] ,
    \sw_124_module_data_out[6] ,
    \sw_124_module_data_out[5] ,
    \sw_124_module_data_out[4] ,
    \sw_124_module_data_out[3] ,
    \sw_124_module_data_out[2] ,
    \sw_124_module_data_out[1] ,
    \sw_124_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_125 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_125_module_data_in[7] ,
    \sw_125_module_data_in[6] ,
    \sw_125_module_data_in[5] ,
    \sw_125_module_data_in[4] ,
    \sw_125_module_data_in[3] ,
    \sw_125_module_data_in[2] ,
    \sw_125_module_data_in[1] ,
    \sw_125_module_data_in[0] }),
    .io_out({\sw_125_module_data_out[7] ,
    \sw_125_module_data_out[6] ,
    \sw_125_module_data_out[5] ,
    \sw_125_module_data_out[4] ,
    \sw_125_module_data_out[3] ,
    \sw_125_module_data_out[2] ,
    \sw_125_module_data_out[1] ,
    \sw_125_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_126 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_126_module_data_in[7] ,
    \sw_126_module_data_in[6] ,
    \sw_126_module_data_in[5] ,
    \sw_126_module_data_in[4] ,
    \sw_126_module_data_in[3] ,
    \sw_126_module_data_in[2] ,
    \sw_126_module_data_in[1] ,
    \sw_126_module_data_in[0] }),
    .io_out({\sw_126_module_data_out[7] ,
    \sw_126_module_data_out[6] ,
    \sw_126_module_data_out[5] ,
    \sw_126_module_data_out[4] ,
    \sw_126_module_data_out[3] ,
    \sw_126_module_data_out[2] ,
    \sw_126_module_data_out[1] ,
    \sw_126_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_127 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_127_module_data_in[7] ,
    \sw_127_module_data_in[6] ,
    \sw_127_module_data_in[5] ,
    \sw_127_module_data_in[4] ,
    \sw_127_module_data_in[3] ,
    \sw_127_module_data_in[2] ,
    \sw_127_module_data_in[1] ,
    \sw_127_module_data_in[0] }),
    .io_out({\sw_127_module_data_out[7] ,
    \sw_127_module_data_out[6] ,
    \sw_127_module_data_out[5] ,
    \sw_127_module_data_out[4] ,
    \sw_127_module_data_out[3] ,
    \sw_127_module_data_out[2] ,
    \sw_127_module_data_out[1] ,
    \sw_127_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_128 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_128_module_data_in[7] ,
    \sw_128_module_data_in[6] ,
    \sw_128_module_data_in[5] ,
    \sw_128_module_data_in[4] ,
    \sw_128_module_data_in[3] ,
    \sw_128_module_data_in[2] ,
    \sw_128_module_data_in[1] ,
    \sw_128_module_data_in[0] }),
    .io_out({\sw_128_module_data_out[7] ,
    \sw_128_module_data_out[6] ,
    \sw_128_module_data_out[5] ,
    \sw_128_module_data_out[4] ,
    \sw_128_module_data_out[3] ,
    \sw_128_module_data_out[2] ,
    \sw_128_module_data_out[1] ,
    \sw_128_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_129 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_129_module_data_in[7] ,
    \sw_129_module_data_in[6] ,
    \sw_129_module_data_in[5] ,
    \sw_129_module_data_in[4] ,
    \sw_129_module_data_in[3] ,
    \sw_129_module_data_in[2] ,
    \sw_129_module_data_in[1] ,
    \sw_129_module_data_in[0] }),
    .io_out({\sw_129_module_data_out[7] ,
    \sw_129_module_data_out[6] ,
    \sw_129_module_data_out[5] ,
    \sw_129_module_data_out[4] ,
    \sw_129_module_data_out[3] ,
    \sw_129_module_data_out[2] ,
    \sw_129_module_data_out[1] ,
    \sw_129_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_130 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_130_module_data_in[7] ,
    \sw_130_module_data_in[6] ,
    \sw_130_module_data_in[5] ,
    \sw_130_module_data_in[4] ,
    \sw_130_module_data_in[3] ,
    \sw_130_module_data_in[2] ,
    \sw_130_module_data_in[1] ,
    \sw_130_module_data_in[0] }),
    .io_out({\sw_130_module_data_out[7] ,
    \sw_130_module_data_out[6] ,
    \sw_130_module_data_out[5] ,
    \sw_130_module_data_out[4] ,
    \sw_130_module_data_out[3] ,
    \sw_130_module_data_out[2] ,
    \sw_130_module_data_out[1] ,
    \sw_130_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_131 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_131_module_data_in[7] ,
    \sw_131_module_data_in[6] ,
    \sw_131_module_data_in[5] ,
    \sw_131_module_data_in[4] ,
    \sw_131_module_data_in[3] ,
    \sw_131_module_data_in[2] ,
    \sw_131_module_data_in[1] ,
    \sw_131_module_data_in[0] }),
    .io_out({\sw_131_module_data_out[7] ,
    \sw_131_module_data_out[6] ,
    \sw_131_module_data_out[5] ,
    \sw_131_module_data_out[4] ,
    \sw_131_module_data_out[3] ,
    \sw_131_module_data_out[2] ,
    \sw_131_module_data_out[1] ,
    \sw_131_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_132 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_132_module_data_in[7] ,
    \sw_132_module_data_in[6] ,
    \sw_132_module_data_in[5] ,
    \sw_132_module_data_in[4] ,
    \sw_132_module_data_in[3] ,
    \sw_132_module_data_in[2] ,
    \sw_132_module_data_in[1] ,
    \sw_132_module_data_in[0] }),
    .io_out({\sw_132_module_data_out[7] ,
    \sw_132_module_data_out[6] ,
    \sw_132_module_data_out[5] ,
    \sw_132_module_data_out[4] ,
    \sw_132_module_data_out[3] ,
    \sw_132_module_data_out[2] ,
    \sw_132_module_data_out[1] ,
    \sw_132_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_133 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_133_module_data_in[7] ,
    \sw_133_module_data_in[6] ,
    \sw_133_module_data_in[5] ,
    \sw_133_module_data_in[4] ,
    \sw_133_module_data_in[3] ,
    \sw_133_module_data_in[2] ,
    \sw_133_module_data_in[1] ,
    \sw_133_module_data_in[0] }),
    .io_out({\sw_133_module_data_out[7] ,
    \sw_133_module_data_out[6] ,
    \sw_133_module_data_out[5] ,
    \sw_133_module_data_out[4] ,
    \sw_133_module_data_out[3] ,
    \sw_133_module_data_out[2] ,
    \sw_133_module_data_out[1] ,
    \sw_133_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_134 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_134_module_data_in[7] ,
    \sw_134_module_data_in[6] ,
    \sw_134_module_data_in[5] ,
    \sw_134_module_data_in[4] ,
    \sw_134_module_data_in[3] ,
    \sw_134_module_data_in[2] ,
    \sw_134_module_data_in[1] ,
    \sw_134_module_data_in[0] }),
    .io_out({\sw_134_module_data_out[7] ,
    \sw_134_module_data_out[6] ,
    \sw_134_module_data_out[5] ,
    \sw_134_module_data_out[4] ,
    \sw_134_module_data_out[3] ,
    \sw_134_module_data_out[2] ,
    \sw_134_module_data_out[1] ,
    \sw_134_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_135 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_135_module_data_in[7] ,
    \sw_135_module_data_in[6] ,
    \sw_135_module_data_in[5] ,
    \sw_135_module_data_in[4] ,
    \sw_135_module_data_in[3] ,
    \sw_135_module_data_in[2] ,
    \sw_135_module_data_in[1] ,
    \sw_135_module_data_in[0] }),
    .io_out({\sw_135_module_data_out[7] ,
    \sw_135_module_data_out[6] ,
    \sw_135_module_data_out[5] ,
    \sw_135_module_data_out[4] ,
    \sw_135_module_data_out[3] ,
    \sw_135_module_data_out[2] ,
    \sw_135_module_data_out[1] ,
    \sw_135_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_136 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_136_module_data_in[7] ,
    \sw_136_module_data_in[6] ,
    \sw_136_module_data_in[5] ,
    \sw_136_module_data_in[4] ,
    \sw_136_module_data_in[3] ,
    \sw_136_module_data_in[2] ,
    \sw_136_module_data_in[1] ,
    \sw_136_module_data_in[0] }),
    .io_out({\sw_136_module_data_out[7] ,
    \sw_136_module_data_out[6] ,
    \sw_136_module_data_out[5] ,
    \sw_136_module_data_out[4] ,
    \sw_136_module_data_out[3] ,
    \sw_136_module_data_out[2] ,
    \sw_136_module_data_out[1] ,
    \sw_136_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_137 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_137_module_data_in[7] ,
    \sw_137_module_data_in[6] ,
    \sw_137_module_data_in[5] ,
    \sw_137_module_data_in[4] ,
    \sw_137_module_data_in[3] ,
    \sw_137_module_data_in[2] ,
    \sw_137_module_data_in[1] ,
    \sw_137_module_data_in[0] }),
    .io_out({\sw_137_module_data_out[7] ,
    \sw_137_module_data_out[6] ,
    \sw_137_module_data_out[5] ,
    \sw_137_module_data_out[4] ,
    \sw_137_module_data_out[3] ,
    \sw_137_module_data_out[2] ,
    \sw_137_module_data_out[1] ,
    \sw_137_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_138 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_138_module_data_in[7] ,
    \sw_138_module_data_in[6] ,
    \sw_138_module_data_in[5] ,
    \sw_138_module_data_in[4] ,
    \sw_138_module_data_in[3] ,
    \sw_138_module_data_in[2] ,
    \sw_138_module_data_in[1] ,
    \sw_138_module_data_in[0] }),
    .io_out({\sw_138_module_data_out[7] ,
    \sw_138_module_data_out[6] ,
    \sw_138_module_data_out[5] ,
    \sw_138_module_data_out[4] ,
    \sw_138_module_data_out[3] ,
    \sw_138_module_data_out[2] ,
    \sw_138_module_data_out[1] ,
    \sw_138_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_139 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_139_module_data_in[7] ,
    \sw_139_module_data_in[6] ,
    \sw_139_module_data_in[5] ,
    \sw_139_module_data_in[4] ,
    \sw_139_module_data_in[3] ,
    \sw_139_module_data_in[2] ,
    \sw_139_module_data_in[1] ,
    \sw_139_module_data_in[0] }),
    .io_out({\sw_139_module_data_out[7] ,
    \sw_139_module_data_out[6] ,
    \sw_139_module_data_out[5] ,
    \sw_139_module_data_out[4] ,
    \sw_139_module_data_out[3] ,
    \sw_139_module_data_out[2] ,
    \sw_139_module_data_out[1] ,
    \sw_139_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_140 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_140_module_data_in[7] ,
    \sw_140_module_data_in[6] ,
    \sw_140_module_data_in[5] ,
    \sw_140_module_data_in[4] ,
    \sw_140_module_data_in[3] ,
    \sw_140_module_data_in[2] ,
    \sw_140_module_data_in[1] ,
    \sw_140_module_data_in[0] }),
    .io_out({\sw_140_module_data_out[7] ,
    \sw_140_module_data_out[6] ,
    \sw_140_module_data_out[5] ,
    \sw_140_module_data_out[4] ,
    \sw_140_module_data_out[3] ,
    \sw_140_module_data_out[2] ,
    \sw_140_module_data_out[1] ,
    \sw_140_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_141 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_141_module_data_in[7] ,
    \sw_141_module_data_in[6] ,
    \sw_141_module_data_in[5] ,
    \sw_141_module_data_in[4] ,
    \sw_141_module_data_in[3] ,
    \sw_141_module_data_in[2] ,
    \sw_141_module_data_in[1] ,
    \sw_141_module_data_in[0] }),
    .io_out({\sw_141_module_data_out[7] ,
    \sw_141_module_data_out[6] ,
    \sw_141_module_data_out[5] ,
    \sw_141_module_data_out[4] ,
    \sw_141_module_data_out[3] ,
    \sw_141_module_data_out[2] ,
    \sw_141_module_data_out[1] ,
    \sw_141_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_142 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_142_module_data_in[7] ,
    \sw_142_module_data_in[6] ,
    \sw_142_module_data_in[5] ,
    \sw_142_module_data_in[4] ,
    \sw_142_module_data_in[3] ,
    \sw_142_module_data_in[2] ,
    \sw_142_module_data_in[1] ,
    \sw_142_module_data_in[0] }),
    .io_out({\sw_142_module_data_out[7] ,
    \sw_142_module_data_out[6] ,
    \sw_142_module_data_out[5] ,
    \sw_142_module_data_out[4] ,
    \sw_142_module_data_out[3] ,
    \sw_142_module_data_out[2] ,
    \sw_142_module_data_out[1] ,
    \sw_142_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_143 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_143_module_data_in[7] ,
    \sw_143_module_data_in[6] ,
    \sw_143_module_data_in[5] ,
    \sw_143_module_data_in[4] ,
    \sw_143_module_data_in[3] ,
    \sw_143_module_data_in[2] ,
    \sw_143_module_data_in[1] ,
    \sw_143_module_data_in[0] }),
    .io_out({\sw_143_module_data_out[7] ,
    \sw_143_module_data_out[6] ,
    \sw_143_module_data_out[5] ,
    \sw_143_module_data_out[4] ,
    \sw_143_module_data_out[3] ,
    \sw_143_module_data_out[2] ,
    \sw_143_module_data_out[1] ,
    \sw_143_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_144 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_144_module_data_in[7] ,
    \sw_144_module_data_in[6] ,
    \sw_144_module_data_in[5] ,
    \sw_144_module_data_in[4] ,
    \sw_144_module_data_in[3] ,
    \sw_144_module_data_in[2] ,
    \sw_144_module_data_in[1] ,
    \sw_144_module_data_in[0] }),
    .io_out({\sw_144_module_data_out[7] ,
    \sw_144_module_data_out[6] ,
    \sw_144_module_data_out[5] ,
    \sw_144_module_data_out[4] ,
    \sw_144_module_data_out[3] ,
    \sw_144_module_data_out[2] ,
    \sw_144_module_data_out[1] ,
    \sw_144_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_145 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_145_module_data_in[7] ,
    \sw_145_module_data_in[6] ,
    \sw_145_module_data_in[5] ,
    \sw_145_module_data_in[4] ,
    \sw_145_module_data_in[3] ,
    \sw_145_module_data_in[2] ,
    \sw_145_module_data_in[1] ,
    \sw_145_module_data_in[0] }),
    .io_out({\sw_145_module_data_out[7] ,
    \sw_145_module_data_out[6] ,
    \sw_145_module_data_out[5] ,
    \sw_145_module_data_out[4] ,
    \sw_145_module_data_out[3] ,
    \sw_145_module_data_out[2] ,
    \sw_145_module_data_out[1] ,
    \sw_145_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_146 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_146_module_data_in[7] ,
    \sw_146_module_data_in[6] ,
    \sw_146_module_data_in[5] ,
    \sw_146_module_data_in[4] ,
    \sw_146_module_data_in[3] ,
    \sw_146_module_data_in[2] ,
    \sw_146_module_data_in[1] ,
    \sw_146_module_data_in[0] }),
    .io_out({\sw_146_module_data_out[7] ,
    \sw_146_module_data_out[6] ,
    \sw_146_module_data_out[5] ,
    \sw_146_module_data_out[4] ,
    \sw_146_module_data_out[3] ,
    \sw_146_module_data_out[2] ,
    \sw_146_module_data_out[1] ,
    \sw_146_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_147 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_147_module_data_in[7] ,
    \sw_147_module_data_in[6] ,
    \sw_147_module_data_in[5] ,
    \sw_147_module_data_in[4] ,
    \sw_147_module_data_in[3] ,
    \sw_147_module_data_in[2] ,
    \sw_147_module_data_in[1] ,
    \sw_147_module_data_in[0] }),
    .io_out({\sw_147_module_data_out[7] ,
    \sw_147_module_data_out[6] ,
    \sw_147_module_data_out[5] ,
    \sw_147_module_data_out[4] ,
    \sw_147_module_data_out[3] ,
    \sw_147_module_data_out[2] ,
    \sw_147_module_data_out[1] ,
    \sw_147_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_148 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_148_module_data_in[7] ,
    \sw_148_module_data_in[6] ,
    \sw_148_module_data_in[5] ,
    \sw_148_module_data_in[4] ,
    \sw_148_module_data_in[3] ,
    \sw_148_module_data_in[2] ,
    \sw_148_module_data_in[1] ,
    \sw_148_module_data_in[0] }),
    .io_out({\sw_148_module_data_out[7] ,
    \sw_148_module_data_out[6] ,
    \sw_148_module_data_out[5] ,
    \sw_148_module_data_out[4] ,
    \sw_148_module_data_out[3] ,
    \sw_148_module_data_out[2] ,
    \sw_148_module_data_out[1] ,
    \sw_148_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_149 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_149_module_data_in[7] ,
    \sw_149_module_data_in[6] ,
    \sw_149_module_data_in[5] ,
    \sw_149_module_data_in[4] ,
    \sw_149_module_data_in[3] ,
    \sw_149_module_data_in[2] ,
    \sw_149_module_data_in[1] ,
    \sw_149_module_data_in[0] }),
    .io_out({\sw_149_module_data_out[7] ,
    \sw_149_module_data_out[6] ,
    \sw_149_module_data_out[5] ,
    \sw_149_module_data_out[4] ,
    \sw_149_module_data_out[3] ,
    \sw_149_module_data_out[2] ,
    \sw_149_module_data_out[1] ,
    \sw_149_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_150 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_150_module_data_in[7] ,
    \sw_150_module_data_in[6] ,
    \sw_150_module_data_in[5] ,
    \sw_150_module_data_in[4] ,
    \sw_150_module_data_in[3] ,
    \sw_150_module_data_in[2] ,
    \sw_150_module_data_in[1] ,
    \sw_150_module_data_in[0] }),
    .io_out({\sw_150_module_data_out[7] ,
    \sw_150_module_data_out[6] ,
    \sw_150_module_data_out[5] ,
    \sw_150_module_data_out[4] ,
    \sw_150_module_data_out[3] ,
    \sw_150_module_data_out[2] ,
    \sw_150_module_data_out[1] ,
    \sw_150_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_151 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_151_module_data_in[7] ,
    \sw_151_module_data_in[6] ,
    \sw_151_module_data_in[5] ,
    \sw_151_module_data_in[4] ,
    \sw_151_module_data_in[3] ,
    \sw_151_module_data_in[2] ,
    \sw_151_module_data_in[1] ,
    \sw_151_module_data_in[0] }),
    .io_out({\sw_151_module_data_out[7] ,
    \sw_151_module_data_out[6] ,
    \sw_151_module_data_out[5] ,
    \sw_151_module_data_out[4] ,
    \sw_151_module_data_out[3] ,
    \sw_151_module_data_out[2] ,
    \sw_151_module_data_out[1] ,
    \sw_151_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_152 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_152_module_data_in[7] ,
    \sw_152_module_data_in[6] ,
    \sw_152_module_data_in[5] ,
    \sw_152_module_data_in[4] ,
    \sw_152_module_data_in[3] ,
    \sw_152_module_data_in[2] ,
    \sw_152_module_data_in[1] ,
    \sw_152_module_data_in[0] }),
    .io_out({\sw_152_module_data_out[7] ,
    \sw_152_module_data_out[6] ,
    \sw_152_module_data_out[5] ,
    \sw_152_module_data_out[4] ,
    \sw_152_module_data_out[3] ,
    \sw_152_module_data_out[2] ,
    \sw_152_module_data_out[1] ,
    \sw_152_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_153 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_153_module_data_in[7] ,
    \sw_153_module_data_in[6] ,
    \sw_153_module_data_in[5] ,
    \sw_153_module_data_in[4] ,
    \sw_153_module_data_in[3] ,
    \sw_153_module_data_in[2] ,
    \sw_153_module_data_in[1] ,
    \sw_153_module_data_in[0] }),
    .io_out({\sw_153_module_data_out[7] ,
    \sw_153_module_data_out[6] ,
    \sw_153_module_data_out[5] ,
    \sw_153_module_data_out[4] ,
    \sw_153_module_data_out[3] ,
    \sw_153_module_data_out[2] ,
    \sw_153_module_data_out[1] ,
    \sw_153_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_154 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_154_module_data_in[7] ,
    \sw_154_module_data_in[6] ,
    \sw_154_module_data_in[5] ,
    \sw_154_module_data_in[4] ,
    \sw_154_module_data_in[3] ,
    \sw_154_module_data_in[2] ,
    \sw_154_module_data_in[1] ,
    \sw_154_module_data_in[0] }),
    .io_out({\sw_154_module_data_out[7] ,
    \sw_154_module_data_out[6] ,
    \sw_154_module_data_out[5] ,
    \sw_154_module_data_out[4] ,
    \sw_154_module_data_out[3] ,
    \sw_154_module_data_out[2] ,
    \sw_154_module_data_out[1] ,
    \sw_154_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_155 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_155_module_data_in[7] ,
    \sw_155_module_data_in[6] ,
    \sw_155_module_data_in[5] ,
    \sw_155_module_data_in[4] ,
    \sw_155_module_data_in[3] ,
    \sw_155_module_data_in[2] ,
    \sw_155_module_data_in[1] ,
    \sw_155_module_data_in[0] }),
    .io_out({\sw_155_module_data_out[7] ,
    \sw_155_module_data_out[6] ,
    \sw_155_module_data_out[5] ,
    \sw_155_module_data_out[4] ,
    \sw_155_module_data_out[3] ,
    \sw_155_module_data_out[2] ,
    \sw_155_module_data_out[1] ,
    \sw_155_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_156 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_156_module_data_in[7] ,
    \sw_156_module_data_in[6] ,
    \sw_156_module_data_in[5] ,
    \sw_156_module_data_in[4] ,
    \sw_156_module_data_in[3] ,
    \sw_156_module_data_in[2] ,
    \sw_156_module_data_in[1] ,
    \sw_156_module_data_in[0] }),
    .io_out({\sw_156_module_data_out[7] ,
    \sw_156_module_data_out[6] ,
    \sw_156_module_data_out[5] ,
    \sw_156_module_data_out[4] ,
    \sw_156_module_data_out[3] ,
    \sw_156_module_data_out[2] ,
    \sw_156_module_data_out[1] ,
    \sw_156_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_157 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_157_module_data_in[7] ,
    \sw_157_module_data_in[6] ,
    \sw_157_module_data_in[5] ,
    \sw_157_module_data_in[4] ,
    \sw_157_module_data_in[3] ,
    \sw_157_module_data_in[2] ,
    \sw_157_module_data_in[1] ,
    \sw_157_module_data_in[0] }),
    .io_out({\sw_157_module_data_out[7] ,
    \sw_157_module_data_out[6] ,
    \sw_157_module_data_out[5] ,
    \sw_157_module_data_out[4] ,
    \sw_157_module_data_out[3] ,
    \sw_157_module_data_out[2] ,
    \sw_157_module_data_out[1] ,
    \sw_157_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_158 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_158_module_data_in[7] ,
    \sw_158_module_data_in[6] ,
    \sw_158_module_data_in[5] ,
    \sw_158_module_data_in[4] ,
    \sw_158_module_data_in[3] ,
    \sw_158_module_data_in[2] ,
    \sw_158_module_data_in[1] ,
    \sw_158_module_data_in[0] }),
    .io_out({\sw_158_module_data_out[7] ,
    \sw_158_module_data_out[6] ,
    \sw_158_module_data_out[5] ,
    \sw_158_module_data_out[4] ,
    \sw_158_module_data_out[3] ,
    \sw_158_module_data_out[2] ,
    \sw_158_module_data_out[1] ,
    \sw_158_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_159 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_159_module_data_in[7] ,
    \sw_159_module_data_in[6] ,
    \sw_159_module_data_in[5] ,
    \sw_159_module_data_in[4] ,
    \sw_159_module_data_in[3] ,
    \sw_159_module_data_in[2] ,
    \sw_159_module_data_in[1] ,
    \sw_159_module_data_in[0] }),
    .io_out({\sw_159_module_data_out[7] ,
    \sw_159_module_data_out[6] ,
    \sw_159_module_data_out[5] ,
    \sw_159_module_data_out[4] ,
    \sw_159_module_data_out[3] ,
    \sw_159_module_data_out[2] ,
    \sw_159_module_data_out[1] ,
    \sw_159_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_160 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_160_module_data_in[7] ,
    \sw_160_module_data_in[6] ,
    \sw_160_module_data_in[5] ,
    \sw_160_module_data_in[4] ,
    \sw_160_module_data_in[3] ,
    \sw_160_module_data_in[2] ,
    \sw_160_module_data_in[1] ,
    \sw_160_module_data_in[0] }),
    .io_out({\sw_160_module_data_out[7] ,
    \sw_160_module_data_out[6] ,
    \sw_160_module_data_out[5] ,
    \sw_160_module_data_out[4] ,
    \sw_160_module_data_out[3] ,
    \sw_160_module_data_out[2] ,
    \sw_160_module_data_out[1] ,
    \sw_160_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_161 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_161_module_data_in[7] ,
    \sw_161_module_data_in[6] ,
    \sw_161_module_data_in[5] ,
    \sw_161_module_data_in[4] ,
    \sw_161_module_data_in[3] ,
    \sw_161_module_data_in[2] ,
    \sw_161_module_data_in[1] ,
    \sw_161_module_data_in[0] }),
    .io_out({\sw_161_module_data_out[7] ,
    \sw_161_module_data_out[6] ,
    \sw_161_module_data_out[5] ,
    \sw_161_module_data_out[4] ,
    \sw_161_module_data_out[3] ,
    \sw_161_module_data_out[2] ,
    \sw_161_module_data_out[1] ,
    \sw_161_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_162 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_162_module_data_in[7] ,
    \sw_162_module_data_in[6] ,
    \sw_162_module_data_in[5] ,
    \sw_162_module_data_in[4] ,
    \sw_162_module_data_in[3] ,
    \sw_162_module_data_in[2] ,
    \sw_162_module_data_in[1] ,
    \sw_162_module_data_in[0] }),
    .io_out({\sw_162_module_data_out[7] ,
    \sw_162_module_data_out[6] ,
    \sw_162_module_data_out[5] ,
    \sw_162_module_data_out[4] ,
    \sw_162_module_data_out[3] ,
    \sw_162_module_data_out[2] ,
    \sw_162_module_data_out[1] ,
    \sw_162_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_163 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_163_module_data_in[7] ,
    \sw_163_module_data_in[6] ,
    \sw_163_module_data_in[5] ,
    \sw_163_module_data_in[4] ,
    \sw_163_module_data_in[3] ,
    \sw_163_module_data_in[2] ,
    \sw_163_module_data_in[1] ,
    \sw_163_module_data_in[0] }),
    .io_out({\sw_163_module_data_out[7] ,
    \sw_163_module_data_out[6] ,
    \sw_163_module_data_out[5] ,
    \sw_163_module_data_out[4] ,
    \sw_163_module_data_out[3] ,
    \sw_163_module_data_out[2] ,
    \sw_163_module_data_out[1] ,
    \sw_163_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_164 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_164_module_data_in[7] ,
    \sw_164_module_data_in[6] ,
    \sw_164_module_data_in[5] ,
    \sw_164_module_data_in[4] ,
    \sw_164_module_data_in[3] ,
    \sw_164_module_data_in[2] ,
    \sw_164_module_data_in[1] ,
    \sw_164_module_data_in[0] }),
    .io_out({\sw_164_module_data_out[7] ,
    \sw_164_module_data_out[6] ,
    \sw_164_module_data_out[5] ,
    \sw_164_module_data_out[4] ,
    \sw_164_module_data_out[3] ,
    \sw_164_module_data_out[2] ,
    \sw_164_module_data_out[1] ,
    \sw_164_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_165 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_165_module_data_in[7] ,
    \sw_165_module_data_in[6] ,
    \sw_165_module_data_in[5] ,
    \sw_165_module_data_in[4] ,
    \sw_165_module_data_in[3] ,
    \sw_165_module_data_in[2] ,
    \sw_165_module_data_in[1] ,
    \sw_165_module_data_in[0] }),
    .io_out({\sw_165_module_data_out[7] ,
    \sw_165_module_data_out[6] ,
    \sw_165_module_data_out[5] ,
    \sw_165_module_data_out[4] ,
    \sw_165_module_data_out[3] ,
    \sw_165_module_data_out[2] ,
    \sw_165_module_data_out[1] ,
    \sw_165_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_166 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_166_module_data_in[7] ,
    \sw_166_module_data_in[6] ,
    \sw_166_module_data_in[5] ,
    \sw_166_module_data_in[4] ,
    \sw_166_module_data_in[3] ,
    \sw_166_module_data_in[2] ,
    \sw_166_module_data_in[1] ,
    \sw_166_module_data_in[0] }),
    .io_out({\sw_166_module_data_out[7] ,
    \sw_166_module_data_out[6] ,
    \sw_166_module_data_out[5] ,
    \sw_166_module_data_out[4] ,
    \sw_166_module_data_out[3] ,
    \sw_166_module_data_out[2] ,
    \sw_166_module_data_out[1] ,
    \sw_166_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_167 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_167_module_data_in[7] ,
    \sw_167_module_data_in[6] ,
    \sw_167_module_data_in[5] ,
    \sw_167_module_data_in[4] ,
    \sw_167_module_data_in[3] ,
    \sw_167_module_data_in[2] ,
    \sw_167_module_data_in[1] ,
    \sw_167_module_data_in[0] }),
    .io_out({\sw_167_module_data_out[7] ,
    \sw_167_module_data_out[6] ,
    \sw_167_module_data_out[5] ,
    \sw_167_module_data_out[4] ,
    \sw_167_module_data_out[3] ,
    \sw_167_module_data_out[2] ,
    \sw_167_module_data_out[1] ,
    \sw_167_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_168 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_168_module_data_in[7] ,
    \sw_168_module_data_in[6] ,
    \sw_168_module_data_in[5] ,
    \sw_168_module_data_in[4] ,
    \sw_168_module_data_in[3] ,
    \sw_168_module_data_in[2] ,
    \sw_168_module_data_in[1] ,
    \sw_168_module_data_in[0] }),
    .io_out({\sw_168_module_data_out[7] ,
    \sw_168_module_data_out[6] ,
    \sw_168_module_data_out[5] ,
    \sw_168_module_data_out[4] ,
    \sw_168_module_data_out[3] ,
    \sw_168_module_data_out[2] ,
    \sw_168_module_data_out[1] ,
    \sw_168_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_169 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_169_module_data_in[7] ,
    \sw_169_module_data_in[6] ,
    \sw_169_module_data_in[5] ,
    \sw_169_module_data_in[4] ,
    \sw_169_module_data_in[3] ,
    \sw_169_module_data_in[2] ,
    \sw_169_module_data_in[1] ,
    \sw_169_module_data_in[0] }),
    .io_out({\sw_169_module_data_out[7] ,
    \sw_169_module_data_out[6] ,
    \sw_169_module_data_out[5] ,
    \sw_169_module_data_out[4] ,
    \sw_169_module_data_out[3] ,
    \sw_169_module_data_out[2] ,
    \sw_169_module_data_out[1] ,
    \sw_169_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_170 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_170_module_data_in[7] ,
    \sw_170_module_data_in[6] ,
    \sw_170_module_data_in[5] ,
    \sw_170_module_data_in[4] ,
    \sw_170_module_data_in[3] ,
    \sw_170_module_data_in[2] ,
    \sw_170_module_data_in[1] ,
    \sw_170_module_data_in[0] }),
    .io_out({\sw_170_module_data_out[7] ,
    \sw_170_module_data_out[6] ,
    \sw_170_module_data_out[5] ,
    \sw_170_module_data_out[4] ,
    \sw_170_module_data_out[3] ,
    \sw_170_module_data_out[2] ,
    \sw_170_module_data_out[1] ,
    \sw_170_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_171 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_171_module_data_in[7] ,
    \sw_171_module_data_in[6] ,
    \sw_171_module_data_in[5] ,
    \sw_171_module_data_in[4] ,
    \sw_171_module_data_in[3] ,
    \sw_171_module_data_in[2] ,
    \sw_171_module_data_in[1] ,
    \sw_171_module_data_in[0] }),
    .io_out({\sw_171_module_data_out[7] ,
    \sw_171_module_data_out[6] ,
    \sw_171_module_data_out[5] ,
    \sw_171_module_data_out[4] ,
    \sw_171_module_data_out[3] ,
    \sw_171_module_data_out[2] ,
    \sw_171_module_data_out[1] ,
    \sw_171_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_172 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_172_module_data_in[7] ,
    \sw_172_module_data_in[6] ,
    \sw_172_module_data_in[5] ,
    \sw_172_module_data_in[4] ,
    \sw_172_module_data_in[3] ,
    \sw_172_module_data_in[2] ,
    \sw_172_module_data_in[1] ,
    \sw_172_module_data_in[0] }),
    .io_out({\sw_172_module_data_out[7] ,
    \sw_172_module_data_out[6] ,
    \sw_172_module_data_out[5] ,
    \sw_172_module_data_out[4] ,
    \sw_172_module_data_out[3] ,
    \sw_172_module_data_out[2] ,
    \sw_172_module_data_out[1] ,
    \sw_172_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_173 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_173_module_data_in[7] ,
    \sw_173_module_data_in[6] ,
    \sw_173_module_data_in[5] ,
    \sw_173_module_data_in[4] ,
    \sw_173_module_data_in[3] ,
    \sw_173_module_data_in[2] ,
    \sw_173_module_data_in[1] ,
    \sw_173_module_data_in[0] }),
    .io_out({\sw_173_module_data_out[7] ,
    \sw_173_module_data_out[6] ,
    \sw_173_module_data_out[5] ,
    \sw_173_module_data_out[4] ,
    \sw_173_module_data_out[3] ,
    \sw_173_module_data_out[2] ,
    \sw_173_module_data_out[1] ,
    \sw_173_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_174 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_174_module_data_in[7] ,
    \sw_174_module_data_in[6] ,
    \sw_174_module_data_in[5] ,
    \sw_174_module_data_in[4] ,
    \sw_174_module_data_in[3] ,
    \sw_174_module_data_in[2] ,
    \sw_174_module_data_in[1] ,
    \sw_174_module_data_in[0] }),
    .io_out({\sw_174_module_data_out[7] ,
    \sw_174_module_data_out[6] ,
    \sw_174_module_data_out[5] ,
    \sw_174_module_data_out[4] ,
    \sw_174_module_data_out[3] ,
    \sw_174_module_data_out[2] ,
    \sw_174_module_data_out[1] ,
    \sw_174_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_175 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_175_module_data_in[7] ,
    \sw_175_module_data_in[6] ,
    \sw_175_module_data_in[5] ,
    \sw_175_module_data_in[4] ,
    \sw_175_module_data_in[3] ,
    \sw_175_module_data_in[2] ,
    \sw_175_module_data_in[1] ,
    \sw_175_module_data_in[0] }),
    .io_out({\sw_175_module_data_out[7] ,
    \sw_175_module_data_out[6] ,
    \sw_175_module_data_out[5] ,
    \sw_175_module_data_out[4] ,
    \sw_175_module_data_out[3] ,
    \sw_175_module_data_out[2] ,
    \sw_175_module_data_out[1] ,
    \sw_175_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_176 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_176_module_data_in[7] ,
    \sw_176_module_data_in[6] ,
    \sw_176_module_data_in[5] ,
    \sw_176_module_data_in[4] ,
    \sw_176_module_data_in[3] ,
    \sw_176_module_data_in[2] ,
    \sw_176_module_data_in[1] ,
    \sw_176_module_data_in[0] }),
    .io_out({\sw_176_module_data_out[7] ,
    \sw_176_module_data_out[6] ,
    \sw_176_module_data_out[5] ,
    \sw_176_module_data_out[4] ,
    \sw_176_module_data_out[3] ,
    \sw_176_module_data_out[2] ,
    \sw_176_module_data_out[1] ,
    \sw_176_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_177 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_177_module_data_in[7] ,
    \sw_177_module_data_in[6] ,
    \sw_177_module_data_in[5] ,
    \sw_177_module_data_in[4] ,
    \sw_177_module_data_in[3] ,
    \sw_177_module_data_in[2] ,
    \sw_177_module_data_in[1] ,
    \sw_177_module_data_in[0] }),
    .io_out({\sw_177_module_data_out[7] ,
    \sw_177_module_data_out[6] ,
    \sw_177_module_data_out[5] ,
    \sw_177_module_data_out[4] ,
    \sw_177_module_data_out[3] ,
    \sw_177_module_data_out[2] ,
    \sw_177_module_data_out[1] ,
    \sw_177_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_178 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_178_module_data_in[7] ,
    \sw_178_module_data_in[6] ,
    \sw_178_module_data_in[5] ,
    \sw_178_module_data_in[4] ,
    \sw_178_module_data_in[3] ,
    \sw_178_module_data_in[2] ,
    \sw_178_module_data_in[1] ,
    \sw_178_module_data_in[0] }),
    .io_out({\sw_178_module_data_out[7] ,
    \sw_178_module_data_out[6] ,
    \sw_178_module_data_out[5] ,
    \sw_178_module_data_out[4] ,
    \sw_178_module_data_out[3] ,
    \sw_178_module_data_out[2] ,
    \sw_178_module_data_out[1] ,
    \sw_178_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_179 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_179_module_data_in[7] ,
    \sw_179_module_data_in[6] ,
    \sw_179_module_data_in[5] ,
    \sw_179_module_data_in[4] ,
    \sw_179_module_data_in[3] ,
    \sw_179_module_data_in[2] ,
    \sw_179_module_data_in[1] ,
    \sw_179_module_data_in[0] }),
    .io_out({\sw_179_module_data_out[7] ,
    \sw_179_module_data_out[6] ,
    \sw_179_module_data_out[5] ,
    \sw_179_module_data_out[4] ,
    \sw_179_module_data_out[3] ,
    \sw_179_module_data_out[2] ,
    \sw_179_module_data_out[1] ,
    \sw_179_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_180 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_180_module_data_in[7] ,
    \sw_180_module_data_in[6] ,
    \sw_180_module_data_in[5] ,
    \sw_180_module_data_in[4] ,
    \sw_180_module_data_in[3] ,
    \sw_180_module_data_in[2] ,
    \sw_180_module_data_in[1] ,
    \sw_180_module_data_in[0] }),
    .io_out({\sw_180_module_data_out[7] ,
    \sw_180_module_data_out[6] ,
    \sw_180_module_data_out[5] ,
    \sw_180_module_data_out[4] ,
    \sw_180_module_data_out[3] ,
    \sw_180_module_data_out[2] ,
    \sw_180_module_data_out[1] ,
    \sw_180_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_181 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_181_module_data_in[7] ,
    \sw_181_module_data_in[6] ,
    \sw_181_module_data_in[5] ,
    \sw_181_module_data_in[4] ,
    \sw_181_module_data_in[3] ,
    \sw_181_module_data_in[2] ,
    \sw_181_module_data_in[1] ,
    \sw_181_module_data_in[0] }),
    .io_out({\sw_181_module_data_out[7] ,
    \sw_181_module_data_out[6] ,
    \sw_181_module_data_out[5] ,
    \sw_181_module_data_out[4] ,
    \sw_181_module_data_out[3] ,
    \sw_181_module_data_out[2] ,
    \sw_181_module_data_out[1] ,
    \sw_181_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_182 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_182_module_data_in[7] ,
    \sw_182_module_data_in[6] ,
    \sw_182_module_data_in[5] ,
    \sw_182_module_data_in[4] ,
    \sw_182_module_data_in[3] ,
    \sw_182_module_data_in[2] ,
    \sw_182_module_data_in[1] ,
    \sw_182_module_data_in[0] }),
    .io_out({\sw_182_module_data_out[7] ,
    \sw_182_module_data_out[6] ,
    \sw_182_module_data_out[5] ,
    \sw_182_module_data_out[4] ,
    \sw_182_module_data_out[3] ,
    \sw_182_module_data_out[2] ,
    \sw_182_module_data_out[1] ,
    \sw_182_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_183 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_183_module_data_in[7] ,
    \sw_183_module_data_in[6] ,
    \sw_183_module_data_in[5] ,
    \sw_183_module_data_in[4] ,
    \sw_183_module_data_in[3] ,
    \sw_183_module_data_in[2] ,
    \sw_183_module_data_in[1] ,
    \sw_183_module_data_in[0] }),
    .io_out({\sw_183_module_data_out[7] ,
    \sw_183_module_data_out[6] ,
    \sw_183_module_data_out[5] ,
    \sw_183_module_data_out[4] ,
    \sw_183_module_data_out[3] ,
    \sw_183_module_data_out[2] ,
    \sw_183_module_data_out[1] ,
    \sw_183_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_184 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_184_module_data_in[7] ,
    \sw_184_module_data_in[6] ,
    \sw_184_module_data_in[5] ,
    \sw_184_module_data_in[4] ,
    \sw_184_module_data_in[3] ,
    \sw_184_module_data_in[2] ,
    \sw_184_module_data_in[1] ,
    \sw_184_module_data_in[0] }),
    .io_out({\sw_184_module_data_out[7] ,
    \sw_184_module_data_out[6] ,
    \sw_184_module_data_out[5] ,
    \sw_184_module_data_out[4] ,
    \sw_184_module_data_out[3] ,
    \sw_184_module_data_out[2] ,
    \sw_184_module_data_out[1] ,
    \sw_184_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_185 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_185_module_data_in[7] ,
    \sw_185_module_data_in[6] ,
    \sw_185_module_data_in[5] ,
    \sw_185_module_data_in[4] ,
    \sw_185_module_data_in[3] ,
    \sw_185_module_data_in[2] ,
    \sw_185_module_data_in[1] ,
    \sw_185_module_data_in[0] }),
    .io_out({\sw_185_module_data_out[7] ,
    \sw_185_module_data_out[6] ,
    \sw_185_module_data_out[5] ,
    \sw_185_module_data_out[4] ,
    \sw_185_module_data_out[3] ,
    \sw_185_module_data_out[2] ,
    \sw_185_module_data_out[1] ,
    \sw_185_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_186 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_186_module_data_in[7] ,
    \sw_186_module_data_in[6] ,
    \sw_186_module_data_in[5] ,
    \sw_186_module_data_in[4] ,
    \sw_186_module_data_in[3] ,
    \sw_186_module_data_in[2] ,
    \sw_186_module_data_in[1] ,
    \sw_186_module_data_in[0] }),
    .io_out({\sw_186_module_data_out[7] ,
    \sw_186_module_data_out[6] ,
    \sw_186_module_data_out[5] ,
    \sw_186_module_data_out[4] ,
    \sw_186_module_data_out[3] ,
    \sw_186_module_data_out[2] ,
    \sw_186_module_data_out[1] ,
    \sw_186_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_187 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_187_module_data_in[7] ,
    \sw_187_module_data_in[6] ,
    \sw_187_module_data_in[5] ,
    \sw_187_module_data_in[4] ,
    \sw_187_module_data_in[3] ,
    \sw_187_module_data_in[2] ,
    \sw_187_module_data_in[1] ,
    \sw_187_module_data_in[0] }),
    .io_out({\sw_187_module_data_out[7] ,
    \sw_187_module_data_out[6] ,
    \sw_187_module_data_out[5] ,
    \sw_187_module_data_out[4] ,
    \sw_187_module_data_out[3] ,
    \sw_187_module_data_out[2] ,
    \sw_187_module_data_out[1] ,
    \sw_187_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_188 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_188_module_data_in[7] ,
    \sw_188_module_data_in[6] ,
    \sw_188_module_data_in[5] ,
    \sw_188_module_data_in[4] ,
    \sw_188_module_data_in[3] ,
    \sw_188_module_data_in[2] ,
    \sw_188_module_data_in[1] ,
    \sw_188_module_data_in[0] }),
    .io_out({\sw_188_module_data_out[7] ,
    \sw_188_module_data_out[6] ,
    \sw_188_module_data_out[5] ,
    \sw_188_module_data_out[4] ,
    \sw_188_module_data_out[3] ,
    \sw_188_module_data_out[2] ,
    \sw_188_module_data_out[1] ,
    \sw_188_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_189 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_189_module_data_in[7] ,
    \sw_189_module_data_in[6] ,
    \sw_189_module_data_in[5] ,
    \sw_189_module_data_in[4] ,
    \sw_189_module_data_in[3] ,
    \sw_189_module_data_in[2] ,
    \sw_189_module_data_in[1] ,
    \sw_189_module_data_in[0] }),
    .io_out({\sw_189_module_data_out[7] ,
    \sw_189_module_data_out[6] ,
    \sw_189_module_data_out[5] ,
    \sw_189_module_data_out[4] ,
    \sw_189_module_data_out[3] ,
    \sw_189_module_data_out[2] ,
    \sw_189_module_data_out[1] ,
    \sw_189_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_190 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_190_module_data_in[7] ,
    \sw_190_module_data_in[6] ,
    \sw_190_module_data_in[5] ,
    \sw_190_module_data_in[4] ,
    \sw_190_module_data_in[3] ,
    \sw_190_module_data_in[2] ,
    \sw_190_module_data_in[1] ,
    \sw_190_module_data_in[0] }),
    .io_out({\sw_190_module_data_out[7] ,
    \sw_190_module_data_out[6] ,
    \sw_190_module_data_out[5] ,
    \sw_190_module_data_out[4] ,
    \sw_190_module_data_out[3] ,
    \sw_190_module_data_out[2] ,
    \sw_190_module_data_out[1] ,
    \sw_190_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_191 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_191_module_data_in[7] ,
    \sw_191_module_data_in[6] ,
    \sw_191_module_data_in[5] ,
    \sw_191_module_data_in[4] ,
    \sw_191_module_data_in[3] ,
    \sw_191_module_data_in[2] ,
    \sw_191_module_data_in[1] ,
    \sw_191_module_data_in[0] }),
    .io_out({\sw_191_module_data_out[7] ,
    \sw_191_module_data_out[6] ,
    \sw_191_module_data_out[5] ,
    \sw_191_module_data_out[4] ,
    \sw_191_module_data_out[3] ,
    \sw_191_module_data_out[2] ,
    \sw_191_module_data_out[1] ,
    \sw_191_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_192 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_192_module_data_in[7] ,
    \sw_192_module_data_in[6] ,
    \sw_192_module_data_in[5] ,
    \sw_192_module_data_in[4] ,
    \sw_192_module_data_in[3] ,
    \sw_192_module_data_in[2] ,
    \sw_192_module_data_in[1] ,
    \sw_192_module_data_in[0] }),
    .io_out({\sw_192_module_data_out[7] ,
    \sw_192_module_data_out[6] ,
    \sw_192_module_data_out[5] ,
    \sw_192_module_data_out[4] ,
    \sw_192_module_data_out[3] ,
    \sw_192_module_data_out[2] ,
    \sw_192_module_data_out[1] ,
    \sw_192_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_193 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_193_module_data_in[7] ,
    \sw_193_module_data_in[6] ,
    \sw_193_module_data_in[5] ,
    \sw_193_module_data_in[4] ,
    \sw_193_module_data_in[3] ,
    \sw_193_module_data_in[2] ,
    \sw_193_module_data_in[1] ,
    \sw_193_module_data_in[0] }),
    .io_out({\sw_193_module_data_out[7] ,
    \sw_193_module_data_out[6] ,
    \sw_193_module_data_out[5] ,
    \sw_193_module_data_out[4] ,
    \sw_193_module_data_out[3] ,
    \sw_193_module_data_out[2] ,
    \sw_193_module_data_out[1] ,
    \sw_193_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_194 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_194_module_data_in[7] ,
    \sw_194_module_data_in[6] ,
    \sw_194_module_data_in[5] ,
    \sw_194_module_data_in[4] ,
    \sw_194_module_data_in[3] ,
    \sw_194_module_data_in[2] ,
    \sw_194_module_data_in[1] ,
    \sw_194_module_data_in[0] }),
    .io_out({\sw_194_module_data_out[7] ,
    \sw_194_module_data_out[6] ,
    \sw_194_module_data_out[5] ,
    \sw_194_module_data_out[4] ,
    \sw_194_module_data_out[3] ,
    \sw_194_module_data_out[2] ,
    \sw_194_module_data_out[1] ,
    \sw_194_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_195 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_195_module_data_in[7] ,
    \sw_195_module_data_in[6] ,
    \sw_195_module_data_in[5] ,
    \sw_195_module_data_in[4] ,
    \sw_195_module_data_in[3] ,
    \sw_195_module_data_in[2] ,
    \sw_195_module_data_in[1] ,
    \sw_195_module_data_in[0] }),
    .io_out({\sw_195_module_data_out[7] ,
    \sw_195_module_data_out[6] ,
    \sw_195_module_data_out[5] ,
    \sw_195_module_data_out[4] ,
    \sw_195_module_data_out[3] ,
    \sw_195_module_data_out[2] ,
    \sw_195_module_data_out[1] ,
    \sw_195_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_196 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_196_module_data_in[7] ,
    \sw_196_module_data_in[6] ,
    \sw_196_module_data_in[5] ,
    \sw_196_module_data_in[4] ,
    \sw_196_module_data_in[3] ,
    \sw_196_module_data_in[2] ,
    \sw_196_module_data_in[1] ,
    \sw_196_module_data_in[0] }),
    .io_out({\sw_196_module_data_out[7] ,
    \sw_196_module_data_out[6] ,
    \sw_196_module_data_out[5] ,
    \sw_196_module_data_out[4] ,
    \sw_196_module_data_out[3] ,
    \sw_196_module_data_out[2] ,
    \sw_196_module_data_out[1] ,
    \sw_196_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_197 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_197_module_data_in[7] ,
    \sw_197_module_data_in[6] ,
    \sw_197_module_data_in[5] ,
    \sw_197_module_data_in[4] ,
    \sw_197_module_data_in[3] ,
    \sw_197_module_data_in[2] ,
    \sw_197_module_data_in[1] ,
    \sw_197_module_data_in[0] }),
    .io_out({\sw_197_module_data_out[7] ,
    \sw_197_module_data_out[6] ,
    \sw_197_module_data_out[5] ,
    \sw_197_module_data_out[4] ,
    \sw_197_module_data_out[3] ,
    \sw_197_module_data_out[2] ,
    \sw_197_module_data_out[1] ,
    \sw_197_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_198 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_198_module_data_in[7] ,
    \sw_198_module_data_in[6] ,
    \sw_198_module_data_in[5] ,
    \sw_198_module_data_in[4] ,
    \sw_198_module_data_in[3] ,
    \sw_198_module_data_in[2] ,
    \sw_198_module_data_in[1] ,
    \sw_198_module_data_in[0] }),
    .io_out({\sw_198_module_data_out[7] ,
    \sw_198_module_data_out[6] ,
    \sw_198_module_data_out[5] ,
    \sw_198_module_data_out[4] ,
    \sw_198_module_data_out[3] ,
    \sw_198_module_data_out[2] ,
    \sw_198_module_data_out[1] ,
    \sw_198_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_199 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_199_module_data_in[7] ,
    \sw_199_module_data_in[6] ,
    \sw_199_module_data_in[5] ,
    \sw_199_module_data_in[4] ,
    \sw_199_module_data_in[3] ,
    \sw_199_module_data_in[2] ,
    \sw_199_module_data_in[1] ,
    \sw_199_module_data_in[0] }),
    .io_out({\sw_199_module_data_out[7] ,
    \sw_199_module_data_out[6] ,
    \sw_199_module_data_out[5] ,
    \sw_199_module_data_out[4] ,
    \sw_199_module_data_out[3] ,
    \sw_199_module_data_out[2] ,
    \sw_199_module_data_out[1] ,
    \sw_199_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_200 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_200_module_data_in[7] ,
    \sw_200_module_data_in[6] ,
    \sw_200_module_data_in[5] ,
    \sw_200_module_data_in[4] ,
    \sw_200_module_data_in[3] ,
    \sw_200_module_data_in[2] ,
    \sw_200_module_data_in[1] ,
    \sw_200_module_data_in[0] }),
    .io_out({\sw_200_module_data_out[7] ,
    \sw_200_module_data_out[6] ,
    \sw_200_module_data_out[5] ,
    \sw_200_module_data_out[4] ,
    \sw_200_module_data_out[3] ,
    \sw_200_module_data_out[2] ,
    \sw_200_module_data_out[1] ,
    \sw_200_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_201 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_201_module_data_in[7] ,
    \sw_201_module_data_in[6] ,
    \sw_201_module_data_in[5] ,
    \sw_201_module_data_in[4] ,
    \sw_201_module_data_in[3] ,
    \sw_201_module_data_in[2] ,
    \sw_201_module_data_in[1] ,
    \sw_201_module_data_in[0] }),
    .io_out({\sw_201_module_data_out[7] ,
    \sw_201_module_data_out[6] ,
    \sw_201_module_data_out[5] ,
    \sw_201_module_data_out[4] ,
    \sw_201_module_data_out[3] ,
    \sw_201_module_data_out[2] ,
    \sw_201_module_data_out[1] ,
    \sw_201_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_202 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_202_module_data_in[7] ,
    \sw_202_module_data_in[6] ,
    \sw_202_module_data_in[5] ,
    \sw_202_module_data_in[4] ,
    \sw_202_module_data_in[3] ,
    \sw_202_module_data_in[2] ,
    \sw_202_module_data_in[1] ,
    \sw_202_module_data_in[0] }),
    .io_out({\sw_202_module_data_out[7] ,
    \sw_202_module_data_out[6] ,
    \sw_202_module_data_out[5] ,
    \sw_202_module_data_out[4] ,
    \sw_202_module_data_out[3] ,
    \sw_202_module_data_out[2] ,
    \sw_202_module_data_out[1] ,
    \sw_202_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_203 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_203_module_data_in[7] ,
    \sw_203_module_data_in[6] ,
    \sw_203_module_data_in[5] ,
    \sw_203_module_data_in[4] ,
    \sw_203_module_data_in[3] ,
    \sw_203_module_data_in[2] ,
    \sw_203_module_data_in[1] ,
    \sw_203_module_data_in[0] }),
    .io_out({\sw_203_module_data_out[7] ,
    \sw_203_module_data_out[6] ,
    \sw_203_module_data_out[5] ,
    \sw_203_module_data_out[4] ,
    \sw_203_module_data_out[3] ,
    \sw_203_module_data_out[2] ,
    \sw_203_module_data_out[1] ,
    \sw_203_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_204 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_204_module_data_in[7] ,
    \sw_204_module_data_in[6] ,
    \sw_204_module_data_in[5] ,
    \sw_204_module_data_in[4] ,
    \sw_204_module_data_in[3] ,
    \sw_204_module_data_in[2] ,
    \sw_204_module_data_in[1] ,
    \sw_204_module_data_in[0] }),
    .io_out({\sw_204_module_data_out[7] ,
    \sw_204_module_data_out[6] ,
    \sw_204_module_data_out[5] ,
    \sw_204_module_data_out[4] ,
    \sw_204_module_data_out[3] ,
    \sw_204_module_data_out[2] ,
    \sw_204_module_data_out[1] ,
    \sw_204_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_205 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_205_module_data_in[7] ,
    \sw_205_module_data_in[6] ,
    \sw_205_module_data_in[5] ,
    \sw_205_module_data_in[4] ,
    \sw_205_module_data_in[3] ,
    \sw_205_module_data_in[2] ,
    \sw_205_module_data_in[1] ,
    \sw_205_module_data_in[0] }),
    .io_out({\sw_205_module_data_out[7] ,
    \sw_205_module_data_out[6] ,
    \sw_205_module_data_out[5] ,
    \sw_205_module_data_out[4] ,
    \sw_205_module_data_out[3] ,
    \sw_205_module_data_out[2] ,
    \sw_205_module_data_out[1] ,
    \sw_205_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_206 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_206_module_data_in[7] ,
    \sw_206_module_data_in[6] ,
    \sw_206_module_data_in[5] ,
    \sw_206_module_data_in[4] ,
    \sw_206_module_data_in[3] ,
    \sw_206_module_data_in[2] ,
    \sw_206_module_data_in[1] ,
    \sw_206_module_data_in[0] }),
    .io_out({\sw_206_module_data_out[7] ,
    \sw_206_module_data_out[6] ,
    \sw_206_module_data_out[5] ,
    \sw_206_module_data_out[4] ,
    \sw_206_module_data_out[3] ,
    \sw_206_module_data_out[2] ,
    \sw_206_module_data_out[1] ,
    \sw_206_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_207 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_207_module_data_in[7] ,
    \sw_207_module_data_in[6] ,
    \sw_207_module_data_in[5] ,
    \sw_207_module_data_in[4] ,
    \sw_207_module_data_in[3] ,
    \sw_207_module_data_in[2] ,
    \sw_207_module_data_in[1] ,
    \sw_207_module_data_in[0] }),
    .io_out({\sw_207_module_data_out[7] ,
    \sw_207_module_data_out[6] ,
    \sw_207_module_data_out[5] ,
    \sw_207_module_data_out[4] ,
    \sw_207_module_data_out[3] ,
    \sw_207_module_data_out[2] ,
    \sw_207_module_data_out[1] ,
    \sw_207_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_208 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_208_module_data_in[7] ,
    \sw_208_module_data_in[6] ,
    \sw_208_module_data_in[5] ,
    \sw_208_module_data_in[4] ,
    \sw_208_module_data_in[3] ,
    \sw_208_module_data_in[2] ,
    \sw_208_module_data_in[1] ,
    \sw_208_module_data_in[0] }),
    .io_out({\sw_208_module_data_out[7] ,
    \sw_208_module_data_out[6] ,
    \sw_208_module_data_out[5] ,
    \sw_208_module_data_out[4] ,
    \sw_208_module_data_out[3] ,
    \sw_208_module_data_out[2] ,
    \sw_208_module_data_out[1] ,
    \sw_208_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_209 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_209_module_data_in[7] ,
    \sw_209_module_data_in[6] ,
    \sw_209_module_data_in[5] ,
    \sw_209_module_data_in[4] ,
    \sw_209_module_data_in[3] ,
    \sw_209_module_data_in[2] ,
    \sw_209_module_data_in[1] ,
    \sw_209_module_data_in[0] }),
    .io_out({\sw_209_module_data_out[7] ,
    \sw_209_module_data_out[6] ,
    \sw_209_module_data_out[5] ,
    \sw_209_module_data_out[4] ,
    \sw_209_module_data_out[3] ,
    \sw_209_module_data_out[2] ,
    \sw_209_module_data_out[1] ,
    \sw_209_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_210 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_210_module_data_in[7] ,
    \sw_210_module_data_in[6] ,
    \sw_210_module_data_in[5] ,
    \sw_210_module_data_in[4] ,
    \sw_210_module_data_in[3] ,
    \sw_210_module_data_in[2] ,
    \sw_210_module_data_in[1] ,
    \sw_210_module_data_in[0] }),
    .io_out({\sw_210_module_data_out[7] ,
    \sw_210_module_data_out[6] ,
    \sw_210_module_data_out[5] ,
    \sw_210_module_data_out[4] ,
    \sw_210_module_data_out[3] ,
    \sw_210_module_data_out[2] ,
    \sw_210_module_data_out[1] ,
    \sw_210_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_211 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_211_module_data_in[7] ,
    \sw_211_module_data_in[6] ,
    \sw_211_module_data_in[5] ,
    \sw_211_module_data_in[4] ,
    \sw_211_module_data_in[3] ,
    \sw_211_module_data_in[2] ,
    \sw_211_module_data_in[1] ,
    \sw_211_module_data_in[0] }),
    .io_out({\sw_211_module_data_out[7] ,
    \sw_211_module_data_out[6] ,
    \sw_211_module_data_out[5] ,
    \sw_211_module_data_out[4] ,
    \sw_211_module_data_out[3] ,
    \sw_211_module_data_out[2] ,
    \sw_211_module_data_out[1] ,
    \sw_211_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_212 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_212_module_data_in[7] ,
    \sw_212_module_data_in[6] ,
    \sw_212_module_data_in[5] ,
    \sw_212_module_data_in[4] ,
    \sw_212_module_data_in[3] ,
    \sw_212_module_data_in[2] ,
    \sw_212_module_data_in[1] ,
    \sw_212_module_data_in[0] }),
    .io_out({\sw_212_module_data_out[7] ,
    \sw_212_module_data_out[6] ,
    \sw_212_module_data_out[5] ,
    \sw_212_module_data_out[4] ,
    \sw_212_module_data_out[3] ,
    \sw_212_module_data_out[2] ,
    \sw_212_module_data_out[1] ,
    \sw_212_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_213 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_213_module_data_in[7] ,
    \sw_213_module_data_in[6] ,
    \sw_213_module_data_in[5] ,
    \sw_213_module_data_in[4] ,
    \sw_213_module_data_in[3] ,
    \sw_213_module_data_in[2] ,
    \sw_213_module_data_in[1] ,
    \sw_213_module_data_in[0] }),
    .io_out({\sw_213_module_data_out[7] ,
    \sw_213_module_data_out[6] ,
    \sw_213_module_data_out[5] ,
    \sw_213_module_data_out[4] ,
    \sw_213_module_data_out[3] ,
    \sw_213_module_data_out[2] ,
    \sw_213_module_data_out[1] ,
    \sw_213_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_214 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_214_module_data_in[7] ,
    \sw_214_module_data_in[6] ,
    \sw_214_module_data_in[5] ,
    \sw_214_module_data_in[4] ,
    \sw_214_module_data_in[3] ,
    \sw_214_module_data_in[2] ,
    \sw_214_module_data_in[1] ,
    \sw_214_module_data_in[0] }),
    .io_out({\sw_214_module_data_out[7] ,
    \sw_214_module_data_out[6] ,
    \sw_214_module_data_out[5] ,
    \sw_214_module_data_out[4] ,
    \sw_214_module_data_out[3] ,
    \sw_214_module_data_out[2] ,
    \sw_214_module_data_out[1] ,
    \sw_214_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_215 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_215_module_data_in[7] ,
    \sw_215_module_data_in[6] ,
    \sw_215_module_data_in[5] ,
    \sw_215_module_data_in[4] ,
    \sw_215_module_data_in[3] ,
    \sw_215_module_data_in[2] ,
    \sw_215_module_data_in[1] ,
    \sw_215_module_data_in[0] }),
    .io_out({\sw_215_module_data_out[7] ,
    \sw_215_module_data_out[6] ,
    \sw_215_module_data_out[5] ,
    \sw_215_module_data_out[4] ,
    \sw_215_module_data_out[3] ,
    \sw_215_module_data_out[2] ,
    \sw_215_module_data_out[1] ,
    \sw_215_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_216 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_216_module_data_in[7] ,
    \sw_216_module_data_in[6] ,
    \sw_216_module_data_in[5] ,
    \sw_216_module_data_in[4] ,
    \sw_216_module_data_in[3] ,
    \sw_216_module_data_in[2] ,
    \sw_216_module_data_in[1] ,
    \sw_216_module_data_in[0] }),
    .io_out({\sw_216_module_data_out[7] ,
    \sw_216_module_data_out[6] ,
    \sw_216_module_data_out[5] ,
    \sw_216_module_data_out[4] ,
    \sw_216_module_data_out[3] ,
    \sw_216_module_data_out[2] ,
    \sw_216_module_data_out[1] ,
    \sw_216_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_217 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_217_module_data_in[7] ,
    \sw_217_module_data_in[6] ,
    \sw_217_module_data_in[5] ,
    \sw_217_module_data_in[4] ,
    \sw_217_module_data_in[3] ,
    \sw_217_module_data_in[2] ,
    \sw_217_module_data_in[1] ,
    \sw_217_module_data_in[0] }),
    .io_out({\sw_217_module_data_out[7] ,
    \sw_217_module_data_out[6] ,
    \sw_217_module_data_out[5] ,
    \sw_217_module_data_out[4] ,
    \sw_217_module_data_out[3] ,
    \sw_217_module_data_out[2] ,
    \sw_217_module_data_out[1] ,
    \sw_217_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_218 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_218_module_data_in[7] ,
    \sw_218_module_data_in[6] ,
    \sw_218_module_data_in[5] ,
    \sw_218_module_data_in[4] ,
    \sw_218_module_data_in[3] ,
    \sw_218_module_data_in[2] ,
    \sw_218_module_data_in[1] ,
    \sw_218_module_data_in[0] }),
    .io_out({\sw_218_module_data_out[7] ,
    \sw_218_module_data_out[6] ,
    \sw_218_module_data_out[5] ,
    \sw_218_module_data_out[4] ,
    \sw_218_module_data_out[3] ,
    \sw_218_module_data_out[2] ,
    \sw_218_module_data_out[1] ,
    \sw_218_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_219 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_219_module_data_in[7] ,
    \sw_219_module_data_in[6] ,
    \sw_219_module_data_in[5] ,
    \sw_219_module_data_in[4] ,
    \sw_219_module_data_in[3] ,
    \sw_219_module_data_in[2] ,
    \sw_219_module_data_in[1] ,
    \sw_219_module_data_in[0] }),
    .io_out({\sw_219_module_data_out[7] ,
    \sw_219_module_data_out[6] ,
    \sw_219_module_data_out[5] ,
    \sw_219_module_data_out[4] ,
    \sw_219_module_data_out[3] ,
    \sw_219_module_data_out[2] ,
    \sw_219_module_data_out[1] ,
    \sw_219_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_220 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_220_module_data_in[7] ,
    \sw_220_module_data_in[6] ,
    \sw_220_module_data_in[5] ,
    \sw_220_module_data_in[4] ,
    \sw_220_module_data_in[3] ,
    \sw_220_module_data_in[2] ,
    \sw_220_module_data_in[1] ,
    \sw_220_module_data_in[0] }),
    .io_out({\sw_220_module_data_out[7] ,
    \sw_220_module_data_out[6] ,
    \sw_220_module_data_out[5] ,
    \sw_220_module_data_out[4] ,
    \sw_220_module_data_out[3] ,
    \sw_220_module_data_out[2] ,
    \sw_220_module_data_out[1] ,
    \sw_220_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_221 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_221_module_data_in[7] ,
    \sw_221_module_data_in[6] ,
    \sw_221_module_data_in[5] ,
    \sw_221_module_data_in[4] ,
    \sw_221_module_data_in[3] ,
    \sw_221_module_data_in[2] ,
    \sw_221_module_data_in[1] ,
    \sw_221_module_data_in[0] }),
    .io_out({\sw_221_module_data_out[7] ,
    \sw_221_module_data_out[6] ,
    \sw_221_module_data_out[5] ,
    \sw_221_module_data_out[4] ,
    \sw_221_module_data_out[3] ,
    \sw_221_module_data_out[2] ,
    \sw_221_module_data_out[1] ,
    \sw_221_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_222 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_222_module_data_in[7] ,
    \sw_222_module_data_in[6] ,
    \sw_222_module_data_in[5] ,
    \sw_222_module_data_in[4] ,
    \sw_222_module_data_in[3] ,
    \sw_222_module_data_in[2] ,
    \sw_222_module_data_in[1] ,
    \sw_222_module_data_in[0] }),
    .io_out({\sw_222_module_data_out[7] ,
    \sw_222_module_data_out[6] ,
    \sw_222_module_data_out[5] ,
    \sw_222_module_data_out[4] ,
    \sw_222_module_data_out[3] ,
    \sw_222_module_data_out[2] ,
    \sw_222_module_data_out[1] ,
    \sw_222_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_223 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_223_module_data_in[7] ,
    \sw_223_module_data_in[6] ,
    \sw_223_module_data_in[5] ,
    \sw_223_module_data_in[4] ,
    \sw_223_module_data_in[3] ,
    \sw_223_module_data_in[2] ,
    \sw_223_module_data_in[1] ,
    \sw_223_module_data_in[0] }),
    .io_out({\sw_223_module_data_out[7] ,
    \sw_223_module_data_out[6] ,
    \sw_223_module_data_out[5] ,
    \sw_223_module_data_out[4] ,
    \sw_223_module_data_out[3] ,
    \sw_223_module_data_out[2] ,
    \sw_223_module_data_out[1] ,
    \sw_223_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_224 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_224_module_data_in[7] ,
    \sw_224_module_data_in[6] ,
    \sw_224_module_data_in[5] ,
    \sw_224_module_data_in[4] ,
    \sw_224_module_data_in[3] ,
    \sw_224_module_data_in[2] ,
    \sw_224_module_data_in[1] ,
    \sw_224_module_data_in[0] }),
    .io_out({\sw_224_module_data_out[7] ,
    \sw_224_module_data_out[6] ,
    \sw_224_module_data_out[5] ,
    \sw_224_module_data_out[4] ,
    \sw_224_module_data_out[3] ,
    \sw_224_module_data_out[2] ,
    \sw_224_module_data_out[1] ,
    \sw_224_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_225 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_225_module_data_in[7] ,
    \sw_225_module_data_in[6] ,
    \sw_225_module_data_in[5] ,
    \sw_225_module_data_in[4] ,
    \sw_225_module_data_in[3] ,
    \sw_225_module_data_in[2] ,
    \sw_225_module_data_in[1] ,
    \sw_225_module_data_in[0] }),
    .io_out({\sw_225_module_data_out[7] ,
    \sw_225_module_data_out[6] ,
    \sw_225_module_data_out[5] ,
    \sw_225_module_data_out[4] ,
    \sw_225_module_data_out[3] ,
    \sw_225_module_data_out[2] ,
    \sw_225_module_data_out[1] ,
    \sw_225_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_226 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_226_module_data_in[7] ,
    \sw_226_module_data_in[6] ,
    \sw_226_module_data_in[5] ,
    \sw_226_module_data_in[4] ,
    \sw_226_module_data_in[3] ,
    \sw_226_module_data_in[2] ,
    \sw_226_module_data_in[1] ,
    \sw_226_module_data_in[0] }),
    .io_out({\sw_226_module_data_out[7] ,
    \sw_226_module_data_out[6] ,
    \sw_226_module_data_out[5] ,
    \sw_226_module_data_out[4] ,
    \sw_226_module_data_out[3] ,
    \sw_226_module_data_out[2] ,
    \sw_226_module_data_out[1] ,
    \sw_226_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_227 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_227_module_data_in[7] ,
    \sw_227_module_data_in[6] ,
    \sw_227_module_data_in[5] ,
    \sw_227_module_data_in[4] ,
    \sw_227_module_data_in[3] ,
    \sw_227_module_data_in[2] ,
    \sw_227_module_data_in[1] ,
    \sw_227_module_data_in[0] }),
    .io_out({\sw_227_module_data_out[7] ,
    \sw_227_module_data_out[6] ,
    \sw_227_module_data_out[5] ,
    \sw_227_module_data_out[4] ,
    \sw_227_module_data_out[3] ,
    \sw_227_module_data_out[2] ,
    \sw_227_module_data_out[1] ,
    \sw_227_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_228 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_228_module_data_in[7] ,
    \sw_228_module_data_in[6] ,
    \sw_228_module_data_in[5] ,
    \sw_228_module_data_in[4] ,
    \sw_228_module_data_in[3] ,
    \sw_228_module_data_in[2] ,
    \sw_228_module_data_in[1] ,
    \sw_228_module_data_in[0] }),
    .io_out({\sw_228_module_data_out[7] ,
    \sw_228_module_data_out[6] ,
    \sw_228_module_data_out[5] ,
    \sw_228_module_data_out[4] ,
    \sw_228_module_data_out[3] ,
    \sw_228_module_data_out[2] ,
    \sw_228_module_data_out[1] ,
    \sw_228_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_229 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_229_module_data_in[7] ,
    \sw_229_module_data_in[6] ,
    \sw_229_module_data_in[5] ,
    \sw_229_module_data_in[4] ,
    \sw_229_module_data_in[3] ,
    \sw_229_module_data_in[2] ,
    \sw_229_module_data_in[1] ,
    \sw_229_module_data_in[0] }),
    .io_out({\sw_229_module_data_out[7] ,
    \sw_229_module_data_out[6] ,
    \sw_229_module_data_out[5] ,
    \sw_229_module_data_out[4] ,
    \sw_229_module_data_out[3] ,
    \sw_229_module_data_out[2] ,
    \sw_229_module_data_out[1] ,
    \sw_229_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_230 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_230_module_data_in[7] ,
    \sw_230_module_data_in[6] ,
    \sw_230_module_data_in[5] ,
    \sw_230_module_data_in[4] ,
    \sw_230_module_data_in[3] ,
    \sw_230_module_data_in[2] ,
    \sw_230_module_data_in[1] ,
    \sw_230_module_data_in[0] }),
    .io_out({\sw_230_module_data_out[7] ,
    \sw_230_module_data_out[6] ,
    \sw_230_module_data_out[5] ,
    \sw_230_module_data_out[4] ,
    \sw_230_module_data_out[3] ,
    \sw_230_module_data_out[2] ,
    \sw_230_module_data_out[1] ,
    \sw_230_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_231 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_231_module_data_in[7] ,
    \sw_231_module_data_in[6] ,
    \sw_231_module_data_in[5] ,
    \sw_231_module_data_in[4] ,
    \sw_231_module_data_in[3] ,
    \sw_231_module_data_in[2] ,
    \sw_231_module_data_in[1] ,
    \sw_231_module_data_in[0] }),
    .io_out({\sw_231_module_data_out[7] ,
    \sw_231_module_data_out[6] ,
    \sw_231_module_data_out[5] ,
    \sw_231_module_data_out[4] ,
    \sw_231_module_data_out[3] ,
    \sw_231_module_data_out[2] ,
    \sw_231_module_data_out[1] ,
    \sw_231_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_232 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_232_module_data_in[7] ,
    \sw_232_module_data_in[6] ,
    \sw_232_module_data_in[5] ,
    \sw_232_module_data_in[4] ,
    \sw_232_module_data_in[3] ,
    \sw_232_module_data_in[2] ,
    \sw_232_module_data_in[1] ,
    \sw_232_module_data_in[0] }),
    .io_out({\sw_232_module_data_out[7] ,
    \sw_232_module_data_out[6] ,
    \sw_232_module_data_out[5] ,
    \sw_232_module_data_out[4] ,
    \sw_232_module_data_out[3] ,
    \sw_232_module_data_out[2] ,
    \sw_232_module_data_out[1] ,
    \sw_232_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_233 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_233_module_data_in[7] ,
    \sw_233_module_data_in[6] ,
    \sw_233_module_data_in[5] ,
    \sw_233_module_data_in[4] ,
    \sw_233_module_data_in[3] ,
    \sw_233_module_data_in[2] ,
    \sw_233_module_data_in[1] ,
    \sw_233_module_data_in[0] }),
    .io_out({\sw_233_module_data_out[7] ,
    \sw_233_module_data_out[6] ,
    \sw_233_module_data_out[5] ,
    \sw_233_module_data_out[4] ,
    \sw_233_module_data_out[3] ,
    \sw_233_module_data_out[2] ,
    \sw_233_module_data_out[1] ,
    \sw_233_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_234 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_234_module_data_in[7] ,
    \sw_234_module_data_in[6] ,
    \sw_234_module_data_in[5] ,
    \sw_234_module_data_in[4] ,
    \sw_234_module_data_in[3] ,
    \sw_234_module_data_in[2] ,
    \sw_234_module_data_in[1] ,
    \sw_234_module_data_in[0] }),
    .io_out({\sw_234_module_data_out[7] ,
    \sw_234_module_data_out[6] ,
    \sw_234_module_data_out[5] ,
    \sw_234_module_data_out[4] ,
    \sw_234_module_data_out[3] ,
    \sw_234_module_data_out[2] ,
    \sw_234_module_data_out[1] ,
    \sw_234_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_235 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_235_module_data_in[7] ,
    \sw_235_module_data_in[6] ,
    \sw_235_module_data_in[5] ,
    \sw_235_module_data_in[4] ,
    \sw_235_module_data_in[3] ,
    \sw_235_module_data_in[2] ,
    \sw_235_module_data_in[1] ,
    \sw_235_module_data_in[0] }),
    .io_out({\sw_235_module_data_out[7] ,
    \sw_235_module_data_out[6] ,
    \sw_235_module_data_out[5] ,
    \sw_235_module_data_out[4] ,
    \sw_235_module_data_out[3] ,
    \sw_235_module_data_out[2] ,
    \sw_235_module_data_out[1] ,
    \sw_235_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_236 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_236_module_data_in[7] ,
    \sw_236_module_data_in[6] ,
    \sw_236_module_data_in[5] ,
    \sw_236_module_data_in[4] ,
    \sw_236_module_data_in[3] ,
    \sw_236_module_data_in[2] ,
    \sw_236_module_data_in[1] ,
    \sw_236_module_data_in[0] }),
    .io_out({\sw_236_module_data_out[7] ,
    \sw_236_module_data_out[6] ,
    \sw_236_module_data_out[5] ,
    \sw_236_module_data_out[4] ,
    \sw_236_module_data_out[3] ,
    \sw_236_module_data_out[2] ,
    \sw_236_module_data_out[1] ,
    \sw_236_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_237 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_237_module_data_in[7] ,
    \sw_237_module_data_in[6] ,
    \sw_237_module_data_in[5] ,
    \sw_237_module_data_in[4] ,
    \sw_237_module_data_in[3] ,
    \sw_237_module_data_in[2] ,
    \sw_237_module_data_in[1] ,
    \sw_237_module_data_in[0] }),
    .io_out({\sw_237_module_data_out[7] ,
    \sw_237_module_data_out[6] ,
    \sw_237_module_data_out[5] ,
    \sw_237_module_data_out[4] ,
    \sw_237_module_data_out[3] ,
    \sw_237_module_data_out[2] ,
    \sw_237_module_data_out[1] ,
    \sw_237_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_238 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_238_module_data_in[7] ,
    \sw_238_module_data_in[6] ,
    \sw_238_module_data_in[5] ,
    \sw_238_module_data_in[4] ,
    \sw_238_module_data_in[3] ,
    \sw_238_module_data_in[2] ,
    \sw_238_module_data_in[1] ,
    \sw_238_module_data_in[0] }),
    .io_out({\sw_238_module_data_out[7] ,
    \sw_238_module_data_out[6] ,
    \sw_238_module_data_out[5] ,
    \sw_238_module_data_out[4] ,
    \sw_238_module_data_out[3] ,
    \sw_238_module_data_out[2] ,
    \sw_238_module_data_out[1] ,
    \sw_238_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_239 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_239_module_data_in[7] ,
    \sw_239_module_data_in[6] ,
    \sw_239_module_data_in[5] ,
    \sw_239_module_data_in[4] ,
    \sw_239_module_data_in[3] ,
    \sw_239_module_data_in[2] ,
    \sw_239_module_data_in[1] ,
    \sw_239_module_data_in[0] }),
    .io_out({\sw_239_module_data_out[7] ,
    \sw_239_module_data_out[6] ,
    \sw_239_module_data_out[5] ,
    \sw_239_module_data_out[4] ,
    \sw_239_module_data_out[3] ,
    \sw_239_module_data_out[2] ,
    \sw_239_module_data_out[1] ,
    \sw_239_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_240 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_240_module_data_in[7] ,
    \sw_240_module_data_in[6] ,
    \sw_240_module_data_in[5] ,
    \sw_240_module_data_in[4] ,
    \sw_240_module_data_in[3] ,
    \sw_240_module_data_in[2] ,
    \sw_240_module_data_in[1] ,
    \sw_240_module_data_in[0] }),
    .io_out({\sw_240_module_data_out[7] ,
    \sw_240_module_data_out[6] ,
    \sw_240_module_data_out[5] ,
    \sw_240_module_data_out[4] ,
    \sw_240_module_data_out[3] ,
    \sw_240_module_data_out[2] ,
    \sw_240_module_data_out[1] ,
    \sw_240_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_241 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_241_module_data_in[7] ,
    \sw_241_module_data_in[6] ,
    \sw_241_module_data_in[5] ,
    \sw_241_module_data_in[4] ,
    \sw_241_module_data_in[3] ,
    \sw_241_module_data_in[2] ,
    \sw_241_module_data_in[1] ,
    \sw_241_module_data_in[0] }),
    .io_out({\sw_241_module_data_out[7] ,
    \sw_241_module_data_out[6] ,
    \sw_241_module_data_out[5] ,
    \sw_241_module_data_out[4] ,
    \sw_241_module_data_out[3] ,
    \sw_241_module_data_out[2] ,
    \sw_241_module_data_out[1] ,
    \sw_241_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_242 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_242_module_data_in[7] ,
    \sw_242_module_data_in[6] ,
    \sw_242_module_data_in[5] ,
    \sw_242_module_data_in[4] ,
    \sw_242_module_data_in[3] ,
    \sw_242_module_data_in[2] ,
    \sw_242_module_data_in[1] ,
    \sw_242_module_data_in[0] }),
    .io_out({\sw_242_module_data_out[7] ,
    \sw_242_module_data_out[6] ,
    \sw_242_module_data_out[5] ,
    \sw_242_module_data_out[4] ,
    \sw_242_module_data_out[3] ,
    \sw_242_module_data_out[2] ,
    \sw_242_module_data_out[1] ,
    \sw_242_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_243 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_243_module_data_in[7] ,
    \sw_243_module_data_in[6] ,
    \sw_243_module_data_in[5] ,
    \sw_243_module_data_in[4] ,
    \sw_243_module_data_in[3] ,
    \sw_243_module_data_in[2] ,
    \sw_243_module_data_in[1] ,
    \sw_243_module_data_in[0] }),
    .io_out({\sw_243_module_data_out[7] ,
    \sw_243_module_data_out[6] ,
    \sw_243_module_data_out[5] ,
    \sw_243_module_data_out[4] ,
    \sw_243_module_data_out[3] ,
    \sw_243_module_data_out[2] ,
    \sw_243_module_data_out[1] ,
    \sw_243_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_244 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_244_module_data_in[7] ,
    \sw_244_module_data_in[6] ,
    \sw_244_module_data_in[5] ,
    \sw_244_module_data_in[4] ,
    \sw_244_module_data_in[3] ,
    \sw_244_module_data_in[2] ,
    \sw_244_module_data_in[1] ,
    \sw_244_module_data_in[0] }),
    .io_out({\sw_244_module_data_out[7] ,
    \sw_244_module_data_out[6] ,
    \sw_244_module_data_out[5] ,
    \sw_244_module_data_out[4] ,
    \sw_244_module_data_out[3] ,
    \sw_244_module_data_out[2] ,
    \sw_244_module_data_out[1] ,
    \sw_244_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_245 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_245_module_data_in[7] ,
    \sw_245_module_data_in[6] ,
    \sw_245_module_data_in[5] ,
    \sw_245_module_data_in[4] ,
    \sw_245_module_data_in[3] ,
    \sw_245_module_data_in[2] ,
    \sw_245_module_data_in[1] ,
    \sw_245_module_data_in[0] }),
    .io_out({\sw_245_module_data_out[7] ,
    \sw_245_module_data_out[6] ,
    \sw_245_module_data_out[5] ,
    \sw_245_module_data_out[4] ,
    \sw_245_module_data_out[3] ,
    \sw_245_module_data_out[2] ,
    \sw_245_module_data_out[1] ,
    \sw_245_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_246 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_246_module_data_in[7] ,
    \sw_246_module_data_in[6] ,
    \sw_246_module_data_in[5] ,
    \sw_246_module_data_in[4] ,
    \sw_246_module_data_in[3] ,
    \sw_246_module_data_in[2] ,
    \sw_246_module_data_in[1] ,
    \sw_246_module_data_in[0] }),
    .io_out({\sw_246_module_data_out[7] ,
    \sw_246_module_data_out[6] ,
    \sw_246_module_data_out[5] ,
    \sw_246_module_data_out[4] ,
    \sw_246_module_data_out[3] ,
    \sw_246_module_data_out[2] ,
    \sw_246_module_data_out[1] ,
    \sw_246_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_247 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_247_module_data_in[7] ,
    \sw_247_module_data_in[6] ,
    \sw_247_module_data_in[5] ,
    \sw_247_module_data_in[4] ,
    \sw_247_module_data_in[3] ,
    \sw_247_module_data_in[2] ,
    \sw_247_module_data_in[1] ,
    \sw_247_module_data_in[0] }),
    .io_out({\sw_247_module_data_out[7] ,
    \sw_247_module_data_out[6] ,
    \sw_247_module_data_out[5] ,
    \sw_247_module_data_out[4] ,
    \sw_247_module_data_out[3] ,
    \sw_247_module_data_out[2] ,
    \sw_247_module_data_out[1] ,
    \sw_247_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_248 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_248_module_data_in[7] ,
    \sw_248_module_data_in[6] ,
    \sw_248_module_data_in[5] ,
    \sw_248_module_data_in[4] ,
    \sw_248_module_data_in[3] ,
    \sw_248_module_data_in[2] ,
    \sw_248_module_data_in[1] ,
    \sw_248_module_data_in[0] }),
    .io_out({\sw_248_module_data_out[7] ,
    \sw_248_module_data_out[6] ,
    \sw_248_module_data_out[5] ,
    \sw_248_module_data_out[4] ,
    \sw_248_module_data_out[3] ,
    \sw_248_module_data_out[2] ,
    \sw_248_module_data_out[1] ,
    \sw_248_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_249 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_249_module_data_in[7] ,
    \sw_249_module_data_in[6] ,
    \sw_249_module_data_in[5] ,
    \sw_249_module_data_in[4] ,
    \sw_249_module_data_in[3] ,
    \sw_249_module_data_in[2] ,
    \sw_249_module_data_in[1] ,
    \sw_249_module_data_in[0] }),
    .io_out({\sw_249_module_data_out[7] ,
    \sw_249_module_data_out[6] ,
    \sw_249_module_data_out[5] ,
    \sw_249_module_data_out[4] ,
    \sw_249_module_data_out[3] ,
    \sw_249_module_data_out[2] ,
    \sw_249_module_data_out[1] ,
    \sw_249_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_250 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_250_module_data_in[7] ,
    \sw_250_module_data_in[6] ,
    \sw_250_module_data_in[5] ,
    \sw_250_module_data_in[4] ,
    \sw_250_module_data_in[3] ,
    \sw_250_module_data_in[2] ,
    \sw_250_module_data_in[1] ,
    \sw_250_module_data_in[0] }),
    .io_out({\sw_250_module_data_out[7] ,
    \sw_250_module_data_out[6] ,
    \sw_250_module_data_out[5] ,
    \sw_250_module_data_out[4] ,
    \sw_250_module_data_out[3] ,
    \sw_250_module_data_out[2] ,
    \sw_250_module_data_out[1] ,
    \sw_250_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_251 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_251_module_data_in[7] ,
    \sw_251_module_data_in[6] ,
    \sw_251_module_data_in[5] ,
    \sw_251_module_data_in[4] ,
    \sw_251_module_data_in[3] ,
    \sw_251_module_data_in[2] ,
    \sw_251_module_data_in[1] ,
    \sw_251_module_data_in[0] }),
    .io_out({\sw_251_module_data_out[7] ,
    \sw_251_module_data_out[6] ,
    \sw_251_module_data_out[5] ,
    \sw_251_module_data_out[4] ,
    \sw_251_module_data_out[3] ,
    \sw_251_module_data_out[2] ,
    \sw_251_module_data_out[1] ,
    \sw_251_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_252 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_252_module_data_in[7] ,
    \sw_252_module_data_in[6] ,
    \sw_252_module_data_in[5] ,
    \sw_252_module_data_in[4] ,
    \sw_252_module_data_in[3] ,
    \sw_252_module_data_in[2] ,
    \sw_252_module_data_in[1] ,
    \sw_252_module_data_in[0] }),
    .io_out({\sw_252_module_data_out[7] ,
    \sw_252_module_data_out[6] ,
    \sw_252_module_data_out[5] ,
    \sw_252_module_data_out[4] ,
    \sw_252_module_data_out[3] ,
    \sw_252_module_data_out[2] ,
    \sw_252_module_data_out[1] ,
    \sw_252_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_253 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_253_module_data_in[7] ,
    \sw_253_module_data_in[6] ,
    \sw_253_module_data_in[5] ,
    \sw_253_module_data_in[4] ,
    \sw_253_module_data_in[3] ,
    \sw_253_module_data_in[2] ,
    \sw_253_module_data_in[1] ,
    \sw_253_module_data_in[0] }),
    .io_out({\sw_253_module_data_out[7] ,
    \sw_253_module_data_out[6] ,
    \sw_253_module_data_out[5] ,
    \sw_253_module_data_out[4] ,
    \sw_253_module_data_out[3] ,
    \sw_253_module_data_out[2] ,
    \sw_253_module_data_out[1] ,
    \sw_253_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_254 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_254_module_data_in[7] ,
    \sw_254_module_data_in[6] ,
    \sw_254_module_data_in[5] ,
    \sw_254_module_data_in[4] ,
    \sw_254_module_data_in[3] ,
    \sw_254_module_data_in[2] ,
    \sw_254_module_data_in[1] ,
    \sw_254_module_data_in[0] }),
    .io_out({\sw_254_module_data_out[7] ,
    \sw_254_module_data_out[6] ,
    \sw_254_module_data_out[5] ,
    \sw_254_module_data_out[4] ,
    \sw_254_module_data_out[3] ,
    \sw_254_module_data_out[2] ,
    \sw_254_module_data_out[1] ,
    \sw_254_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_255 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_255_module_data_in[7] ,
    \sw_255_module_data_in[6] ,
    \sw_255_module_data_in[5] ,
    \sw_255_module_data_in[4] ,
    \sw_255_module_data_in[3] ,
    \sw_255_module_data_in[2] ,
    \sw_255_module_data_in[1] ,
    \sw_255_module_data_in[0] }),
    .io_out({\sw_255_module_data_out[7] ,
    \sw_255_module_data_out[6] ,
    \sw_255_module_data_out[5] ,
    \sw_255_module_data_out[4] ,
    \sw_255_module_data_out[3] ,
    \sw_255_module_data_out[2] ,
    \sw_255_module_data_out[1] ,
    \sw_255_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_256 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_256_module_data_in[7] ,
    \sw_256_module_data_in[6] ,
    \sw_256_module_data_in[5] ,
    \sw_256_module_data_in[4] ,
    \sw_256_module_data_in[3] ,
    \sw_256_module_data_in[2] ,
    \sw_256_module_data_in[1] ,
    \sw_256_module_data_in[0] }),
    .io_out({\sw_256_module_data_out[7] ,
    \sw_256_module_data_out[6] ,
    \sw_256_module_data_out[5] ,
    \sw_256_module_data_out[4] ,
    \sw_256_module_data_out[3] ,
    \sw_256_module_data_out[2] ,
    \sw_256_module_data_out[1] ,
    \sw_256_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_257 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_257_module_data_in[7] ,
    \sw_257_module_data_in[6] ,
    \sw_257_module_data_in[5] ,
    \sw_257_module_data_in[4] ,
    \sw_257_module_data_in[3] ,
    \sw_257_module_data_in[2] ,
    \sw_257_module_data_in[1] ,
    \sw_257_module_data_in[0] }),
    .io_out({\sw_257_module_data_out[7] ,
    \sw_257_module_data_out[6] ,
    \sw_257_module_data_out[5] ,
    \sw_257_module_data_out[4] ,
    \sw_257_module_data_out[3] ,
    \sw_257_module_data_out[2] ,
    \sw_257_module_data_out[1] ,
    \sw_257_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_258 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_258_module_data_in[7] ,
    \sw_258_module_data_in[6] ,
    \sw_258_module_data_in[5] ,
    \sw_258_module_data_in[4] ,
    \sw_258_module_data_in[3] ,
    \sw_258_module_data_in[2] ,
    \sw_258_module_data_in[1] ,
    \sw_258_module_data_in[0] }),
    .io_out({\sw_258_module_data_out[7] ,
    \sw_258_module_data_out[6] ,
    \sw_258_module_data_out[5] ,
    \sw_258_module_data_out[4] ,
    \sw_258_module_data_out[3] ,
    \sw_258_module_data_out[2] ,
    \sw_258_module_data_out[1] ,
    \sw_258_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_259 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_259_module_data_in[7] ,
    \sw_259_module_data_in[6] ,
    \sw_259_module_data_in[5] ,
    \sw_259_module_data_in[4] ,
    \sw_259_module_data_in[3] ,
    \sw_259_module_data_in[2] ,
    \sw_259_module_data_in[1] ,
    \sw_259_module_data_in[0] }),
    .io_out({\sw_259_module_data_out[7] ,
    \sw_259_module_data_out[6] ,
    \sw_259_module_data_out[5] ,
    \sw_259_module_data_out[4] ,
    \sw_259_module_data_out[3] ,
    \sw_259_module_data_out[2] ,
    \sw_259_module_data_out[1] ,
    \sw_259_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_260 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_260_module_data_in[7] ,
    \sw_260_module_data_in[6] ,
    \sw_260_module_data_in[5] ,
    \sw_260_module_data_in[4] ,
    \sw_260_module_data_in[3] ,
    \sw_260_module_data_in[2] ,
    \sw_260_module_data_in[1] ,
    \sw_260_module_data_in[0] }),
    .io_out({\sw_260_module_data_out[7] ,
    \sw_260_module_data_out[6] ,
    \sw_260_module_data_out[5] ,
    \sw_260_module_data_out[4] ,
    \sw_260_module_data_out[3] ,
    \sw_260_module_data_out[2] ,
    \sw_260_module_data_out[1] ,
    \sw_260_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_261 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_261_module_data_in[7] ,
    \sw_261_module_data_in[6] ,
    \sw_261_module_data_in[5] ,
    \sw_261_module_data_in[4] ,
    \sw_261_module_data_in[3] ,
    \sw_261_module_data_in[2] ,
    \sw_261_module_data_in[1] ,
    \sw_261_module_data_in[0] }),
    .io_out({\sw_261_module_data_out[7] ,
    \sw_261_module_data_out[6] ,
    \sw_261_module_data_out[5] ,
    \sw_261_module_data_out[4] ,
    \sw_261_module_data_out[3] ,
    \sw_261_module_data_out[2] ,
    \sw_261_module_data_out[1] ,
    \sw_261_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_262 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_262_module_data_in[7] ,
    \sw_262_module_data_in[6] ,
    \sw_262_module_data_in[5] ,
    \sw_262_module_data_in[4] ,
    \sw_262_module_data_in[3] ,
    \sw_262_module_data_in[2] ,
    \sw_262_module_data_in[1] ,
    \sw_262_module_data_in[0] }),
    .io_out({\sw_262_module_data_out[7] ,
    \sw_262_module_data_out[6] ,
    \sw_262_module_data_out[5] ,
    \sw_262_module_data_out[4] ,
    \sw_262_module_data_out[3] ,
    \sw_262_module_data_out[2] ,
    \sw_262_module_data_out[1] ,
    \sw_262_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_263 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_263_module_data_in[7] ,
    \sw_263_module_data_in[6] ,
    \sw_263_module_data_in[5] ,
    \sw_263_module_data_in[4] ,
    \sw_263_module_data_in[3] ,
    \sw_263_module_data_in[2] ,
    \sw_263_module_data_in[1] ,
    \sw_263_module_data_in[0] }),
    .io_out({\sw_263_module_data_out[7] ,
    \sw_263_module_data_out[6] ,
    \sw_263_module_data_out[5] ,
    \sw_263_module_data_out[4] ,
    \sw_263_module_data_out[3] ,
    \sw_263_module_data_out[2] ,
    \sw_263_module_data_out[1] ,
    \sw_263_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_264 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_264_module_data_in[7] ,
    \sw_264_module_data_in[6] ,
    \sw_264_module_data_in[5] ,
    \sw_264_module_data_in[4] ,
    \sw_264_module_data_in[3] ,
    \sw_264_module_data_in[2] ,
    \sw_264_module_data_in[1] ,
    \sw_264_module_data_in[0] }),
    .io_out({\sw_264_module_data_out[7] ,
    \sw_264_module_data_out[6] ,
    \sw_264_module_data_out[5] ,
    \sw_264_module_data_out[4] ,
    \sw_264_module_data_out[3] ,
    \sw_264_module_data_out[2] ,
    \sw_264_module_data_out[1] ,
    \sw_264_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_265 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_265_module_data_in[7] ,
    \sw_265_module_data_in[6] ,
    \sw_265_module_data_in[5] ,
    \sw_265_module_data_in[4] ,
    \sw_265_module_data_in[3] ,
    \sw_265_module_data_in[2] ,
    \sw_265_module_data_in[1] ,
    \sw_265_module_data_in[0] }),
    .io_out({\sw_265_module_data_out[7] ,
    \sw_265_module_data_out[6] ,
    \sw_265_module_data_out[5] ,
    \sw_265_module_data_out[4] ,
    \sw_265_module_data_out[3] ,
    \sw_265_module_data_out[2] ,
    \sw_265_module_data_out[1] ,
    \sw_265_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_266 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_266_module_data_in[7] ,
    \sw_266_module_data_in[6] ,
    \sw_266_module_data_in[5] ,
    \sw_266_module_data_in[4] ,
    \sw_266_module_data_in[3] ,
    \sw_266_module_data_in[2] ,
    \sw_266_module_data_in[1] ,
    \sw_266_module_data_in[0] }),
    .io_out({\sw_266_module_data_out[7] ,
    \sw_266_module_data_out[6] ,
    \sw_266_module_data_out[5] ,
    \sw_266_module_data_out[4] ,
    \sw_266_module_data_out[3] ,
    \sw_266_module_data_out[2] ,
    \sw_266_module_data_out[1] ,
    \sw_266_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_267 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_267_module_data_in[7] ,
    \sw_267_module_data_in[6] ,
    \sw_267_module_data_in[5] ,
    \sw_267_module_data_in[4] ,
    \sw_267_module_data_in[3] ,
    \sw_267_module_data_in[2] ,
    \sw_267_module_data_in[1] ,
    \sw_267_module_data_in[0] }),
    .io_out({\sw_267_module_data_out[7] ,
    \sw_267_module_data_out[6] ,
    \sw_267_module_data_out[5] ,
    \sw_267_module_data_out[4] ,
    \sw_267_module_data_out[3] ,
    \sw_267_module_data_out[2] ,
    \sw_267_module_data_out[1] ,
    \sw_267_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_268 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_268_module_data_in[7] ,
    \sw_268_module_data_in[6] ,
    \sw_268_module_data_in[5] ,
    \sw_268_module_data_in[4] ,
    \sw_268_module_data_in[3] ,
    \sw_268_module_data_in[2] ,
    \sw_268_module_data_in[1] ,
    \sw_268_module_data_in[0] }),
    .io_out({\sw_268_module_data_out[7] ,
    \sw_268_module_data_out[6] ,
    \sw_268_module_data_out[5] ,
    \sw_268_module_data_out[4] ,
    \sw_268_module_data_out[3] ,
    \sw_268_module_data_out[2] ,
    \sw_268_module_data_out[1] ,
    \sw_268_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_269 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_269_module_data_in[7] ,
    \sw_269_module_data_in[6] ,
    \sw_269_module_data_in[5] ,
    \sw_269_module_data_in[4] ,
    \sw_269_module_data_in[3] ,
    \sw_269_module_data_in[2] ,
    \sw_269_module_data_in[1] ,
    \sw_269_module_data_in[0] }),
    .io_out({\sw_269_module_data_out[7] ,
    \sw_269_module_data_out[6] ,
    \sw_269_module_data_out[5] ,
    \sw_269_module_data_out[4] ,
    \sw_269_module_data_out[3] ,
    \sw_269_module_data_out[2] ,
    \sw_269_module_data_out[1] ,
    \sw_269_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_270 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_270_module_data_in[7] ,
    \sw_270_module_data_in[6] ,
    \sw_270_module_data_in[5] ,
    \sw_270_module_data_in[4] ,
    \sw_270_module_data_in[3] ,
    \sw_270_module_data_in[2] ,
    \sw_270_module_data_in[1] ,
    \sw_270_module_data_in[0] }),
    .io_out({\sw_270_module_data_out[7] ,
    \sw_270_module_data_out[6] ,
    \sw_270_module_data_out[5] ,
    \sw_270_module_data_out[4] ,
    \sw_270_module_data_out[3] ,
    \sw_270_module_data_out[2] ,
    \sw_270_module_data_out[1] ,
    \sw_270_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_271 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_271_module_data_in[7] ,
    \sw_271_module_data_in[6] ,
    \sw_271_module_data_in[5] ,
    \sw_271_module_data_in[4] ,
    \sw_271_module_data_in[3] ,
    \sw_271_module_data_in[2] ,
    \sw_271_module_data_in[1] ,
    \sw_271_module_data_in[0] }),
    .io_out({\sw_271_module_data_out[7] ,
    \sw_271_module_data_out[6] ,
    \sw_271_module_data_out[5] ,
    \sw_271_module_data_out[4] ,
    \sw_271_module_data_out[3] ,
    \sw_271_module_data_out[2] ,
    \sw_271_module_data_out[1] ,
    \sw_271_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_272 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_272_module_data_in[7] ,
    \sw_272_module_data_in[6] ,
    \sw_272_module_data_in[5] ,
    \sw_272_module_data_in[4] ,
    \sw_272_module_data_in[3] ,
    \sw_272_module_data_in[2] ,
    \sw_272_module_data_in[1] ,
    \sw_272_module_data_in[0] }),
    .io_out({\sw_272_module_data_out[7] ,
    \sw_272_module_data_out[6] ,
    \sw_272_module_data_out[5] ,
    \sw_272_module_data_out[4] ,
    \sw_272_module_data_out[3] ,
    \sw_272_module_data_out[2] ,
    \sw_272_module_data_out[1] ,
    \sw_272_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_273 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_273_module_data_in[7] ,
    \sw_273_module_data_in[6] ,
    \sw_273_module_data_in[5] ,
    \sw_273_module_data_in[4] ,
    \sw_273_module_data_in[3] ,
    \sw_273_module_data_in[2] ,
    \sw_273_module_data_in[1] ,
    \sw_273_module_data_in[0] }),
    .io_out({\sw_273_module_data_out[7] ,
    \sw_273_module_data_out[6] ,
    \sw_273_module_data_out[5] ,
    \sw_273_module_data_out[4] ,
    \sw_273_module_data_out[3] ,
    \sw_273_module_data_out[2] ,
    \sw_273_module_data_out[1] ,
    \sw_273_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_274 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_274_module_data_in[7] ,
    \sw_274_module_data_in[6] ,
    \sw_274_module_data_in[5] ,
    \sw_274_module_data_in[4] ,
    \sw_274_module_data_in[3] ,
    \sw_274_module_data_in[2] ,
    \sw_274_module_data_in[1] ,
    \sw_274_module_data_in[0] }),
    .io_out({\sw_274_module_data_out[7] ,
    \sw_274_module_data_out[6] ,
    \sw_274_module_data_out[5] ,
    \sw_274_module_data_out[4] ,
    \sw_274_module_data_out[3] ,
    \sw_274_module_data_out[2] ,
    \sw_274_module_data_out[1] ,
    \sw_274_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_275 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_275_module_data_in[7] ,
    \sw_275_module_data_in[6] ,
    \sw_275_module_data_in[5] ,
    \sw_275_module_data_in[4] ,
    \sw_275_module_data_in[3] ,
    \sw_275_module_data_in[2] ,
    \sw_275_module_data_in[1] ,
    \sw_275_module_data_in[0] }),
    .io_out({\sw_275_module_data_out[7] ,
    \sw_275_module_data_out[6] ,
    \sw_275_module_data_out[5] ,
    \sw_275_module_data_out[4] ,
    \sw_275_module_data_out[3] ,
    \sw_275_module_data_out[2] ,
    \sw_275_module_data_out[1] ,
    \sw_275_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_276 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_276_module_data_in[7] ,
    \sw_276_module_data_in[6] ,
    \sw_276_module_data_in[5] ,
    \sw_276_module_data_in[4] ,
    \sw_276_module_data_in[3] ,
    \sw_276_module_data_in[2] ,
    \sw_276_module_data_in[1] ,
    \sw_276_module_data_in[0] }),
    .io_out({\sw_276_module_data_out[7] ,
    \sw_276_module_data_out[6] ,
    \sw_276_module_data_out[5] ,
    \sw_276_module_data_out[4] ,
    \sw_276_module_data_out[3] ,
    \sw_276_module_data_out[2] ,
    \sw_276_module_data_out[1] ,
    \sw_276_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_277 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_277_module_data_in[7] ,
    \sw_277_module_data_in[6] ,
    \sw_277_module_data_in[5] ,
    \sw_277_module_data_in[4] ,
    \sw_277_module_data_in[3] ,
    \sw_277_module_data_in[2] ,
    \sw_277_module_data_in[1] ,
    \sw_277_module_data_in[0] }),
    .io_out({\sw_277_module_data_out[7] ,
    \sw_277_module_data_out[6] ,
    \sw_277_module_data_out[5] ,
    \sw_277_module_data_out[4] ,
    \sw_277_module_data_out[3] ,
    \sw_277_module_data_out[2] ,
    \sw_277_module_data_out[1] ,
    \sw_277_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_278 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_278_module_data_in[7] ,
    \sw_278_module_data_in[6] ,
    \sw_278_module_data_in[5] ,
    \sw_278_module_data_in[4] ,
    \sw_278_module_data_in[3] ,
    \sw_278_module_data_in[2] ,
    \sw_278_module_data_in[1] ,
    \sw_278_module_data_in[0] }),
    .io_out({\sw_278_module_data_out[7] ,
    \sw_278_module_data_out[6] ,
    \sw_278_module_data_out[5] ,
    \sw_278_module_data_out[4] ,
    \sw_278_module_data_out[3] ,
    \sw_278_module_data_out[2] ,
    \sw_278_module_data_out[1] ,
    \sw_278_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_279 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_279_module_data_in[7] ,
    \sw_279_module_data_in[6] ,
    \sw_279_module_data_in[5] ,
    \sw_279_module_data_in[4] ,
    \sw_279_module_data_in[3] ,
    \sw_279_module_data_in[2] ,
    \sw_279_module_data_in[1] ,
    \sw_279_module_data_in[0] }),
    .io_out({\sw_279_module_data_out[7] ,
    \sw_279_module_data_out[6] ,
    \sw_279_module_data_out[5] ,
    \sw_279_module_data_out[4] ,
    \sw_279_module_data_out[3] ,
    \sw_279_module_data_out[2] ,
    \sw_279_module_data_out[1] ,
    \sw_279_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_280 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_280_module_data_in[7] ,
    \sw_280_module_data_in[6] ,
    \sw_280_module_data_in[5] ,
    \sw_280_module_data_in[4] ,
    \sw_280_module_data_in[3] ,
    \sw_280_module_data_in[2] ,
    \sw_280_module_data_in[1] ,
    \sw_280_module_data_in[0] }),
    .io_out({\sw_280_module_data_out[7] ,
    \sw_280_module_data_out[6] ,
    \sw_280_module_data_out[5] ,
    \sw_280_module_data_out[4] ,
    \sw_280_module_data_out[3] ,
    \sw_280_module_data_out[2] ,
    \sw_280_module_data_out[1] ,
    \sw_280_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_281 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_281_module_data_in[7] ,
    \sw_281_module_data_in[6] ,
    \sw_281_module_data_in[5] ,
    \sw_281_module_data_in[4] ,
    \sw_281_module_data_in[3] ,
    \sw_281_module_data_in[2] ,
    \sw_281_module_data_in[1] ,
    \sw_281_module_data_in[0] }),
    .io_out({\sw_281_module_data_out[7] ,
    \sw_281_module_data_out[6] ,
    \sw_281_module_data_out[5] ,
    \sw_281_module_data_out[4] ,
    \sw_281_module_data_out[3] ,
    \sw_281_module_data_out[2] ,
    \sw_281_module_data_out[1] ,
    \sw_281_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_282 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_282_module_data_in[7] ,
    \sw_282_module_data_in[6] ,
    \sw_282_module_data_in[5] ,
    \sw_282_module_data_in[4] ,
    \sw_282_module_data_in[3] ,
    \sw_282_module_data_in[2] ,
    \sw_282_module_data_in[1] ,
    \sw_282_module_data_in[0] }),
    .io_out({\sw_282_module_data_out[7] ,
    \sw_282_module_data_out[6] ,
    \sw_282_module_data_out[5] ,
    \sw_282_module_data_out[4] ,
    \sw_282_module_data_out[3] ,
    \sw_282_module_data_out[2] ,
    \sw_282_module_data_out[1] ,
    \sw_282_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_283 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_283_module_data_in[7] ,
    \sw_283_module_data_in[6] ,
    \sw_283_module_data_in[5] ,
    \sw_283_module_data_in[4] ,
    \sw_283_module_data_in[3] ,
    \sw_283_module_data_in[2] ,
    \sw_283_module_data_in[1] ,
    \sw_283_module_data_in[0] }),
    .io_out({\sw_283_module_data_out[7] ,
    \sw_283_module_data_out[6] ,
    \sw_283_module_data_out[5] ,
    \sw_283_module_data_out[4] ,
    \sw_283_module_data_out[3] ,
    \sw_283_module_data_out[2] ,
    \sw_283_module_data_out[1] ,
    \sw_283_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_284 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_284_module_data_in[7] ,
    \sw_284_module_data_in[6] ,
    \sw_284_module_data_in[5] ,
    \sw_284_module_data_in[4] ,
    \sw_284_module_data_in[3] ,
    \sw_284_module_data_in[2] ,
    \sw_284_module_data_in[1] ,
    \sw_284_module_data_in[0] }),
    .io_out({\sw_284_module_data_out[7] ,
    \sw_284_module_data_out[6] ,
    \sw_284_module_data_out[5] ,
    \sw_284_module_data_out[4] ,
    \sw_284_module_data_out[3] ,
    \sw_284_module_data_out[2] ,
    \sw_284_module_data_out[1] ,
    \sw_284_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_285 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_285_module_data_in[7] ,
    \sw_285_module_data_in[6] ,
    \sw_285_module_data_in[5] ,
    \sw_285_module_data_in[4] ,
    \sw_285_module_data_in[3] ,
    \sw_285_module_data_in[2] ,
    \sw_285_module_data_in[1] ,
    \sw_285_module_data_in[0] }),
    .io_out({\sw_285_module_data_out[7] ,
    \sw_285_module_data_out[6] ,
    \sw_285_module_data_out[5] ,
    \sw_285_module_data_out[4] ,
    \sw_285_module_data_out[3] ,
    \sw_285_module_data_out[2] ,
    \sw_285_module_data_out[1] ,
    \sw_285_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_286 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_286_module_data_in[7] ,
    \sw_286_module_data_in[6] ,
    \sw_286_module_data_in[5] ,
    \sw_286_module_data_in[4] ,
    \sw_286_module_data_in[3] ,
    \sw_286_module_data_in[2] ,
    \sw_286_module_data_in[1] ,
    \sw_286_module_data_in[0] }),
    .io_out({\sw_286_module_data_out[7] ,
    \sw_286_module_data_out[6] ,
    \sw_286_module_data_out[5] ,
    \sw_286_module_data_out[4] ,
    \sw_286_module_data_out[3] ,
    \sw_286_module_data_out[2] ,
    \sw_286_module_data_out[1] ,
    \sw_286_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_287 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_287_module_data_in[7] ,
    \sw_287_module_data_in[6] ,
    \sw_287_module_data_in[5] ,
    \sw_287_module_data_in[4] ,
    \sw_287_module_data_in[3] ,
    \sw_287_module_data_in[2] ,
    \sw_287_module_data_in[1] ,
    \sw_287_module_data_in[0] }),
    .io_out({\sw_287_module_data_out[7] ,
    \sw_287_module_data_out[6] ,
    \sw_287_module_data_out[5] ,
    \sw_287_module_data_out[4] ,
    \sw_287_module_data_out[3] ,
    \sw_287_module_data_out[2] ,
    \sw_287_module_data_out[1] ,
    \sw_287_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_288 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_288_module_data_in[7] ,
    \sw_288_module_data_in[6] ,
    \sw_288_module_data_in[5] ,
    \sw_288_module_data_in[4] ,
    \sw_288_module_data_in[3] ,
    \sw_288_module_data_in[2] ,
    \sw_288_module_data_in[1] ,
    \sw_288_module_data_in[0] }),
    .io_out({\sw_288_module_data_out[7] ,
    \sw_288_module_data_out[6] ,
    \sw_288_module_data_out[5] ,
    \sw_288_module_data_out[4] ,
    \sw_288_module_data_out[3] ,
    \sw_288_module_data_out[2] ,
    \sw_288_module_data_out[1] ,
    \sw_288_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_289 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_289_module_data_in[7] ,
    \sw_289_module_data_in[6] ,
    \sw_289_module_data_in[5] ,
    \sw_289_module_data_in[4] ,
    \sw_289_module_data_in[3] ,
    \sw_289_module_data_in[2] ,
    \sw_289_module_data_in[1] ,
    \sw_289_module_data_in[0] }),
    .io_out({\sw_289_module_data_out[7] ,
    \sw_289_module_data_out[6] ,
    \sw_289_module_data_out[5] ,
    \sw_289_module_data_out[4] ,
    \sw_289_module_data_out[3] ,
    \sw_289_module_data_out[2] ,
    \sw_289_module_data_out[1] ,
    \sw_289_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_29 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_029_module_data_in[7] ,
    \sw_029_module_data_in[6] ,
    \sw_029_module_data_in[5] ,
    \sw_029_module_data_in[4] ,
    \sw_029_module_data_in[3] ,
    \sw_029_module_data_in[2] ,
    \sw_029_module_data_in[1] ,
    \sw_029_module_data_in[0] }),
    .io_out({\sw_029_module_data_out[7] ,
    \sw_029_module_data_out[6] ,
    \sw_029_module_data_out[5] ,
    \sw_029_module_data_out[4] ,
    \sw_029_module_data_out[3] ,
    \sw_029_module_data_out[2] ,
    \sw_029_module_data_out[1] ,
    \sw_029_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_290 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_290_module_data_in[7] ,
    \sw_290_module_data_in[6] ,
    \sw_290_module_data_in[5] ,
    \sw_290_module_data_in[4] ,
    \sw_290_module_data_in[3] ,
    \sw_290_module_data_in[2] ,
    \sw_290_module_data_in[1] ,
    \sw_290_module_data_in[0] }),
    .io_out({\sw_290_module_data_out[7] ,
    \sw_290_module_data_out[6] ,
    \sw_290_module_data_out[5] ,
    \sw_290_module_data_out[4] ,
    \sw_290_module_data_out[3] ,
    \sw_290_module_data_out[2] ,
    \sw_290_module_data_out[1] ,
    \sw_290_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_291 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_291_module_data_in[7] ,
    \sw_291_module_data_in[6] ,
    \sw_291_module_data_in[5] ,
    \sw_291_module_data_in[4] ,
    \sw_291_module_data_in[3] ,
    \sw_291_module_data_in[2] ,
    \sw_291_module_data_in[1] ,
    \sw_291_module_data_in[0] }),
    .io_out({\sw_291_module_data_out[7] ,
    \sw_291_module_data_out[6] ,
    \sw_291_module_data_out[5] ,
    \sw_291_module_data_out[4] ,
    \sw_291_module_data_out[3] ,
    \sw_291_module_data_out[2] ,
    \sw_291_module_data_out[1] ,
    \sw_291_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_292 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_292_module_data_in[7] ,
    \sw_292_module_data_in[6] ,
    \sw_292_module_data_in[5] ,
    \sw_292_module_data_in[4] ,
    \sw_292_module_data_in[3] ,
    \sw_292_module_data_in[2] ,
    \sw_292_module_data_in[1] ,
    \sw_292_module_data_in[0] }),
    .io_out({\sw_292_module_data_out[7] ,
    \sw_292_module_data_out[6] ,
    \sw_292_module_data_out[5] ,
    \sw_292_module_data_out[4] ,
    \sw_292_module_data_out[3] ,
    \sw_292_module_data_out[2] ,
    \sw_292_module_data_out[1] ,
    \sw_292_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_293 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_293_module_data_in[7] ,
    \sw_293_module_data_in[6] ,
    \sw_293_module_data_in[5] ,
    \sw_293_module_data_in[4] ,
    \sw_293_module_data_in[3] ,
    \sw_293_module_data_in[2] ,
    \sw_293_module_data_in[1] ,
    \sw_293_module_data_in[0] }),
    .io_out({\sw_293_module_data_out[7] ,
    \sw_293_module_data_out[6] ,
    \sw_293_module_data_out[5] ,
    \sw_293_module_data_out[4] ,
    \sw_293_module_data_out[3] ,
    \sw_293_module_data_out[2] ,
    \sw_293_module_data_out[1] ,
    \sw_293_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_294 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_294_module_data_in[7] ,
    \sw_294_module_data_in[6] ,
    \sw_294_module_data_in[5] ,
    \sw_294_module_data_in[4] ,
    \sw_294_module_data_in[3] ,
    \sw_294_module_data_in[2] ,
    \sw_294_module_data_in[1] ,
    \sw_294_module_data_in[0] }),
    .io_out({\sw_294_module_data_out[7] ,
    \sw_294_module_data_out[6] ,
    \sw_294_module_data_out[5] ,
    \sw_294_module_data_out[4] ,
    \sw_294_module_data_out[3] ,
    \sw_294_module_data_out[2] ,
    \sw_294_module_data_out[1] ,
    \sw_294_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_295 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_295_module_data_in[7] ,
    \sw_295_module_data_in[6] ,
    \sw_295_module_data_in[5] ,
    \sw_295_module_data_in[4] ,
    \sw_295_module_data_in[3] ,
    \sw_295_module_data_in[2] ,
    \sw_295_module_data_in[1] ,
    \sw_295_module_data_in[0] }),
    .io_out({\sw_295_module_data_out[7] ,
    \sw_295_module_data_out[6] ,
    \sw_295_module_data_out[5] ,
    \sw_295_module_data_out[4] ,
    \sw_295_module_data_out[3] ,
    \sw_295_module_data_out[2] ,
    \sw_295_module_data_out[1] ,
    \sw_295_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_296 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_296_module_data_in[7] ,
    \sw_296_module_data_in[6] ,
    \sw_296_module_data_in[5] ,
    \sw_296_module_data_in[4] ,
    \sw_296_module_data_in[3] ,
    \sw_296_module_data_in[2] ,
    \sw_296_module_data_in[1] ,
    \sw_296_module_data_in[0] }),
    .io_out({\sw_296_module_data_out[7] ,
    \sw_296_module_data_out[6] ,
    \sw_296_module_data_out[5] ,
    \sw_296_module_data_out[4] ,
    \sw_296_module_data_out[3] ,
    \sw_296_module_data_out[2] ,
    \sw_296_module_data_out[1] ,
    \sw_296_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_297 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_297_module_data_in[7] ,
    \sw_297_module_data_in[6] ,
    \sw_297_module_data_in[5] ,
    \sw_297_module_data_in[4] ,
    \sw_297_module_data_in[3] ,
    \sw_297_module_data_in[2] ,
    \sw_297_module_data_in[1] ,
    \sw_297_module_data_in[0] }),
    .io_out({\sw_297_module_data_out[7] ,
    \sw_297_module_data_out[6] ,
    \sw_297_module_data_out[5] ,
    \sw_297_module_data_out[4] ,
    \sw_297_module_data_out[3] ,
    \sw_297_module_data_out[2] ,
    \sw_297_module_data_out[1] ,
    \sw_297_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_298 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_298_module_data_in[7] ,
    \sw_298_module_data_in[6] ,
    \sw_298_module_data_in[5] ,
    \sw_298_module_data_in[4] ,
    \sw_298_module_data_in[3] ,
    \sw_298_module_data_in[2] ,
    \sw_298_module_data_in[1] ,
    \sw_298_module_data_in[0] }),
    .io_out({\sw_298_module_data_out[7] ,
    \sw_298_module_data_out[6] ,
    \sw_298_module_data_out[5] ,
    \sw_298_module_data_out[4] ,
    \sw_298_module_data_out[3] ,
    \sw_298_module_data_out[2] ,
    \sw_298_module_data_out[1] ,
    \sw_298_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_299 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_299_module_data_in[7] ,
    \sw_299_module_data_in[6] ,
    \sw_299_module_data_in[5] ,
    \sw_299_module_data_in[4] ,
    \sw_299_module_data_in[3] ,
    \sw_299_module_data_in[2] ,
    \sw_299_module_data_in[1] ,
    \sw_299_module_data_in[0] }),
    .io_out({\sw_299_module_data_out[7] ,
    \sw_299_module_data_out[6] ,
    \sw_299_module_data_out[5] ,
    \sw_299_module_data_out[4] ,
    \sw_299_module_data_out[3] ,
    \sw_299_module_data_out[2] ,
    \sw_299_module_data_out[1] ,
    \sw_299_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_30 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_030_module_data_in[7] ,
    \sw_030_module_data_in[6] ,
    \sw_030_module_data_in[5] ,
    \sw_030_module_data_in[4] ,
    \sw_030_module_data_in[3] ,
    \sw_030_module_data_in[2] ,
    \sw_030_module_data_in[1] ,
    \sw_030_module_data_in[0] }),
    .io_out({\sw_030_module_data_out[7] ,
    \sw_030_module_data_out[6] ,
    \sw_030_module_data_out[5] ,
    \sw_030_module_data_out[4] ,
    \sw_030_module_data_out[3] ,
    \sw_030_module_data_out[2] ,
    \sw_030_module_data_out[1] ,
    \sw_030_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_300 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_300_module_data_in[7] ,
    \sw_300_module_data_in[6] ,
    \sw_300_module_data_in[5] ,
    \sw_300_module_data_in[4] ,
    \sw_300_module_data_in[3] ,
    \sw_300_module_data_in[2] ,
    \sw_300_module_data_in[1] ,
    \sw_300_module_data_in[0] }),
    .io_out({\sw_300_module_data_out[7] ,
    \sw_300_module_data_out[6] ,
    \sw_300_module_data_out[5] ,
    \sw_300_module_data_out[4] ,
    \sw_300_module_data_out[3] ,
    \sw_300_module_data_out[2] ,
    \sw_300_module_data_out[1] ,
    \sw_300_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_301 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_301_module_data_in[7] ,
    \sw_301_module_data_in[6] ,
    \sw_301_module_data_in[5] ,
    \sw_301_module_data_in[4] ,
    \sw_301_module_data_in[3] ,
    \sw_301_module_data_in[2] ,
    \sw_301_module_data_in[1] ,
    \sw_301_module_data_in[0] }),
    .io_out({\sw_301_module_data_out[7] ,
    \sw_301_module_data_out[6] ,
    \sw_301_module_data_out[5] ,
    \sw_301_module_data_out[4] ,
    \sw_301_module_data_out[3] ,
    \sw_301_module_data_out[2] ,
    \sw_301_module_data_out[1] ,
    \sw_301_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_302 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_302_module_data_in[7] ,
    \sw_302_module_data_in[6] ,
    \sw_302_module_data_in[5] ,
    \sw_302_module_data_in[4] ,
    \sw_302_module_data_in[3] ,
    \sw_302_module_data_in[2] ,
    \sw_302_module_data_in[1] ,
    \sw_302_module_data_in[0] }),
    .io_out({\sw_302_module_data_out[7] ,
    \sw_302_module_data_out[6] ,
    \sw_302_module_data_out[5] ,
    \sw_302_module_data_out[4] ,
    \sw_302_module_data_out[3] ,
    \sw_302_module_data_out[2] ,
    \sw_302_module_data_out[1] ,
    \sw_302_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_303 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_303_module_data_in[7] ,
    \sw_303_module_data_in[6] ,
    \sw_303_module_data_in[5] ,
    \sw_303_module_data_in[4] ,
    \sw_303_module_data_in[3] ,
    \sw_303_module_data_in[2] ,
    \sw_303_module_data_in[1] ,
    \sw_303_module_data_in[0] }),
    .io_out({\sw_303_module_data_out[7] ,
    \sw_303_module_data_out[6] ,
    \sw_303_module_data_out[5] ,
    \sw_303_module_data_out[4] ,
    \sw_303_module_data_out[3] ,
    \sw_303_module_data_out[2] ,
    \sw_303_module_data_out[1] ,
    \sw_303_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_304 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_304_module_data_in[7] ,
    \sw_304_module_data_in[6] ,
    \sw_304_module_data_in[5] ,
    \sw_304_module_data_in[4] ,
    \sw_304_module_data_in[3] ,
    \sw_304_module_data_in[2] ,
    \sw_304_module_data_in[1] ,
    \sw_304_module_data_in[0] }),
    .io_out({\sw_304_module_data_out[7] ,
    \sw_304_module_data_out[6] ,
    \sw_304_module_data_out[5] ,
    \sw_304_module_data_out[4] ,
    \sw_304_module_data_out[3] ,
    \sw_304_module_data_out[2] ,
    \sw_304_module_data_out[1] ,
    \sw_304_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_305 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_305_module_data_in[7] ,
    \sw_305_module_data_in[6] ,
    \sw_305_module_data_in[5] ,
    \sw_305_module_data_in[4] ,
    \sw_305_module_data_in[3] ,
    \sw_305_module_data_in[2] ,
    \sw_305_module_data_in[1] ,
    \sw_305_module_data_in[0] }),
    .io_out({\sw_305_module_data_out[7] ,
    \sw_305_module_data_out[6] ,
    \sw_305_module_data_out[5] ,
    \sw_305_module_data_out[4] ,
    \sw_305_module_data_out[3] ,
    \sw_305_module_data_out[2] ,
    \sw_305_module_data_out[1] ,
    \sw_305_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_306 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_306_module_data_in[7] ,
    \sw_306_module_data_in[6] ,
    \sw_306_module_data_in[5] ,
    \sw_306_module_data_in[4] ,
    \sw_306_module_data_in[3] ,
    \sw_306_module_data_in[2] ,
    \sw_306_module_data_in[1] ,
    \sw_306_module_data_in[0] }),
    .io_out({\sw_306_module_data_out[7] ,
    \sw_306_module_data_out[6] ,
    \sw_306_module_data_out[5] ,
    \sw_306_module_data_out[4] ,
    \sw_306_module_data_out[3] ,
    \sw_306_module_data_out[2] ,
    \sw_306_module_data_out[1] ,
    \sw_306_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_307 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_307_module_data_in[7] ,
    \sw_307_module_data_in[6] ,
    \sw_307_module_data_in[5] ,
    \sw_307_module_data_in[4] ,
    \sw_307_module_data_in[3] ,
    \sw_307_module_data_in[2] ,
    \sw_307_module_data_in[1] ,
    \sw_307_module_data_in[0] }),
    .io_out({\sw_307_module_data_out[7] ,
    \sw_307_module_data_out[6] ,
    \sw_307_module_data_out[5] ,
    \sw_307_module_data_out[4] ,
    \sw_307_module_data_out[3] ,
    \sw_307_module_data_out[2] ,
    \sw_307_module_data_out[1] ,
    \sw_307_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_308 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_308_module_data_in[7] ,
    \sw_308_module_data_in[6] ,
    \sw_308_module_data_in[5] ,
    \sw_308_module_data_in[4] ,
    \sw_308_module_data_in[3] ,
    \sw_308_module_data_in[2] ,
    \sw_308_module_data_in[1] ,
    \sw_308_module_data_in[0] }),
    .io_out({\sw_308_module_data_out[7] ,
    \sw_308_module_data_out[6] ,
    \sw_308_module_data_out[5] ,
    \sw_308_module_data_out[4] ,
    \sw_308_module_data_out[3] ,
    \sw_308_module_data_out[2] ,
    \sw_308_module_data_out[1] ,
    \sw_308_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_309 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_309_module_data_in[7] ,
    \sw_309_module_data_in[6] ,
    \sw_309_module_data_in[5] ,
    \sw_309_module_data_in[4] ,
    \sw_309_module_data_in[3] ,
    \sw_309_module_data_in[2] ,
    \sw_309_module_data_in[1] ,
    \sw_309_module_data_in[0] }),
    .io_out({\sw_309_module_data_out[7] ,
    \sw_309_module_data_out[6] ,
    \sw_309_module_data_out[5] ,
    \sw_309_module_data_out[4] ,
    \sw_309_module_data_out[3] ,
    \sw_309_module_data_out[2] ,
    \sw_309_module_data_out[1] ,
    \sw_309_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_31 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_031_module_data_in[7] ,
    \sw_031_module_data_in[6] ,
    \sw_031_module_data_in[5] ,
    \sw_031_module_data_in[4] ,
    \sw_031_module_data_in[3] ,
    \sw_031_module_data_in[2] ,
    \sw_031_module_data_in[1] ,
    \sw_031_module_data_in[0] }),
    .io_out({\sw_031_module_data_out[7] ,
    \sw_031_module_data_out[6] ,
    \sw_031_module_data_out[5] ,
    \sw_031_module_data_out[4] ,
    \sw_031_module_data_out[3] ,
    \sw_031_module_data_out[2] ,
    \sw_031_module_data_out[1] ,
    \sw_031_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_310 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_310_module_data_in[7] ,
    \sw_310_module_data_in[6] ,
    \sw_310_module_data_in[5] ,
    \sw_310_module_data_in[4] ,
    \sw_310_module_data_in[3] ,
    \sw_310_module_data_in[2] ,
    \sw_310_module_data_in[1] ,
    \sw_310_module_data_in[0] }),
    .io_out({\sw_310_module_data_out[7] ,
    \sw_310_module_data_out[6] ,
    \sw_310_module_data_out[5] ,
    \sw_310_module_data_out[4] ,
    \sw_310_module_data_out[3] ,
    \sw_310_module_data_out[2] ,
    \sw_310_module_data_out[1] ,
    \sw_310_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_311 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_311_module_data_in[7] ,
    \sw_311_module_data_in[6] ,
    \sw_311_module_data_in[5] ,
    \sw_311_module_data_in[4] ,
    \sw_311_module_data_in[3] ,
    \sw_311_module_data_in[2] ,
    \sw_311_module_data_in[1] ,
    \sw_311_module_data_in[0] }),
    .io_out({\sw_311_module_data_out[7] ,
    \sw_311_module_data_out[6] ,
    \sw_311_module_data_out[5] ,
    \sw_311_module_data_out[4] ,
    \sw_311_module_data_out[3] ,
    \sw_311_module_data_out[2] ,
    \sw_311_module_data_out[1] ,
    \sw_311_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_312 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_312_module_data_in[7] ,
    \sw_312_module_data_in[6] ,
    \sw_312_module_data_in[5] ,
    \sw_312_module_data_in[4] ,
    \sw_312_module_data_in[3] ,
    \sw_312_module_data_in[2] ,
    \sw_312_module_data_in[1] ,
    \sw_312_module_data_in[0] }),
    .io_out({\sw_312_module_data_out[7] ,
    \sw_312_module_data_out[6] ,
    \sw_312_module_data_out[5] ,
    \sw_312_module_data_out[4] ,
    \sw_312_module_data_out[3] ,
    \sw_312_module_data_out[2] ,
    \sw_312_module_data_out[1] ,
    \sw_312_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_313 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_313_module_data_in[7] ,
    \sw_313_module_data_in[6] ,
    \sw_313_module_data_in[5] ,
    \sw_313_module_data_in[4] ,
    \sw_313_module_data_in[3] ,
    \sw_313_module_data_in[2] ,
    \sw_313_module_data_in[1] ,
    \sw_313_module_data_in[0] }),
    .io_out({\sw_313_module_data_out[7] ,
    \sw_313_module_data_out[6] ,
    \sw_313_module_data_out[5] ,
    \sw_313_module_data_out[4] ,
    \sw_313_module_data_out[3] ,
    \sw_313_module_data_out[2] ,
    \sw_313_module_data_out[1] ,
    \sw_313_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_314 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_314_module_data_in[7] ,
    \sw_314_module_data_in[6] ,
    \sw_314_module_data_in[5] ,
    \sw_314_module_data_in[4] ,
    \sw_314_module_data_in[3] ,
    \sw_314_module_data_in[2] ,
    \sw_314_module_data_in[1] ,
    \sw_314_module_data_in[0] }),
    .io_out({\sw_314_module_data_out[7] ,
    \sw_314_module_data_out[6] ,
    \sw_314_module_data_out[5] ,
    \sw_314_module_data_out[4] ,
    \sw_314_module_data_out[3] ,
    \sw_314_module_data_out[2] ,
    \sw_314_module_data_out[1] ,
    \sw_314_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_315 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_315_module_data_in[7] ,
    \sw_315_module_data_in[6] ,
    \sw_315_module_data_in[5] ,
    \sw_315_module_data_in[4] ,
    \sw_315_module_data_in[3] ,
    \sw_315_module_data_in[2] ,
    \sw_315_module_data_in[1] ,
    \sw_315_module_data_in[0] }),
    .io_out({\sw_315_module_data_out[7] ,
    \sw_315_module_data_out[6] ,
    \sw_315_module_data_out[5] ,
    \sw_315_module_data_out[4] ,
    \sw_315_module_data_out[3] ,
    \sw_315_module_data_out[2] ,
    \sw_315_module_data_out[1] ,
    \sw_315_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_316 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_316_module_data_in[7] ,
    \sw_316_module_data_in[6] ,
    \sw_316_module_data_in[5] ,
    \sw_316_module_data_in[4] ,
    \sw_316_module_data_in[3] ,
    \sw_316_module_data_in[2] ,
    \sw_316_module_data_in[1] ,
    \sw_316_module_data_in[0] }),
    .io_out({\sw_316_module_data_out[7] ,
    \sw_316_module_data_out[6] ,
    \sw_316_module_data_out[5] ,
    \sw_316_module_data_out[4] ,
    \sw_316_module_data_out[3] ,
    \sw_316_module_data_out[2] ,
    \sw_316_module_data_out[1] ,
    \sw_316_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_317 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_317_module_data_in[7] ,
    \sw_317_module_data_in[6] ,
    \sw_317_module_data_in[5] ,
    \sw_317_module_data_in[4] ,
    \sw_317_module_data_in[3] ,
    \sw_317_module_data_in[2] ,
    \sw_317_module_data_in[1] ,
    \sw_317_module_data_in[0] }),
    .io_out({\sw_317_module_data_out[7] ,
    \sw_317_module_data_out[6] ,
    \sw_317_module_data_out[5] ,
    \sw_317_module_data_out[4] ,
    \sw_317_module_data_out[3] ,
    \sw_317_module_data_out[2] ,
    \sw_317_module_data_out[1] ,
    \sw_317_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_318 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_318_module_data_in[7] ,
    \sw_318_module_data_in[6] ,
    \sw_318_module_data_in[5] ,
    \sw_318_module_data_in[4] ,
    \sw_318_module_data_in[3] ,
    \sw_318_module_data_in[2] ,
    \sw_318_module_data_in[1] ,
    \sw_318_module_data_in[0] }),
    .io_out({\sw_318_module_data_out[7] ,
    \sw_318_module_data_out[6] ,
    \sw_318_module_data_out[5] ,
    \sw_318_module_data_out[4] ,
    \sw_318_module_data_out[3] ,
    \sw_318_module_data_out[2] ,
    \sw_318_module_data_out[1] ,
    \sw_318_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_319 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_319_module_data_in[7] ,
    \sw_319_module_data_in[6] ,
    \sw_319_module_data_in[5] ,
    \sw_319_module_data_in[4] ,
    \sw_319_module_data_in[3] ,
    \sw_319_module_data_in[2] ,
    \sw_319_module_data_in[1] ,
    \sw_319_module_data_in[0] }),
    .io_out({\sw_319_module_data_out[7] ,
    \sw_319_module_data_out[6] ,
    \sw_319_module_data_out[5] ,
    \sw_319_module_data_out[4] ,
    \sw_319_module_data_out[3] ,
    \sw_319_module_data_out[2] ,
    \sw_319_module_data_out[1] ,
    \sw_319_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_32 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_032_module_data_in[7] ,
    \sw_032_module_data_in[6] ,
    \sw_032_module_data_in[5] ,
    \sw_032_module_data_in[4] ,
    \sw_032_module_data_in[3] ,
    \sw_032_module_data_in[2] ,
    \sw_032_module_data_in[1] ,
    \sw_032_module_data_in[0] }),
    .io_out({\sw_032_module_data_out[7] ,
    \sw_032_module_data_out[6] ,
    \sw_032_module_data_out[5] ,
    \sw_032_module_data_out[4] ,
    \sw_032_module_data_out[3] ,
    \sw_032_module_data_out[2] ,
    \sw_032_module_data_out[1] ,
    \sw_032_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_320 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_320_module_data_in[7] ,
    \sw_320_module_data_in[6] ,
    \sw_320_module_data_in[5] ,
    \sw_320_module_data_in[4] ,
    \sw_320_module_data_in[3] ,
    \sw_320_module_data_in[2] ,
    \sw_320_module_data_in[1] ,
    \sw_320_module_data_in[0] }),
    .io_out({\sw_320_module_data_out[7] ,
    \sw_320_module_data_out[6] ,
    \sw_320_module_data_out[5] ,
    \sw_320_module_data_out[4] ,
    \sw_320_module_data_out[3] ,
    \sw_320_module_data_out[2] ,
    \sw_320_module_data_out[1] ,
    \sw_320_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_321 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_321_module_data_in[7] ,
    \sw_321_module_data_in[6] ,
    \sw_321_module_data_in[5] ,
    \sw_321_module_data_in[4] ,
    \sw_321_module_data_in[3] ,
    \sw_321_module_data_in[2] ,
    \sw_321_module_data_in[1] ,
    \sw_321_module_data_in[0] }),
    .io_out({\sw_321_module_data_out[7] ,
    \sw_321_module_data_out[6] ,
    \sw_321_module_data_out[5] ,
    \sw_321_module_data_out[4] ,
    \sw_321_module_data_out[3] ,
    \sw_321_module_data_out[2] ,
    \sw_321_module_data_out[1] ,
    \sw_321_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_322 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_322_module_data_in[7] ,
    \sw_322_module_data_in[6] ,
    \sw_322_module_data_in[5] ,
    \sw_322_module_data_in[4] ,
    \sw_322_module_data_in[3] ,
    \sw_322_module_data_in[2] ,
    \sw_322_module_data_in[1] ,
    \sw_322_module_data_in[0] }),
    .io_out({\sw_322_module_data_out[7] ,
    \sw_322_module_data_out[6] ,
    \sw_322_module_data_out[5] ,
    \sw_322_module_data_out[4] ,
    \sw_322_module_data_out[3] ,
    \sw_322_module_data_out[2] ,
    \sw_322_module_data_out[1] ,
    \sw_322_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_323 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_323_module_data_in[7] ,
    \sw_323_module_data_in[6] ,
    \sw_323_module_data_in[5] ,
    \sw_323_module_data_in[4] ,
    \sw_323_module_data_in[3] ,
    \sw_323_module_data_in[2] ,
    \sw_323_module_data_in[1] ,
    \sw_323_module_data_in[0] }),
    .io_out({\sw_323_module_data_out[7] ,
    \sw_323_module_data_out[6] ,
    \sw_323_module_data_out[5] ,
    \sw_323_module_data_out[4] ,
    \sw_323_module_data_out[3] ,
    \sw_323_module_data_out[2] ,
    \sw_323_module_data_out[1] ,
    \sw_323_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_324 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_324_module_data_in[7] ,
    \sw_324_module_data_in[6] ,
    \sw_324_module_data_in[5] ,
    \sw_324_module_data_in[4] ,
    \sw_324_module_data_in[3] ,
    \sw_324_module_data_in[2] ,
    \sw_324_module_data_in[1] ,
    \sw_324_module_data_in[0] }),
    .io_out({\sw_324_module_data_out[7] ,
    \sw_324_module_data_out[6] ,
    \sw_324_module_data_out[5] ,
    \sw_324_module_data_out[4] ,
    \sw_324_module_data_out[3] ,
    \sw_324_module_data_out[2] ,
    \sw_324_module_data_out[1] ,
    \sw_324_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_325 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_325_module_data_in[7] ,
    \sw_325_module_data_in[6] ,
    \sw_325_module_data_in[5] ,
    \sw_325_module_data_in[4] ,
    \sw_325_module_data_in[3] ,
    \sw_325_module_data_in[2] ,
    \sw_325_module_data_in[1] ,
    \sw_325_module_data_in[0] }),
    .io_out({\sw_325_module_data_out[7] ,
    \sw_325_module_data_out[6] ,
    \sw_325_module_data_out[5] ,
    \sw_325_module_data_out[4] ,
    \sw_325_module_data_out[3] ,
    \sw_325_module_data_out[2] ,
    \sw_325_module_data_out[1] ,
    \sw_325_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_326 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_326_module_data_in[7] ,
    \sw_326_module_data_in[6] ,
    \sw_326_module_data_in[5] ,
    \sw_326_module_data_in[4] ,
    \sw_326_module_data_in[3] ,
    \sw_326_module_data_in[2] ,
    \sw_326_module_data_in[1] ,
    \sw_326_module_data_in[0] }),
    .io_out({\sw_326_module_data_out[7] ,
    \sw_326_module_data_out[6] ,
    \sw_326_module_data_out[5] ,
    \sw_326_module_data_out[4] ,
    \sw_326_module_data_out[3] ,
    \sw_326_module_data_out[2] ,
    \sw_326_module_data_out[1] ,
    \sw_326_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_327 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_327_module_data_in[7] ,
    \sw_327_module_data_in[6] ,
    \sw_327_module_data_in[5] ,
    \sw_327_module_data_in[4] ,
    \sw_327_module_data_in[3] ,
    \sw_327_module_data_in[2] ,
    \sw_327_module_data_in[1] ,
    \sw_327_module_data_in[0] }),
    .io_out({\sw_327_module_data_out[7] ,
    \sw_327_module_data_out[6] ,
    \sw_327_module_data_out[5] ,
    \sw_327_module_data_out[4] ,
    \sw_327_module_data_out[3] ,
    \sw_327_module_data_out[2] ,
    \sw_327_module_data_out[1] ,
    \sw_327_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_328 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_328_module_data_in[7] ,
    \sw_328_module_data_in[6] ,
    \sw_328_module_data_in[5] ,
    \sw_328_module_data_in[4] ,
    \sw_328_module_data_in[3] ,
    \sw_328_module_data_in[2] ,
    \sw_328_module_data_in[1] ,
    \sw_328_module_data_in[0] }),
    .io_out({\sw_328_module_data_out[7] ,
    \sw_328_module_data_out[6] ,
    \sw_328_module_data_out[5] ,
    \sw_328_module_data_out[4] ,
    \sw_328_module_data_out[3] ,
    \sw_328_module_data_out[2] ,
    \sw_328_module_data_out[1] ,
    \sw_328_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_329 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_329_module_data_in[7] ,
    \sw_329_module_data_in[6] ,
    \sw_329_module_data_in[5] ,
    \sw_329_module_data_in[4] ,
    \sw_329_module_data_in[3] ,
    \sw_329_module_data_in[2] ,
    \sw_329_module_data_in[1] ,
    \sw_329_module_data_in[0] }),
    .io_out({\sw_329_module_data_out[7] ,
    \sw_329_module_data_out[6] ,
    \sw_329_module_data_out[5] ,
    \sw_329_module_data_out[4] ,
    \sw_329_module_data_out[3] ,
    \sw_329_module_data_out[2] ,
    \sw_329_module_data_out[1] ,
    \sw_329_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_33 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_033_module_data_in[7] ,
    \sw_033_module_data_in[6] ,
    \sw_033_module_data_in[5] ,
    \sw_033_module_data_in[4] ,
    \sw_033_module_data_in[3] ,
    \sw_033_module_data_in[2] ,
    \sw_033_module_data_in[1] ,
    \sw_033_module_data_in[0] }),
    .io_out({\sw_033_module_data_out[7] ,
    \sw_033_module_data_out[6] ,
    \sw_033_module_data_out[5] ,
    \sw_033_module_data_out[4] ,
    \sw_033_module_data_out[3] ,
    \sw_033_module_data_out[2] ,
    \sw_033_module_data_out[1] ,
    \sw_033_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_330 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_330_module_data_in[7] ,
    \sw_330_module_data_in[6] ,
    \sw_330_module_data_in[5] ,
    \sw_330_module_data_in[4] ,
    \sw_330_module_data_in[3] ,
    \sw_330_module_data_in[2] ,
    \sw_330_module_data_in[1] ,
    \sw_330_module_data_in[0] }),
    .io_out({\sw_330_module_data_out[7] ,
    \sw_330_module_data_out[6] ,
    \sw_330_module_data_out[5] ,
    \sw_330_module_data_out[4] ,
    \sw_330_module_data_out[3] ,
    \sw_330_module_data_out[2] ,
    \sw_330_module_data_out[1] ,
    \sw_330_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_331 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_331_module_data_in[7] ,
    \sw_331_module_data_in[6] ,
    \sw_331_module_data_in[5] ,
    \sw_331_module_data_in[4] ,
    \sw_331_module_data_in[3] ,
    \sw_331_module_data_in[2] ,
    \sw_331_module_data_in[1] ,
    \sw_331_module_data_in[0] }),
    .io_out({\sw_331_module_data_out[7] ,
    \sw_331_module_data_out[6] ,
    \sw_331_module_data_out[5] ,
    \sw_331_module_data_out[4] ,
    \sw_331_module_data_out[3] ,
    \sw_331_module_data_out[2] ,
    \sw_331_module_data_out[1] ,
    \sw_331_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_332 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_332_module_data_in[7] ,
    \sw_332_module_data_in[6] ,
    \sw_332_module_data_in[5] ,
    \sw_332_module_data_in[4] ,
    \sw_332_module_data_in[3] ,
    \sw_332_module_data_in[2] ,
    \sw_332_module_data_in[1] ,
    \sw_332_module_data_in[0] }),
    .io_out({\sw_332_module_data_out[7] ,
    \sw_332_module_data_out[6] ,
    \sw_332_module_data_out[5] ,
    \sw_332_module_data_out[4] ,
    \sw_332_module_data_out[3] ,
    \sw_332_module_data_out[2] ,
    \sw_332_module_data_out[1] ,
    \sw_332_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_333 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_333_module_data_in[7] ,
    \sw_333_module_data_in[6] ,
    \sw_333_module_data_in[5] ,
    \sw_333_module_data_in[4] ,
    \sw_333_module_data_in[3] ,
    \sw_333_module_data_in[2] ,
    \sw_333_module_data_in[1] ,
    \sw_333_module_data_in[0] }),
    .io_out({\sw_333_module_data_out[7] ,
    \sw_333_module_data_out[6] ,
    \sw_333_module_data_out[5] ,
    \sw_333_module_data_out[4] ,
    \sw_333_module_data_out[3] ,
    \sw_333_module_data_out[2] ,
    \sw_333_module_data_out[1] ,
    \sw_333_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_334 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_334_module_data_in[7] ,
    \sw_334_module_data_in[6] ,
    \sw_334_module_data_in[5] ,
    \sw_334_module_data_in[4] ,
    \sw_334_module_data_in[3] ,
    \sw_334_module_data_in[2] ,
    \sw_334_module_data_in[1] ,
    \sw_334_module_data_in[0] }),
    .io_out({\sw_334_module_data_out[7] ,
    \sw_334_module_data_out[6] ,
    \sw_334_module_data_out[5] ,
    \sw_334_module_data_out[4] ,
    \sw_334_module_data_out[3] ,
    \sw_334_module_data_out[2] ,
    \sw_334_module_data_out[1] ,
    \sw_334_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_335 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_335_module_data_in[7] ,
    \sw_335_module_data_in[6] ,
    \sw_335_module_data_in[5] ,
    \sw_335_module_data_in[4] ,
    \sw_335_module_data_in[3] ,
    \sw_335_module_data_in[2] ,
    \sw_335_module_data_in[1] ,
    \sw_335_module_data_in[0] }),
    .io_out({\sw_335_module_data_out[7] ,
    \sw_335_module_data_out[6] ,
    \sw_335_module_data_out[5] ,
    \sw_335_module_data_out[4] ,
    \sw_335_module_data_out[3] ,
    \sw_335_module_data_out[2] ,
    \sw_335_module_data_out[1] ,
    \sw_335_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_336 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_336_module_data_in[7] ,
    \sw_336_module_data_in[6] ,
    \sw_336_module_data_in[5] ,
    \sw_336_module_data_in[4] ,
    \sw_336_module_data_in[3] ,
    \sw_336_module_data_in[2] ,
    \sw_336_module_data_in[1] ,
    \sw_336_module_data_in[0] }),
    .io_out({\sw_336_module_data_out[7] ,
    \sw_336_module_data_out[6] ,
    \sw_336_module_data_out[5] ,
    \sw_336_module_data_out[4] ,
    \sw_336_module_data_out[3] ,
    \sw_336_module_data_out[2] ,
    \sw_336_module_data_out[1] ,
    \sw_336_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_337 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_337_module_data_in[7] ,
    \sw_337_module_data_in[6] ,
    \sw_337_module_data_in[5] ,
    \sw_337_module_data_in[4] ,
    \sw_337_module_data_in[3] ,
    \sw_337_module_data_in[2] ,
    \sw_337_module_data_in[1] ,
    \sw_337_module_data_in[0] }),
    .io_out({\sw_337_module_data_out[7] ,
    \sw_337_module_data_out[6] ,
    \sw_337_module_data_out[5] ,
    \sw_337_module_data_out[4] ,
    \sw_337_module_data_out[3] ,
    \sw_337_module_data_out[2] ,
    \sw_337_module_data_out[1] ,
    \sw_337_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_338 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_338_module_data_in[7] ,
    \sw_338_module_data_in[6] ,
    \sw_338_module_data_in[5] ,
    \sw_338_module_data_in[4] ,
    \sw_338_module_data_in[3] ,
    \sw_338_module_data_in[2] ,
    \sw_338_module_data_in[1] ,
    \sw_338_module_data_in[0] }),
    .io_out({\sw_338_module_data_out[7] ,
    \sw_338_module_data_out[6] ,
    \sw_338_module_data_out[5] ,
    \sw_338_module_data_out[4] ,
    \sw_338_module_data_out[3] ,
    \sw_338_module_data_out[2] ,
    \sw_338_module_data_out[1] ,
    \sw_338_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_339 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_339_module_data_in[7] ,
    \sw_339_module_data_in[6] ,
    \sw_339_module_data_in[5] ,
    \sw_339_module_data_in[4] ,
    \sw_339_module_data_in[3] ,
    \sw_339_module_data_in[2] ,
    \sw_339_module_data_in[1] ,
    \sw_339_module_data_in[0] }),
    .io_out({\sw_339_module_data_out[7] ,
    \sw_339_module_data_out[6] ,
    \sw_339_module_data_out[5] ,
    \sw_339_module_data_out[4] ,
    \sw_339_module_data_out[3] ,
    \sw_339_module_data_out[2] ,
    \sw_339_module_data_out[1] ,
    \sw_339_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_34 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_034_module_data_in[7] ,
    \sw_034_module_data_in[6] ,
    \sw_034_module_data_in[5] ,
    \sw_034_module_data_in[4] ,
    \sw_034_module_data_in[3] ,
    \sw_034_module_data_in[2] ,
    \sw_034_module_data_in[1] ,
    \sw_034_module_data_in[0] }),
    .io_out({\sw_034_module_data_out[7] ,
    \sw_034_module_data_out[6] ,
    \sw_034_module_data_out[5] ,
    \sw_034_module_data_out[4] ,
    \sw_034_module_data_out[3] ,
    \sw_034_module_data_out[2] ,
    \sw_034_module_data_out[1] ,
    \sw_034_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_340 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_340_module_data_in[7] ,
    \sw_340_module_data_in[6] ,
    \sw_340_module_data_in[5] ,
    \sw_340_module_data_in[4] ,
    \sw_340_module_data_in[3] ,
    \sw_340_module_data_in[2] ,
    \sw_340_module_data_in[1] ,
    \sw_340_module_data_in[0] }),
    .io_out({\sw_340_module_data_out[7] ,
    \sw_340_module_data_out[6] ,
    \sw_340_module_data_out[5] ,
    \sw_340_module_data_out[4] ,
    \sw_340_module_data_out[3] ,
    \sw_340_module_data_out[2] ,
    \sw_340_module_data_out[1] ,
    \sw_340_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_341 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_341_module_data_in[7] ,
    \sw_341_module_data_in[6] ,
    \sw_341_module_data_in[5] ,
    \sw_341_module_data_in[4] ,
    \sw_341_module_data_in[3] ,
    \sw_341_module_data_in[2] ,
    \sw_341_module_data_in[1] ,
    \sw_341_module_data_in[0] }),
    .io_out({\sw_341_module_data_out[7] ,
    \sw_341_module_data_out[6] ,
    \sw_341_module_data_out[5] ,
    \sw_341_module_data_out[4] ,
    \sw_341_module_data_out[3] ,
    \sw_341_module_data_out[2] ,
    \sw_341_module_data_out[1] ,
    \sw_341_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_342 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_342_module_data_in[7] ,
    \sw_342_module_data_in[6] ,
    \sw_342_module_data_in[5] ,
    \sw_342_module_data_in[4] ,
    \sw_342_module_data_in[3] ,
    \sw_342_module_data_in[2] ,
    \sw_342_module_data_in[1] ,
    \sw_342_module_data_in[0] }),
    .io_out({\sw_342_module_data_out[7] ,
    \sw_342_module_data_out[6] ,
    \sw_342_module_data_out[5] ,
    \sw_342_module_data_out[4] ,
    \sw_342_module_data_out[3] ,
    \sw_342_module_data_out[2] ,
    \sw_342_module_data_out[1] ,
    \sw_342_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_343 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_343_module_data_in[7] ,
    \sw_343_module_data_in[6] ,
    \sw_343_module_data_in[5] ,
    \sw_343_module_data_in[4] ,
    \sw_343_module_data_in[3] ,
    \sw_343_module_data_in[2] ,
    \sw_343_module_data_in[1] ,
    \sw_343_module_data_in[0] }),
    .io_out({\sw_343_module_data_out[7] ,
    \sw_343_module_data_out[6] ,
    \sw_343_module_data_out[5] ,
    \sw_343_module_data_out[4] ,
    \sw_343_module_data_out[3] ,
    \sw_343_module_data_out[2] ,
    \sw_343_module_data_out[1] ,
    \sw_343_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_344 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_344_module_data_in[7] ,
    \sw_344_module_data_in[6] ,
    \sw_344_module_data_in[5] ,
    \sw_344_module_data_in[4] ,
    \sw_344_module_data_in[3] ,
    \sw_344_module_data_in[2] ,
    \sw_344_module_data_in[1] ,
    \sw_344_module_data_in[0] }),
    .io_out({\sw_344_module_data_out[7] ,
    \sw_344_module_data_out[6] ,
    \sw_344_module_data_out[5] ,
    \sw_344_module_data_out[4] ,
    \sw_344_module_data_out[3] ,
    \sw_344_module_data_out[2] ,
    \sw_344_module_data_out[1] ,
    \sw_344_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_345 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_345_module_data_in[7] ,
    \sw_345_module_data_in[6] ,
    \sw_345_module_data_in[5] ,
    \sw_345_module_data_in[4] ,
    \sw_345_module_data_in[3] ,
    \sw_345_module_data_in[2] ,
    \sw_345_module_data_in[1] ,
    \sw_345_module_data_in[0] }),
    .io_out({\sw_345_module_data_out[7] ,
    \sw_345_module_data_out[6] ,
    \sw_345_module_data_out[5] ,
    \sw_345_module_data_out[4] ,
    \sw_345_module_data_out[3] ,
    \sw_345_module_data_out[2] ,
    \sw_345_module_data_out[1] ,
    \sw_345_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_346 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_346_module_data_in[7] ,
    \sw_346_module_data_in[6] ,
    \sw_346_module_data_in[5] ,
    \sw_346_module_data_in[4] ,
    \sw_346_module_data_in[3] ,
    \sw_346_module_data_in[2] ,
    \sw_346_module_data_in[1] ,
    \sw_346_module_data_in[0] }),
    .io_out({\sw_346_module_data_out[7] ,
    \sw_346_module_data_out[6] ,
    \sw_346_module_data_out[5] ,
    \sw_346_module_data_out[4] ,
    \sw_346_module_data_out[3] ,
    \sw_346_module_data_out[2] ,
    \sw_346_module_data_out[1] ,
    \sw_346_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_347 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_347_module_data_in[7] ,
    \sw_347_module_data_in[6] ,
    \sw_347_module_data_in[5] ,
    \sw_347_module_data_in[4] ,
    \sw_347_module_data_in[3] ,
    \sw_347_module_data_in[2] ,
    \sw_347_module_data_in[1] ,
    \sw_347_module_data_in[0] }),
    .io_out({\sw_347_module_data_out[7] ,
    \sw_347_module_data_out[6] ,
    \sw_347_module_data_out[5] ,
    \sw_347_module_data_out[4] ,
    \sw_347_module_data_out[3] ,
    \sw_347_module_data_out[2] ,
    \sw_347_module_data_out[1] ,
    \sw_347_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_348 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_348_module_data_in[7] ,
    \sw_348_module_data_in[6] ,
    \sw_348_module_data_in[5] ,
    \sw_348_module_data_in[4] ,
    \sw_348_module_data_in[3] ,
    \sw_348_module_data_in[2] ,
    \sw_348_module_data_in[1] ,
    \sw_348_module_data_in[0] }),
    .io_out({\sw_348_module_data_out[7] ,
    \sw_348_module_data_out[6] ,
    \sw_348_module_data_out[5] ,
    \sw_348_module_data_out[4] ,
    \sw_348_module_data_out[3] ,
    \sw_348_module_data_out[2] ,
    \sw_348_module_data_out[1] ,
    \sw_348_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_349 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_349_module_data_in[7] ,
    \sw_349_module_data_in[6] ,
    \sw_349_module_data_in[5] ,
    \sw_349_module_data_in[4] ,
    \sw_349_module_data_in[3] ,
    \sw_349_module_data_in[2] ,
    \sw_349_module_data_in[1] ,
    \sw_349_module_data_in[0] }),
    .io_out({\sw_349_module_data_out[7] ,
    \sw_349_module_data_out[6] ,
    \sw_349_module_data_out[5] ,
    \sw_349_module_data_out[4] ,
    \sw_349_module_data_out[3] ,
    \sw_349_module_data_out[2] ,
    \sw_349_module_data_out[1] ,
    \sw_349_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_35 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_035_module_data_in[7] ,
    \sw_035_module_data_in[6] ,
    \sw_035_module_data_in[5] ,
    \sw_035_module_data_in[4] ,
    \sw_035_module_data_in[3] ,
    \sw_035_module_data_in[2] ,
    \sw_035_module_data_in[1] ,
    \sw_035_module_data_in[0] }),
    .io_out({\sw_035_module_data_out[7] ,
    \sw_035_module_data_out[6] ,
    \sw_035_module_data_out[5] ,
    \sw_035_module_data_out[4] ,
    \sw_035_module_data_out[3] ,
    \sw_035_module_data_out[2] ,
    \sw_035_module_data_out[1] ,
    \sw_035_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_350 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_350_module_data_in[7] ,
    \sw_350_module_data_in[6] ,
    \sw_350_module_data_in[5] ,
    \sw_350_module_data_in[4] ,
    \sw_350_module_data_in[3] ,
    \sw_350_module_data_in[2] ,
    \sw_350_module_data_in[1] ,
    \sw_350_module_data_in[0] }),
    .io_out({\sw_350_module_data_out[7] ,
    \sw_350_module_data_out[6] ,
    \sw_350_module_data_out[5] ,
    \sw_350_module_data_out[4] ,
    \sw_350_module_data_out[3] ,
    \sw_350_module_data_out[2] ,
    \sw_350_module_data_out[1] ,
    \sw_350_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_351 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_351_module_data_in[7] ,
    \sw_351_module_data_in[6] ,
    \sw_351_module_data_in[5] ,
    \sw_351_module_data_in[4] ,
    \sw_351_module_data_in[3] ,
    \sw_351_module_data_in[2] ,
    \sw_351_module_data_in[1] ,
    \sw_351_module_data_in[0] }),
    .io_out({\sw_351_module_data_out[7] ,
    \sw_351_module_data_out[6] ,
    \sw_351_module_data_out[5] ,
    \sw_351_module_data_out[4] ,
    \sw_351_module_data_out[3] ,
    \sw_351_module_data_out[2] ,
    \sw_351_module_data_out[1] ,
    \sw_351_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_352 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_352_module_data_in[7] ,
    \sw_352_module_data_in[6] ,
    \sw_352_module_data_in[5] ,
    \sw_352_module_data_in[4] ,
    \sw_352_module_data_in[3] ,
    \sw_352_module_data_in[2] ,
    \sw_352_module_data_in[1] ,
    \sw_352_module_data_in[0] }),
    .io_out({\sw_352_module_data_out[7] ,
    \sw_352_module_data_out[6] ,
    \sw_352_module_data_out[5] ,
    \sw_352_module_data_out[4] ,
    \sw_352_module_data_out[3] ,
    \sw_352_module_data_out[2] ,
    \sw_352_module_data_out[1] ,
    \sw_352_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_353 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_353_module_data_in[7] ,
    \sw_353_module_data_in[6] ,
    \sw_353_module_data_in[5] ,
    \sw_353_module_data_in[4] ,
    \sw_353_module_data_in[3] ,
    \sw_353_module_data_in[2] ,
    \sw_353_module_data_in[1] ,
    \sw_353_module_data_in[0] }),
    .io_out({\sw_353_module_data_out[7] ,
    \sw_353_module_data_out[6] ,
    \sw_353_module_data_out[5] ,
    \sw_353_module_data_out[4] ,
    \sw_353_module_data_out[3] ,
    \sw_353_module_data_out[2] ,
    \sw_353_module_data_out[1] ,
    \sw_353_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_354 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_354_module_data_in[7] ,
    \sw_354_module_data_in[6] ,
    \sw_354_module_data_in[5] ,
    \sw_354_module_data_in[4] ,
    \sw_354_module_data_in[3] ,
    \sw_354_module_data_in[2] ,
    \sw_354_module_data_in[1] ,
    \sw_354_module_data_in[0] }),
    .io_out({\sw_354_module_data_out[7] ,
    \sw_354_module_data_out[6] ,
    \sw_354_module_data_out[5] ,
    \sw_354_module_data_out[4] ,
    \sw_354_module_data_out[3] ,
    \sw_354_module_data_out[2] ,
    \sw_354_module_data_out[1] ,
    \sw_354_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_355 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_355_module_data_in[7] ,
    \sw_355_module_data_in[6] ,
    \sw_355_module_data_in[5] ,
    \sw_355_module_data_in[4] ,
    \sw_355_module_data_in[3] ,
    \sw_355_module_data_in[2] ,
    \sw_355_module_data_in[1] ,
    \sw_355_module_data_in[0] }),
    .io_out({\sw_355_module_data_out[7] ,
    \sw_355_module_data_out[6] ,
    \sw_355_module_data_out[5] ,
    \sw_355_module_data_out[4] ,
    \sw_355_module_data_out[3] ,
    \sw_355_module_data_out[2] ,
    \sw_355_module_data_out[1] ,
    \sw_355_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_356 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_356_module_data_in[7] ,
    \sw_356_module_data_in[6] ,
    \sw_356_module_data_in[5] ,
    \sw_356_module_data_in[4] ,
    \sw_356_module_data_in[3] ,
    \sw_356_module_data_in[2] ,
    \sw_356_module_data_in[1] ,
    \sw_356_module_data_in[0] }),
    .io_out({\sw_356_module_data_out[7] ,
    \sw_356_module_data_out[6] ,
    \sw_356_module_data_out[5] ,
    \sw_356_module_data_out[4] ,
    \sw_356_module_data_out[3] ,
    \sw_356_module_data_out[2] ,
    \sw_356_module_data_out[1] ,
    \sw_356_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_357 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_357_module_data_in[7] ,
    \sw_357_module_data_in[6] ,
    \sw_357_module_data_in[5] ,
    \sw_357_module_data_in[4] ,
    \sw_357_module_data_in[3] ,
    \sw_357_module_data_in[2] ,
    \sw_357_module_data_in[1] ,
    \sw_357_module_data_in[0] }),
    .io_out({\sw_357_module_data_out[7] ,
    \sw_357_module_data_out[6] ,
    \sw_357_module_data_out[5] ,
    \sw_357_module_data_out[4] ,
    \sw_357_module_data_out[3] ,
    \sw_357_module_data_out[2] ,
    \sw_357_module_data_out[1] ,
    \sw_357_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_358 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_358_module_data_in[7] ,
    \sw_358_module_data_in[6] ,
    \sw_358_module_data_in[5] ,
    \sw_358_module_data_in[4] ,
    \sw_358_module_data_in[3] ,
    \sw_358_module_data_in[2] ,
    \sw_358_module_data_in[1] ,
    \sw_358_module_data_in[0] }),
    .io_out({\sw_358_module_data_out[7] ,
    \sw_358_module_data_out[6] ,
    \sw_358_module_data_out[5] ,
    \sw_358_module_data_out[4] ,
    \sw_358_module_data_out[3] ,
    \sw_358_module_data_out[2] ,
    \sw_358_module_data_out[1] ,
    \sw_358_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_359 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_359_module_data_in[7] ,
    \sw_359_module_data_in[6] ,
    \sw_359_module_data_in[5] ,
    \sw_359_module_data_in[4] ,
    \sw_359_module_data_in[3] ,
    \sw_359_module_data_in[2] ,
    \sw_359_module_data_in[1] ,
    \sw_359_module_data_in[0] }),
    .io_out({\sw_359_module_data_out[7] ,
    \sw_359_module_data_out[6] ,
    \sw_359_module_data_out[5] ,
    \sw_359_module_data_out[4] ,
    \sw_359_module_data_out[3] ,
    \sw_359_module_data_out[2] ,
    \sw_359_module_data_out[1] ,
    \sw_359_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_36 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_036_module_data_in[7] ,
    \sw_036_module_data_in[6] ,
    \sw_036_module_data_in[5] ,
    \sw_036_module_data_in[4] ,
    \sw_036_module_data_in[3] ,
    \sw_036_module_data_in[2] ,
    \sw_036_module_data_in[1] ,
    \sw_036_module_data_in[0] }),
    .io_out({\sw_036_module_data_out[7] ,
    \sw_036_module_data_out[6] ,
    \sw_036_module_data_out[5] ,
    \sw_036_module_data_out[4] ,
    \sw_036_module_data_out[3] ,
    \sw_036_module_data_out[2] ,
    \sw_036_module_data_out[1] ,
    \sw_036_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_360 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_360_module_data_in[7] ,
    \sw_360_module_data_in[6] ,
    \sw_360_module_data_in[5] ,
    \sw_360_module_data_in[4] ,
    \sw_360_module_data_in[3] ,
    \sw_360_module_data_in[2] ,
    \sw_360_module_data_in[1] ,
    \sw_360_module_data_in[0] }),
    .io_out({\sw_360_module_data_out[7] ,
    \sw_360_module_data_out[6] ,
    \sw_360_module_data_out[5] ,
    \sw_360_module_data_out[4] ,
    \sw_360_module_data_out[3] ,
    \sw_360_module_data_out[2] ,
    \sw_360_module_data_out[1] ,
    \sw_360_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_361 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_361_module_data_in[7] ,
    \sw_361_module_data_in[6] ,
    \sw_361_module_data_in[5] ,
    \sw_361_module_data_in[4] ,
    \sw_361_module_data_in[3] ,
    \sw_361_module_data_in[2] ,
    \sw_361_module_data_in[1] ,
    \sw_361_module_data_in[0] }),
    .io_out({\sw_361_module_data_out[7] ,
    \sw_361_module_data_out[6] ,
    \sw_361_module_data_out[5] ,
    \sw_361_module_data_out[4] ,
    \sw_361_module_data_out[3] ,
    \sw_361_module_data_out[2] ,
    \sw_361_module_data_out[1] ,
    \sw_361_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_362 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_362_module_data_in[7] ,
    \sw_362_module_data_in[6] ,
    \sw_362_module_data_in[5] ,
    \sw_362_module_data_in[4] ,
    \sw_362_module_data_in[3] ,
    \sw_362_module_data_in[2] ,
    \sw_362_module_data_in[1] ,
    \sw_362_module_data_in[0] }),
    .io_out({\sw_362_module_data_out[7] ,
    \sw_362_module_data_out[6] ,
    \sw_362_module_data_out[5] ,
    \sw_362_module_data_out[4] ,
    \sw_362_module_data_out[3] ,
    \sw_362_module_data_out[2] ,
    \sw_362_module_data_out[1] ,
    \sw_362_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_363 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_363_module_data_in[7] ,
    \sw_363_module_data_in[6] ,
    \sw_363_module_data_in[5] ,
    \sw_363_module_data_in[4] ,
    \sw_363_module_data_in[3] ,
    \sw_363_module_data_in[2] ,
    \sw_363_module_data_in[1] ,
    \sw_363_module_data_in[0] }),
    .io_out({\sw_363_module_data_out[7] ,
    \sw_363_module_data_out[6] ,
    \sw_363_module_data_out[5] ,
    \sw_363_module_data_out[4] ,
    \sw_363_module_data_out[3] ,
    \sw_363_module_data_out[2] ,
    \sw_363_module_data_out[1] ,
    \sw_363_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_364 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_364_module_data_in[7] ,
    \sw_364_module_data_in[6] ,
    \sw_364_module_data_in[5] ,
    \sw_364_module_data_in[4] ,
    \sw_364_module_data_in[3] ,
    \sw_364_module_data_in[2] ,
    \sw_364_module_data_in[1] ,
    \sw_364_module_data_in[0] }),
    .io_out({\sw_364_module_data_out[7] ,
    \sw_364_module_data_out[6] ,
    \sw_364_module_data_out[5] ,
    \sw_364_module_data_out[4] ,
    \sw_364_module_data_out[3] ,
    \sw_364_module_data_out[2] ,
    \sw_364_module_data_out[1] ,
    \sw_364_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_365 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_365_module_data_in[7] ,
    \sw_365_module_data_in[6] ,
    \sw_365_module_data_in[5] ,
    \sw_365_module_data_in[4] ,
    \sw_365_module_data_in[3] ,
    \sw_365_module_data_in[2] ,
    \sw_365_module_data_in[1] ,
    \sw_365_module_data_in[0] }),
    .io_out({\sw_365_module_data_out[7] ,
    \sw_365_module_data_out[6] ,
    \sw_365_module_data_out[5] ,
    \sw_365_module_data_out[4] ,
    \sw_365_module_data_out[3] ,
    \sw_365_module_data_out[2] ,
    \sw_365_module_data_out[1] ,
    \sw_365_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_366 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_366_module_data_in[7] ,
    \sw_366_module_data_in[6] ,
    \sw_366_module_data_in[5] ,
    \sw_366_module_data_in[4] ,
    \sw_366_module_data_in[3] ,
    \sw_366_module_data_in[2] ,
    \sw_366_module_data_in[1] ,
    \sw_366_module_data_in[0] }),
    .io_out({\sw_366_module_data_out[7] ,
    \sw_366_module_data_out[6] ,
    \sw_366_module_data_out[5] ,
    \sw_366_module_data_out[4] ,
    \sw_366_module_data_out[3] ,
    \sw_366_module_data_out[2] ,
    \sw_366_module_data_out[1] ,
    \sw_366_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_367 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_367_module_data_in[7] ,
    \sw_367_module_data_in[6] ,
    \sw_367_module_data_in[5] ,
    \sw_367_module_data_in[4] ,
    \sw_367_module_data_in[3] ,
    \sw_367_module_data_in[2] ,
    \sw_367_module_data_in[1] ,
    \sw_367_module_data_in[0] }),
    .io_out({\sw_367_module_data_out[7] ,
    \sw_367_module_data_out[6] ,
    \sw_367_module_data_out[5] ,
    \sw_367_module_data_out[4] ,
    \sw_367_module_data_out[3] ,
    \sw_367_module_data_out[2] ,
    \sw_367_module_data_out[1] ,
    \sw_367_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_368 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_368_module_data_in[7] ,
    \sw_368_module_data_in[6] ,
    \sw_368_module_data_in[5] ,
    \sw_368_module_data_in[4] ,
    \sw_368_module_data_in[3] ,
    \sw_368_module_data_in[2] ,
    \sw_368_module_data_in[1] ,
    \sw_368_module_data_in[0] }),
    .io_out({\sw_368_module_data_out[7] ,
    \sw_368_module_data_out[6] ,
    \sw_368_module_data_out[5] ,
    \sw_368_module_data_out[4] ,
    \sw_368_module_data_out[3] ,
    \sw_368_module_data_out[2] ,
    \sw_368_module_data_out[1] ,
    \sw_368_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_369 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_369_module_data_in[7] ,
    \sw_369_module_data_in[6] ,
    \sw_369_module_data_in[5] ,
    \sw_369_module_data_in[4] ,
    \sw_369_module_data_in[3] ,
    \sw_369_module_data_in[2] ,
    \sw_369_module_data_in[1] ,
    \sw_369_module_data_in[0] }),
    .io_out({\sw_369_module_data_out[7] ,
    \sw_369_module_data_out[6] ,
    \sw_369_module_data_out[5] ,
    \sw_369_module_data_out[4] ,
    \sw_369_module_data_out[3] ,
    \sw_369_module_data_out[2] ,
    \sw_369_module_data_out[1] ,
    \sw_369_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_37 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_037_module_data_in[7] ,
    \sw_037_module_data_in[6] ,
    \sw_037_module_data_in[5] ,
    \sw_037_module_data_in[4] ,
    \sw_037_module_data_in[3] ,
    \sw_037_module_data_in[2] ,
    \sw_037_module_data_in[1] ,
    \sw_037_module_data_in[0] }),
    .io_out({\sw_037_module_data_out[7] ,
    \sw_037_module_data_out[6] ,
    \sw_037_module_data_out[5] ,
    \sw_037_module_data_out[4] ,
    \sw_037_module_data_out[3] ,
    \sw_037_module_data_out[2] ,
    \sw_037_module_data_out[1] ,
    \sw_037_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_370 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_370_module_data_in[7] ,
    \sw_370_module_data_in[6] ,
    \sw_370_module_data_in[5] ,
    \sw_370_module_data_in[4] ,
    \sw_370_module_data_in[3] ,
    \sw_370_module_data_in[2] ,
    \sw_370_module_data_in[1] ,
    \sw_370_module_data_in[0] }),
    .io_out({\sw_370_module_data_out[7] ,
    \sw_370_module_data_out[6] ,
    \sw_370_module_data_out[5] ,
    \sw_370_module_data_out[4] ,
    \sw_370_module_data_out[3] ,
    \sw_370_module_data_out[2] ,
    \sw_370_module_data_out[1] ,
    \sw_370_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_371 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_371_module_data_in[7] ,
    \sw_371_module_data_in[6] ,
    \sw_371_module_data_in[5] ,
    \sw_371_module_data_in[4] ,
    \sw_371_module_data_in[3] ,
    \sw_371_module_data_in[2] ,
    \sw_371_module_data_in[1] ,
    \sw_371_module_data_in[0] }),
    .io_out({\sw_371_module_data_out[7] ,
    \sw_371_module_data_out[6] ,
    \sw_371_module_data_out[5] ,
    \sw_371_module_data_out[4] ,
    \sw_371_module_data_out[3] ,
    \sw_371_module_data_out[2] ,
    \sw_371_module_data_out[1] ,
    \sw_371_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_372 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_372_module_data_in[7] ,
    \sw_372_module_data_in[6] ,
    \sw_372_module_data_in[5] ,
    \sw_372_module_data_in[4] ,
    \sw_372_module_data_in[3] ,
    \sw_372_module_data_in[2] ,
    \sw_372_module_data_in[1] ,
    \sw_372_module_data_in[0] }),
    .io_out({\sw_372_module_data_out[7] ,
    \sw_372_module_data_out[6] ,
    \sw_372_module_data_out[5] ,
    \sw_372_module_data_out[4] ,
    \sw_372_module_data_out[3] ,
    \sw_372_module_data_out[2] ,
    \sw_372_module_data_out[1] ,
    \sw_372_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_373 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_373_module_data_in[7] ,
    \sw_373_module_data_in[6] ,
    \sw_373_module_data_in[5] ,
    \sw_373_module_data_in[4] ,
    \sw_373_module_data_in[3] ,
    \sw_373_module_data_in[2] ,
    \sw_373_module_data_in[1] ,
    \sw_373_module_data_in[0] }),
    .io_out({\sw_373_module_data_out[7] ,
    \sw_373_module_data_out[6] ,
    \sw_373_module_data_out[5] ,
    \sw_373_module_data_out[4] ,
    \sw_373_module_data_out[3] ,
    \sw_373_module_data_out[2] ,
    \sw_373_module_data_out[1] ,
    \sw_373_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_374 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_374_module_data_in[7] ,
    \sw_374_module_data_in[6] ,
    \sw_374_module_data_in[5] ,
    \sw_374_module_data_in[4] ,
    \sw_374_module_data_in[3] ,
    \sw_374_module_data_in[2] ,
    \sw_374_module_data_in[1] ,
    \sw_374_module_data_in[0] }),
    .io_out({\sw_374_module_data_out[7] ,
    \sw_374_module_data_out[6] ,
    \sw_374_module_data_out[5] ,
    \sw_374_module_data_out[4] ,
    \sw_374_module_data_out[3] ,
    \sw_374_module_data_out[2] ,
    \sw_374_module_data_out[1] ,
    \sw_374_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_375 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_375_module_data_in[7] ,
    \sw_375_module_data_in[6] ,
    \sw_375_module_data_in[5] ,
    \sw_375_module_data_in[4] ,
    \sw_375_module_data_in[3] ,
    \sw_375_module_data_in[2] ,
    \sw_375_module_data_in[1] ,
    \sw_375_module_data_in[0] }),
    .io_out({\sw_375_module_data_out[7] ,
    \sw_375_module_data_out[6] ,
    \sw_375_module_data_out[5] ,
    \sw_375_module_data_out[4] ,
    \sw_375_module_data_out[3] ,
    \sw_375_module_data_out[2] ,
    \sw_375_module_data_out[1] ,
    \sw_375_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_376 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_376_module_data_in[7] ,
    \sw_376_module_data_in[6] ,
    \sw_376_module_data_in[5] ,
    \sw_376_module_data_in[4] ,
    \sw_376_module_data_in[3] ,
    \sw_376_module_data_in[2] ,
    \sw_376_module_data_in[1] ,
    \sw_376_module_data_in[0] }),
    .io_out({\sw_376_module_data_out[7] ,
    \sw_376_module_data_out[6] ,
    \sw_376_module_data_out[5] ,
    \sw_376_module_data_out[4] ,
    \sw_376_module_data_out[3] ,
    \sw_376_module_data_out[2] ,
    \sw_376_module_data_out[1] ,
    \sw_376_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_377 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_377_module_data_in[7] ,
    \sw_377_module_data_in[6] ,
    \sw_377_module_data_in[5] ,
    \sw_377_module_data_in[4] ,
    \sw_377_module_data_in[3] ,
    \sw_377_module_data_in[2] ,
    \sw_377_module_data_in[1] ,
    \sw_377_module_data_in[0] }),
    .io_out({\sw_377_module_data_out[7] ,
    \sw_377_module_data_out[6] ,
    \sw_377_module_data_out[5] ,
    \sw_377_module_data_out[4] ,
    \sw_377_module_data_out[3] ,
    \sw_377_module_data_out[2] ,
    \sw_377_module_data_out[1] ,
    \sw_377_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_378 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_378_module_data_in[7] ,
    \sw_378_module_data_in[6] ,
    \sw_378_module_data_in[5] ,
    \sw_378_module_data_in[4] ,
    \sw_378_module_data_in[3] ,
    \sw_378_module_data_in[2] ,
    \sw_378_module_data_in[1] ,
    \sw_378_module_data_in[0] }),
    .io_out({\sw_378_module_data_out[7] ,
    \sw_378_module_data_out[6] ,
    \sw_378_module_data_out[5] ,
    \sw_378_module_data_out[4] ,
    \sw_378_module_data_out[3] ,
    \sw_378_module_data_out[2] ,
    \sw_378_module_data_out[1] ,
    \sw_378_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_379 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_379_module_data_in[7] ,
    \sw_379_module_data_in[6] ,
    \sw_379_module_data_in[5] ,
    \sw_379_module_data_in[4] ,
    \sw_379_module_data_in[3] ,
    \sw_379_module_data_in[2] ,
    \sw_379_module_data_in[1] ,
    \sw_379_module_data_in[0] }),
    .io_out({\sw_379_module_data_out[7] ,
    \sw_379_module_data_out[6] ,
    \sw_379_module_data_out[5] ,
    \sw_379_module_data_out[4] ,
    \sw_379_module_data_out[3] ,
    \sw_379_module_data_out[2] ,
    \sw_379_module_data_out[1] ,
    \sw_379_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_38 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_038_module_data_in[7] ,
    \sw_038_module_data_in[6] ,
    \sw_038_module_data_in[5] ,
    \sw_038_module_data_in[4] ,
    \sw_038_module_data_in[3] ,
    \sw_038_module_data_in[2] ,
    \sw_038_module_data_in[1] ,
    \sw_038_module_data_in[0] }),
    .io_out({\sw_038_module_data_out[7] ,
    \sw_038_module_data_out[6] ,
    \sw_038_module_data_out[5] ,
    \sw_038_module_data_out[4] ,
    \sw_038_module_data_out[3] ,
    \sw_038_module_data_out[2] ,
    \sw_038_module_data_out[1] ,
    \sw_038_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_380 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_380_module_data_in[7] ,
    \sw_380_module_data_in[6] ,
    \sw_380_module_data_in[5] ,
    \sw_380_module_data_in[4] ,
    \sw_380_module_data_in[3] ,
    \sw_380_module_data_in[2] ,
    \sw_380_module_data_in[1] ,
    \sw_380_module_data_in[0] }),
    .io_out({\sw_380_module_data_out[7] ,
    \sw_380_module_data_out[6] ,
    \sw_380_module_data_out[5] ,
    \sw_380_module_data_out[4] ,
    \sw_380_module_data_out[3] ,
    \sw_380_module_data_out[2] ,
    \sw_380_module_data_out[1] ,
    \sw_380_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_381 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_381_module_data_in[7] ,
    \sw_381_module_data_in[6] ,
    \sw_381_module_data_in[5] ,
    \sw_381_module_data_in[4] ,
    \sw_381_module_data_in[3] ,
    \sw_381_module_data_in[2] ,
    \sw_381_module_data_in[1] ,
    \sw_381_module_data_in[0] }),
    .io_out({\sw_381_module_data_out[7] ,
    \sw_381_module_data_out[6] ,
    \sw_381_module_data_out[5] ,
    \sw_381_module_data_out[4] ,
    \sw_381_module_data_out[3] ,
    \sw_381_module_data_out[2] ,
    \sw_381_module_data_out[1] ,
    \sw_381_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_382 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_382_module_data_in[7] ,
    \sw_382_module_data_in[6] ,
    \sw_382_module_data_in[5] ,
    \sw_382_module_data_in[4] ,
    \sw_382_module_data_in[3] ,
    \sw_382_module_data_in[2] ,
    \sw_382_module_data_in[1] ,
    \sw_382_module_data_in[0] }),
    .io_out({\sw_382_module_data_out[7] ,
    \sw_382_module_data_out[6] ,
    \sw_382_module_data_out[5] ,
    \sw_382_module_data_out[4] ,
    \sw_382_module_data_out[3] ,
    \sw_382_module_data_out[2] ,
    \sw_382_module_data_out[1] ,
    \sw_382_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_383 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_383_module_data_in[7] ,
    \sw_383_module_data_in[6] ,
    \sw_383_module_data_in[5] ,
    \sw_383_module_data_in[4] ,
    \sw_383_module_data_in[3] ,
    \sw_383_module_data_in[2] ,
    \sw_383_module_data_in[1] ,
    \sw_383_module_data_in[0] }),
    .io_out({\sw_383_module_data_out[7] ,
    \sw_383_module_data_out[6] ,
    \sw_383_module_data_out[5] ,
    \sw_383_module_data_out[4] ,
    \sw_383_module_data_out[3] ,
    \sw_383_module_data_out[2] ,
    \sw_383_module_data_out[1] ,
    \sw_383_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_384 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_384_module_data_in[7] ,
    \sw_384_module_data_in[6] ,
    \sw_384_module_data_in[5] ,
    \sw_384_module_data_in[4] ,
    \sw_384_module_data_in[3] ,
    \sw_384_module_data_in[2] ,
    \sw_384_module_data_in[1] ,
    \sw_384_module_data_in[0] }),
    .io_out({\sw_384_module_data_out[7] ,
    \sw_384_module_data_out[6] ,
    \sw_384_module_data_out[5] ,
    \sw_384_module_data_out[4] ,
    \sw_384_module_data_out[3] ,
    \sw_384_module_data_out[2] ,
    \sw_384_module_data_out[1] ,
    \sw_384_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_385 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_385_module_data_in[7] ,
    \sw_385_module_data_in[6] ,
    \sw_385_module_data_in[5] ,
    \sw_385_module_data_in[4] ,
    \sw_385_module_data_in[3] ,
    \sw_385_module_data_in[2] ,
    \sw_385_module_data_in[1] ,
    \sw_385_module_data_in[0] }),
    .io_out({\sw_385_module_data_out[7] ,
    \sw_385_module_data_out[6] ,
    \sw_385_module_data_out[5] ,
    \sw_385_module_data_out[4] ,
    \sw_385_module_data_out[3] ,
    \sw_385_module_data_out[2] ,
    \sw_385_module_data_out[1] ,
    \sw_385_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_386 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_386_module_data_in[7] ,
    \sw_386_module_data_in[6] ,
    \sw_386_module_data_in[5] ,
    \sw_386_module_data_in[4] ,
    \sw_386_module_data_in[3] ,
    \sw_386_module_data_in[2] ,
    \sw_386_module_data_in[1] ,
    \sw_386_module_data_in[0] }),
    .io_out({\sw_386_module_data_out[7] ,
    \sw_386_module_data_out[6] ,
    \sw_386_module_data_out[5] ,
    \sw_386_module_data_out[4] ,
    \sw_386_module_data_out[3] ,
    \sw_386_module_data_out[2] ,
    \sw_386_module_data_out[1] ,
    \sw_386_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_387 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_387_module_data_in[7] ,
    \sw_387_module_data_in[6] ,
    \sw_387_module_data_in[5] ,
    \sw_387_module_data_in[4] ,
    \sw_387_module_data_in[3] ,
    \sw_387_module_data_in[2] ,
    \sw_387_module_data_in[1] ,
    \sw_387_module_data_in[0] }),
    .io_out({\sw_387_module_data_out[7] ,
    \sw_387_module_data_out[6] ,
    \sw_387_module_data_out[5] ,
    \sw_387_module_data_out[4] ,
    \sw_387_module_data_out[3] ,
    \sw_387_module_data_out[2] ,
    \sw_387_module_data_out[1] ,
    \sw_387_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_388 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_388_module_data_in[7] ,
    \sw_388_module_data_in[6] ,
    \sw_388_module_data_in[5] ,
    \sw_388_module_data_in[4] ,
    \sw_388_module_data_in[3] ,
    \sw_388_module_data_in[2] ,
    \sw_388_module_data_in[1] ,
    \sw_388_module_data_in[0] }),
    .io_out({\sw_388_module_data_out[7] ,
    \sw_388_module_data_out[6] ,
    \sw_388_module_data_out[5] ,
    \sw_388_module_data_out[4] ,
    \sw_388_module_data_out[3] ,
    \sw_388_module_data_out[2] ,
    \sw_388_module_data_out[1] ,
    \sw_388_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_389 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_389_module_data_in[7] ,
    \sw_389_module_data_in[6] ,
    \sw_389_module_data_in[5] ,
    \sw_389_module_data_in[4] ,
    \sw_389_module_data_in[3] ,
    \sw_389_module_data_in[2] ,
    \sw_389_module_data_in[1] ,
    \sw_389_module_data_in[0] }),
    .io_out({\sw_389_module_data_out[7] ,
    \sw_389_module_data_out[6] ,
    \sw_389_module_data_out[5] ,
    \sw_389_module_data_out[4] ,
    \sw_389_module_data_out[3] ,
    \sw_389_module_data_out[2] ,
    \sw_389_module_data_out[1] ,
    \sw_389_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_39 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_039_module_data_in[7] ,
    \sw_039_module_data_in[6] ,
    \sw_039_module_data_in[5] ,
    \sw_039_module_data_in[4] ,
    \sw_039_module_data_in[3] ,
    \sw_039_module_data_in[2] ,
    \sw_039_module_data_in[1] ,
    \sw_039_module_data_in[0] }),
    .io_out({\sw_039_module_data_out[7] ,
    \sw_039_module_data_out[6] ,
    \sw_039_module_data_out[5] ,
    \sw_039_module_data_out[4] ,
    \sw_039_module_data_out[3] ,
    \sw_039_module_data_out[2] ,
    \sw_039_module_data_out[1] ,
    \sw_039_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_390 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_390_module_data_in[7] ,
    \sw_390_module_data_in[6] ,
    \sw_390_module_data_in[5] ,
    \sw_390_module_data_in[4] ,
    \sw_390_module_data_in[3] ,
    \sw_390_module_data_in[2] ,
    \sw_390_module_data_in[1] ,
    \sw_390_module_data_in[0] }),
    .io_out({\sw_390_module_data_out[7] ,
    \sw_390_module_data_out[6] ,
    \sw_390_module_data_out[5] ,
    \sw_390_module_data_out[4] ,
    \sw_390_module_data_out[3] ,
    \sw_390_module_data_out[2] ,
    \sw_390_module_data_out[1] ,
    \sw_390_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_391 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_391_module_data_in[7] ,
    \sw_391_module_data_in[6] ,
    \sw_391_module_data_in[5] ,
    \sw_391_module_data_in[4] ,
    \sw_391_module_data_in[3] ,
    \sw_391_module_data_in[2] ,
    \sw_391_module_data_in[1] ,
    \sw_391_module_data_in[0] }),
    .io_out({\sw_391_module_data_out[7] ,
    \sw_391_module_data_out[6] ,
    \sw_391_module_data_out[5] ,
    \sw_391_module_data_out[4] ,
    \sw_391_module_data_out[3] ,
    \sw_391_module_data_out[2] ,
    \sw_391_module_data_out[1] ,
    \sw_391_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_392 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_392_module_data_in[7] ,
    \sw_392_module_data_in[6] ,
    \sw_392_module_data_in[5] ,
    \sw_392_module_data_in[4] ,
    \sw_392_module_data_in[3] ,
    \sw_392_module_data_in[2] ,
    \sw_392_module_data_in[1] ,
    \sw_392_module_data_in[0] }),
    .io_out({\sw_392_module_data_out[7] ,
    \sw_392_module_data_out[6] ,
    \sw_392_module_data_out[5] ,
    \sw_392_module_data_out[4] ,
    \sw_392_module_data_out[3] ,
    \sw_392_module_data_out[2] ,
    \sw_392_module_data_out[1] ,
    \sw_392_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_393 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_393_module_data_in[7] ,
    \sw_393_module_data_in[6] ,
    \sw_393_module_data_in[5] ,
    \sw_393_module_data_in[4] ,
    \sw_393_module_data_in[3] ,
    \sw_393_module_data_in[2] ,
    \sw_393_module_data_in[1] ,
    \sw_393_module_data_in[0] }),
    .io_out({\sw_393_module_data_out[7] ,
    \sw_393_module_data_out[6] ,
    \sw_393_module_data_out[5] ,
    \sw_393_module_data_out[4] ,
    \sw_393_module_data_out[3] ,
    \sw_393_module_data_out[2] ,
    \sw_393_module_data_out[1] ,
    \sw_393_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_394 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_394_module_data_in[7] ,
    \sw_394_module_data_in[6] ,
    \sw_394_module_data_in[5] ,
    \sw_394_module_data_in[4] ,
    \sw_394_module_data_in[3] ,
    \sw_394_module_data_in[2] ,
    \sw_394_module_data_in[1] ,
    \sw_394_module_data_in[0] }),
    .io_out({\sw_394_module_data_out[7] ,
    \sw_394_module_data_out[6] ,
    \sw_394_module_data_out[5] ,
    \sw_394_module_data_out[4] ,
    \sw_394_module_data_out[3] ,
    \sw_394_module_data_out[2] ,
    \sw_394_module_data_out[1] ,
    \sw_394_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_395 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_395_module_data_in[7] ,
    \sw_395_module_data_in[6] ,
    \sw_395_module_data_in[5] ,
    \sw_395_module_data_in[4] ,
    \sw_395_module_data_in[3] ,
    \sw_395_module_data_in[2] ,
    \sw_395_module_data_in[1] ,
    \sw_395_module_data_in[0] }),
    .io_out({\sw_395_module_data_out[7] ,
    \sw_395_module_data_out[6] ,
    \sw_395_module_data_out[5] ,
    \sw_395_module_data_out[4] ,
    \sw_395_module_data_out[3] ,
    \sw_395_module_data_out[2] ,
    \sw_395_module_data_out[1] ,
    \sw_395_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_396 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_396_module_data_in[7] ,
    \sw_396_module_data_in[6] ,
    \sw_396_module_data_in[5] ,
    \sw_396_module_data_in[4] ,
    \sw_396_module_data_in[3] ,
    \sw_396_module_data_in[2] ,
    \sw_396_module_data_in[1] ,
    \sw_396_module_data_in[0] }),
    .io_out({\sw_396_module_data_out[7] ,
    \sw_396_module_data_out[6] ,
    \sw_396_module_data_out[5] ,
    \sw_396_module_data_out[4] ,
    \sw_396_module_data_out[3] ,
    \sw_396_module_data_out[2] ,
    \sw_396_module_data_out[1] ,
    \sw_396_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_397 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_397_module_data_in[7] ,
    \sw_397_module_data_in[6] ,
    \sw_397_module_data_in[5] ,
    \sw_397_module_data_in[4] ,
    \sw_397_module_data_in[3] ,
    \sw_397_module_data_in[2] ,
    \sw_397_module_data_in[1] ,
    \sw_397_module_data_in[0] }),
    .io_out({\sw_397_module_data_out[7] ,
    \sw_397_module_data_out[6] ,
    \sw_397_module_data_out[5] ,
    \sw_397_module_data_out[4] ,
    \sw_397_module_data_out[3] ,
    \sw_397_module_data_out[2] ,
    \sw_397_module_data_out[1] ,
    \sw_397_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_398 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_398_module_data_in[7] ,
    \sw_398_module_data_in[6] ,
    \sw_398_module_data_in[5] ,
    \sw_398_module_data_in[4] ,
    \sw_398_module_data_in[3] ,
    \sw_398_module_data_in[2] ,
    \sw_398_module_data_in[1] ,
    \sw_398_module_data_in[0] }),
    .io_out({\sw_398_module_data_out[7] ,
    \sw_398_module_data_out[6] ,
    \sw_398_module_data_out[5] ,
    \sw_398_module_data_out[4] ,
    \sw_398_module_data_out[3] ,
    \sw_398_module_data_out[2] ,
    \sw_398_module_data_out[1] ,
    \sw_398_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_399 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_399_module_data_in[7] ,
    \sw_399_module_data_in[6] ,
    \sw_399_module_data_in[5] ,
    \sw_399_module_data_in[4] ,
    \sw_399_module_data_in[3] ,
    \sw_399_module_data_in[2] ,
    \sw_399_module_data_in[1] ,
    \sw_399_module_data_in[0] }),
    .io_out({\sw_399_module_data_out[7] ,
    \sw_399_module_data_out[6] ,
    \sw_399_module_data_out[5] ,
    \sw_399_module_data_out[4] ,
    \sw_399_module_data_out[3] ,
    \sw_399_module_data_out[2] ,
    \sw_399_module_data_out[1] ,
    \sw_399_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_40 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_040_module_data_in[7] ,
    \sw_040_module_data_in[6] ,
    \sw_040_module_data_in[5] ,
    \sw_040_module_data_in[4] ,
    \sw_040_module_data_in[3] ,
    \sw_040_module_data_in[2] ,
    \sw_040_module_data_in[1] ,
    \sw_040_module_data_in[0] }),
    .io_out({\sw_040_module_data_out[7] ,
    \sw_040_module_data_out[6] ,
    \sw_040_module_data_out[5] ,
    \sw_040_module_data_out[4] ,
    \sw_040_module_data_out[3] ,
    \sw_040_module_data_out[2] ,
    \sw_040_module_data_out[1] ,
    \sw_040_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_400 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_400_module_data_in[7] ,
    \sw_400_module_data_in[6] ,
    \sw_400_module_data_in[5] ,
    \sw_400_module_data_in[4] ,
    \sw_400_module_data_in[3] ,
    \sw_400_module_data_in[2] ,
    \sw_400_module_data_in[1] ,
    \sw_400_module_data_in[0] }),
    .io_out({\sw_400_module_data_out[7] ,
    \sw_400_module_data_out[6] ,
    \sw_400_module_data_out[5] ,
    \sw_400_module_data_out[4] ,
    \sw_400_module_data_out[3] ,
    \sw_400_module_data_out[2] ,
    \sw_400_module_data_out[1] ,
    \sw_400_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_401 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_401_module_data_in[7] ,
    \sw_401_module_data_in[6] ,
    \sw_401_module_data_in[5] ,
    \sw_401_module_data_in[4] ,
    \sw_401_module_data_in[3] ,
    \sw_401_module_data_in[2] ,
    \sw_401_module_data_in[1] ,
    \sw_401_module_data_in[0] }),
    .io_out({\sw_401_module_data_out[7] ,
    \sw_401_module_data_out[6] ,
    \sw_401_module_data_out[5] ,
    \sw_401_module_data_out[4] ,
    \sw_401_module_data_out[3] ,
    \sw_401_module_data_out[2] ,
    \sw_401_module_data_out[1] ,
    \sw_401_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_402 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_402_module_data_in[7] ,
    \sw_402_module_data_in[6] ,
    \sw_402_module_data_in[5] ,
    \sw_402_module_data_in[4] ,
    \sw_402_module_data_in[3] ,
    \sw_402_module_data_in[2] ,
    \sw_402_module_data_in[1] ,
    \sw_402_module_data_in[0] }),
    .io_out({\sw_402_module_data_out[7] ,
    \sw_402_module_data_out[6] ,
    \sw_402_module_data_out[5] ,
    \sw_402_module_data_out[4] ,
    \sw_402_module_data_out[3] ,
    \sw_402_module_data_out[2] ,
    \sw_402_module_data_out[1] ,
    \sw_402_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_403 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_403_module_data_in[7] ,
    \sw_403_module_data_in[6] ,
    \sw_403_module_data_in[5] ,
    \sw_403_module_data_in[4] ,
    \sw_403_module_data_in[3] ,
    \sw_403_module_data_in[2] ,
    \sw_403_module_data_in[1] ,
    \sw_403_module_data_in[0] }),
    .io_out({\sw_403_module_data_out[7] ,
    \sw_403_module_data_out[6] ,
    \sw_403_module_data_out[5] ,
    \sw_403_module_data_out[4] ,
    \sw_403_module_data_out[3] ,
    \sw_403_module_data_out[2] ,
    \sw_403_module_data_out[1] ,
    \sw_403_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_404 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_404_module_data_in[7] ,
    \sw_404_module_data_in[6] ,
    \sw_404_module_data_in[5] ,
    \sw_404_module_data_in[4] ,
    \sw_404_module_data_in[3] ,
    \sw_404_module_data_in[2] ,
    \sw_404_module_data_in[1] ,
    \sw_404_module_data_in[0] }),
    .io_out({\sw_404_module_data_out[7] ,
    \sw_404_module_data_out[6] ,
    \sw_404_module_data_out[5] ,
    \sw_404_module_data_out[4] ,
    \sw_404_module_data_out[3] ,
    \sw_404_module_data_out[2] ,
    \sw_404_module_data_out[1] ,
    \sw_404_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_405 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_405_module_data_in[7] ,
    \sw_405_module_data_in[6] ,
    \sw_405_module_data_in[5] ,
    \sw_405_module_data_in[4] ,
    \sw_405_module_data_in[3] ,
    \sw_405_module_data_in[2] ,
    \sw_405_module_data_in[1] ,
    \sw_405_module_data_in[0] }),
    .io_out({\sw_405_module_data_out[7] ,
    \sw_405_module_data_out[6] ,
    \sw_405_module_data_out[5] ,
    \sw_405_module_data_out[4] ,
    \sw_405_module_data_out[3] ,
    \sw_405_module_data_out[2] ,
    \sw_405_module_data_out[1] ,
    \sw_405_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_406 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_406_module_data_in[7] ,
    \sw_406_module_data_in[6] ,
    \sw_406_module_data_in[5] ,
    \sw_406_module_data_in[4] ,
    \sw_406_module_data_in[3] ,
    \sw_406_module_data_in[2] ,
    \sw_406_module_data_in[1] ,
    \sw_406_module_data_in[0] }),
    .io_out({\sw_406_module_data_out[7] ,
    \sw_406_module_data_out[6] ,
    \sw_406_module_data_out[5] ,
    \sw_406_module_data_out[4] ,
    \sw_406_module_data_out[3] ,
    \sw_406_module_data_out[2] ,
    \sw_406_module_data_out[1] ,
    \sw_406_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_407 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_407_module_data_in[7] ,
    \sw_407_module_data_in[6] ,
    \sw_407_module_data_in[5] ,
    \sw_407_module_data_in[4] ,
    \sw_407_module_data_in[3] ,
    \sw_407_module_data_in[2] ,
    \sw_407_module_data_in[1] ,
    \sw_407_module_data_in[0] }),
    .io_out({\sw_407_module_data_out[7] ,
    \sw_407_module_data_out[6] ,
    \sw_407_module_data_out[5] ,
    \sw_407_module_data_out[4] ,
    \sw_407_module_data_out[3] ,
    \sw_407_module_data_out[2] ,
    \sw_407_module_data_out[1] ,
    \sw_407_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_408 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_408_module_data_in[7] ,
    \sw_408_module_data_in[6] ,
    \sw_408_module_data_in[5] ,
    \sw_408_module_data_in[4] ,
    \sw_408_module_data_in[3] ,
    \sw_408_module_data_in[2] ,
    \sw_408_module_data_in[1] ,
    \sw_408_module_data_in[0] }),
    .io_out({\sw_408_module_data_out[7] ,
    \sw_408_module_data_out[6] ,
    \sw_408_module_data_out[5] ,
    \sw_408_module_data_out[4] ,
    \sw_408_module_data_out[3] ,
    \sw_408_module_data_out[2] ,
    \sw_408_module_data_out[1] ,
    \sw_408_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_409 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_409_module_data_in[7] ,
    \sw_409_module_data_in[6] ,
    \sw_409_module_data_in[5] ,
    \sw_409_module_data_in[4] ,
    \sw_409_module_data_in[3] ,
    \sw_409_module_data_in[2] ,
    \sw_409_module_data_in[1] ,
    \sw_409_module_data_in[0] }),
    .io_out({\sw_409_module_data_out[7] ,
    \sw_409_module_data_out[6] ,
    \sw_409_module_data_out[5] ,
    \sw_409_module_data_out[4] ,
    \sw_409_module_data_out[3] ,
    \sw_409_module_data_out[2] ,
    \sw_409_module_data_out[1] ,
    \sw_409_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_41 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_041_module_data_in[7] ,
    \sw_041_module_data_in[6] ,
    \sw_041_module_data_in[5] ,
    \sw_041_module_data_in[4] ,
    \sw_041_module_data_in[3] ,
    \sw_041_module_data_in[2] ,
    \sw_041_module_data_in[1] ,
    \sw_041_module_data_in[0] }),
    .io_out({\sw_041_module_data_out[7] ,
    \sw_041_module_data_out[6] ,
    \sw_041_module_data_out[5] ,
    \sw_041_module_data_out[4] ,
    \sw_041_module_data_out[3] ,
    \sw_041_module_data_out[2] ,
    \sw_041_module_data_out[1] ,
    \sw_041_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_410 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_410_module_data_in[7] ,
    \sw_410_module_data_in[6] ,
    \sw_410_module_data_in[5] ,
    \sw_410_module_data_in[4] ,
    \sw_410_module_data_in[3] ,
    \sw_410_module_data_in[2] ,
    \sw_410_module_data_in[1] ,
    \sw_410_module_data_in[0] }),
    .io_out({\sw_410_module_data_out[7] ,
    \sw_410_module_data_out[6] ,
    \sw_410_module_data_out[5] ,
    \sw_410_module_data_out[4] ,
    \sw_410_module_data_out[3] ,
    \sw_410_module_data_out[2] ,
    \sw_410_module_data_out[1] ,
    \sw_410_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_411 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_411_module_data_in[7] ,
    \sw_411_module_data_in[6] ,
    \sw_411_module_data_in[5] ,
    \sw_411_module_data_in[4] ,
    \sw_411_module_data_in[3] ,
    \sw_411_module_data_in[2] ,
    \sw_411_module_data_in[1] ,
    \sw_411_module_data_in[0] }),
    .io_out({\sw_411_module_data_out[7] ,
    \sw_411_module_data_out[6] ,
    \sw_411_module_data_out[5] ,
    \sw_411_module_data_out[4] ,
    \sw_411_module_data_out[3] ,
    \sw_411_module_data_out[2] ,
    \sw_411_module_data_out[1] ,
    \sw_411_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_412 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_412_module_data_in[7] ,
    \sw_412_module_data_in[6] ,
    \sw_412_module_data_in[5] ,
    \sw_412_module_data_in[4] ,
    \sw_412_module_data_in[3] ,
    \sw_412_module_data_in[2] ,
    \sw_412_module_data_in[1] ,
    \sw_412_module_data_in[0] }),
    .io_out({\sw_412_module_data_out[7] ,
    \sw_412_module_data_out[6] ,
    \sw_412_module_data_out[5] ,
    \sw_412_module_data_out[4] ,
    \sw_412_module_data_out[3] ,
    \sw_412_module_data_out[2] ,
    \sw_412_module_data_out[1] ,
    \sw_412_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_413 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_413_module_data_in[7] ,
    \sw_413_module_data_in[6] ,
    \sw_413_module_data_in[5] ,
    \sw_413_module_data_in[4] ,
    \sw_413_module_data_in[3] ,
    \sw_413_module_data_in[2] ,
    \sw_413_module_data_in[1] ,
    \sw_413_module_data_in[0] }),
    .io_out({\sw_413_module_data_out[7] ,
    \sw_413_module_data_out[6] ,
    \sw_413_module_data_out[5] ,
    \sw_413_module_data_out[4] ,
    \sw_413_module_data_out[3] ,
    \sw_413_module_data_out[2] ,
    \sw_413_module_data_out[1] ,
    \sw_413_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_414 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_414_module_data_in[7] ,
    \sw_414_module_data_in[6] ,
    \sw_414_module_data_in[5] ,
    \sw_414_module_data_in[4] ,
    \sw_414_module_data_in[3] ,
    \sw_414_module_data_in[2] ,
    \sw_414_module_data_in[1] ,
    \sw_414_module_data_in[0] }),
    .io_out({\sw_414_module_data_out[7] ,
    \sw_414_module_data_out[6] ,
    \sw_414_module_data_out[5] ,
    \sw_414_module_data_out[4] ,
    \sw_414_module_data_out[3] ,
    \sw_414_module_data_out[2] ,
    \sw_414_module_data_out[1] ,
    \sw_414_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_415 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_415_module_data_in[7] ,
    \sw_415_module_data_in[6] ,
    \sw_415_module_data_in[5] ,
    \sw_415_module_data_in[4] ,
    \sw_415_module_data_in[3] ,
    \sw_415_module_data_in[2] ,
    \sw_415_module_data_in[1] ,
    \sw_415_module_data_in[0] }),
    .io_out({\sw_415_module_data_out[7] ,
    \sw_415_module_data_out[6] ,
    \sw_415_module_data_out[5] ,
    \sw_415_module_data_out[4] ,
    \sw_415_module_data_out[3] ,
    \sw_415_module_data_out[2] ,
    \sw_415_module_data_out[1] ,
    \sw_415_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_416 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_416_module_data_in[7] ,
    \sw_416_module_data_in[6] ,
    \sw_416_module_data_in[5] ,
    \sw_416_module_data_in[4] ,
    \sw_416_module_data_in[3] ,
    \sw_416_module_data_in[2] ,
    \sw_416_module_data_in[1] ,
    \sw_416_module_data_in[0] }),
    .io_out({\sw_416_module_data_out[7] ,
    \sw_416_module_data_out[6] ,
    \sw_416_module_data_out[5] ,
    \sw_416_module_data_out[4] ,
    \sw_416_module_data_out[3] ,
    \sw_416_module_data_out[2] ,
    \sw_416_module_data_out[1] ,
    \sw_416_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_417 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_417_module_data_in[7] ,
    \sw_417_module_data_in[6] ,
    \sw_417_module_data_in[5] ,
    \sw_417_module_data_in[4] ,
    \sw_417_module_data_in[3] ,
    \sw_417_module_data_in[2] ,
    \sw_417_module_data_in[1] ,
    \sw_417_module_data_in[0] }),
    .io_out({\sw_417_module_data_out[7] ,
    \sw_417_module_data_out[6] ,
    \sw_417_module_data_out[5] ,
    \sw_417_module_data_out[4] ,
    \sw_417_module_data_out[3] ,
    \sw_417_module_data_out[2] ,
    \sw_417_module_data_out[1] ,
    \sw_417_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_418 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_418_module_data_in[7] ,
    \sw_418_module_data_in[6] ,
    \sw_418_module_data_in[5] ,
    \sw_418_module_data_in[4] ,
    \sw_418_module_data_in[3] ,
    \sw_418_module_data_in[2] ,
    \sw_418_module_data_in[1] ,
    \sw_418_module_data_in[0] }),
    .io_out({\sw_418_module_data_out[7] ,
    \sw_418_module_data_out[6] ,
    \sw_418_module_data_out[5] ,
    \sw_418_module_data_out[4] ,
    \sw_418_module_data_out[3] ,
    \sw_418_module_data_out[2] ,
    \sw_418_module_data_out[1] ,
    \sw_418_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_419 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_419_module_data_in[7] ,
    \sw_419_module_data_in[6] ,
    \sw_419_module_data_in[5] ,
    \sw_419_module_data_in[4] ,
    \sw_419_module_data_in[3] ,
    \sw_419_module_data_in[2] ,
    \sw_419_module_data_in[1] ,
    \sw_419_module_data_in[0] }),
    .io_out({\sw_419_module_data_out[7] ,
    \sw_419_module_data_out[6] ,
    \sw_419_module_data_out[5] ,
    \sw_419_module_data_out[4] ,
    \sw_419_module_data_out[3] ,
    \sw_419_module_data_out[2] ,
    \sw_419_module_data_out[1] ,
    \sw_419_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_42 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_042_module_data_in[7] ,
    \sw_042_module_data_in[6] ,
    \sw_042_module_data_in[5] ,
    \sw_042_module_data_in[4] ,
    \sw_042_module_data_in[3] ,
    \sw_042_module_data_in[2] ,
    \sw_042_module_data_in[1] ,
    \sw_042_module_data_in[0] }),
    .io_out({\sw_042_module_data_out[7] ,
    \sw_042_module_data_out[6] ,
    \sw_042_module_data_out[5] ,
    \sw_042_module_data_out[4] ,
    \sw_042_module_data_out[3] ,
    \sw_042_module_data_out[2] ,
    \sw_042_module_data_out[1] ,
    \sw_042_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_420 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_420_module_data_in[7] ,
    \sw_420_module_data_in[6] ,
    \sw_420_module_data_in[5] ,
    \sw_420_module_data_in[4] ,
    \sw_420_module_data_in[3] ,
    \sw_420_module_data_in[2] ,
    \sw_420_module_data_in[1] ,
    \sw_420_module_data_in[0] }),
    .io_out({\sw_420_module_data_out[7] ,
    \sw_420_module_data_out[6] ,
    \sw_420_module_data_out[5] ,
    \sw_420_module_data_out[4] ,
    \sw_420_module_data_out[3] ,
    \sw_420_module_data_out[2] ,
    \sw_420_module_data_out[1] ,
    \sw_420_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_421 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_421_module_data_in[7] ,
    \sw_421_module_data_in[6] ,
    \sw_421_module_data_in[5] ,
    \sw_421_module_data_in[4] ,
    \sw_421_module_data_in[3] ,
    \sw_421_module_data_in[2] ,
    \sw_421_module_data_in[1] ,
    \sw_421_module_data_in[0] }),
    .io_out({\sw_421_module_data_out[7] ,
    \sw_421_module_data_out[6] ,
    \sw_421_module_data_out[5] ,
    \sw_421_module_data_out[4] ,
    \sw_421_module_data_out[3] ,
    \sw_421_module_data_out[2] ,
    \sw_421_module_data_out[1] ,
    \sw_421_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_422 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_422_module_data_in[7] ,
    \sw_422_module_data_in[6] ,
    \sw_422_module_data_in[5] ,
    \sw_422_module_data_in[4] ,
    \sw_422_module_data_in[3] ,
    \sw_422_module_data_in[2] ,
    \sw_422_module_data_in[1] ,
    \sw_422_module_data_in[0] }),
    .io_out({\sw_422_module_data_out[7] ,
    \sw_422_module_data_out[6] ,
    \sw_422_module_data_out[5] ,
    \sw_422_module_data_out[4] ,
    \sw_422_module_data_out[3] ,
    \sw_422_module_data_out[2] ,
    \sw_422_module_data_out[1] ,
    \sw_422_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_423 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_423_module_data_in[7] ,
    \sw_423_module_data_in[6] ,
    \sw_423_module_data_in[5] ,
    \sw_423_module_data_in[4] ,
    \sw_423_module_data_in[3] ,
    \sw_423_module_data_in[2] ,
    \sw_423_module_data_in[1] ,
    \sw_423_module_data_in[0] }),
    .io_out({\sw_423_module_data_out[7] ,
    \sw_423_module_data_out[6] ,
    \sw_423_module_data_out[5] ,
    \sw_423_module_data_out[4] ,
    \sw_423_module_data_out[3] ,
    \sw_423_module_data_out[2] ,
    \sw_423_module_data_out[1] ,
    \sw_423_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_424 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_424_module_data_in[7] ,
    \sw_424_module_data_in[6] ,
    \sw_424_module_data_in[5] ,
    \sw_424_module_data_in[4] ,
    \sw_424_module_data_in[3] ,
    \sw_424_module_data_in[2] ,
    \sw_424_module_data_in[1] ,
    \sw_424_module_data_in[0] }),
    .io_out({\sw_424_module_data_out[7] ,
    \sw_424_module_data_out[6] ,
    \sw_424_module_data_out[5] ,
    \sw_424_module_data_out[4] ,
    \sw_424_module_data_out[3] ,
    \sw_424_module_data_out[2] ,
    \sw_424_module_data_out[1] ,
    \sw_424_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_425 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_425_module_data_in[7] ,
    \sw_425_module_data_in[6] ,
    \sw_425_module_data_in[5] ,
    \sw_425_module_data_in[4] ,
    \sw_425_module_data_in[3] ,
    \sw_425_module_data_in[2] ,
    \sw_425_module_data_in[1] ,
    \sw_425_module_data_in[0] }),
    .io_out({\sw_425_module_data_out[7] ,
    \sw_425_module_data_out[6] ,
    \sw_425_module_data_out[5] ,
    \sw_425_module_data_out[4] ,
    \sw_425_module_data_out[3] ,
    \sw_425_module_data_out[2] ,
    \sw_425_module_data_out[1] ,
    \sw_425_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_426 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_426_module_data_in[7] ,
    \sw_426_module_data_in[6] ,
    \sw_426_module_data_in[5] ,
    \sw_426_module_data_in[4] ,
    \sw_426_module_data_in[3] ,
    \sw_426_module_data_in[2] ,
    \sw_426_module_data_in[1] ,
    \sw_426_module_data_in[0] }),
    .io_out({\sw_426_module_data_out[7] ,
    \sw_426_module_data_out[6] ,
    \sw_426_module_data_out[5] ,
    \sw_426_module_data_out[4] ,
    \sw_426_module_data_out[3] ,
    \sw_426_module_data_out[2] ,
    \sw_426_module_data_out[1] ,
    \sw_426_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_427 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_427_module_data_in[7] ,
    \sw_427_module_data_in[6] ,
    \sw_427_module_data_in[5] ,
    \sw_427_module_data_in[4] ,
    \sw_427_module_data_in[3] ,
    \sw_427_module_data_in[2] ,
    \sw_427_module_data_in[1] ,
    \sw_427_module_data_in[0] }),
    .io_out({\sw_427_module_data_out[7] ,
    \sw_427_module_data_out[6] ,
    \sw_427_module_data_out[5] ,
    \sw_427_module_data_out[4] ,
    \sw_427_module_data_out[3] ,
    \sw_427_module_data_out[2] ,
    \sw_427_module_data_out[1] ,
    \sw_427_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_428 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_428_module_data_in[7] ,
    \sw_428_module_data_in[6] ,
    \sw_428_module_data_in[5] ,
    \sw_428_module_data_in[4] ,
    \sw_428_module_data_in[3] ,
    \sw_428_module_data_in[2] ,
    \sw_428_module_data_in[1] ,
    \sw_428_module_data_in[0] }),
    .io_out({\sw_428_module_data_out[7] ,
    \sw_428_module_data_out[6] ,
    \sw_428_module_data_out[5] ,
    \sw_428_module_data_out[4] ,
    \sw_428_module_data_out[3] ,
    \sw_428_module_data_out[2] ,
    \sw_428_module_data_out[1] ,
    \sw_428_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_429 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_429_module_data_in[7] ,
    \sw_429_module_data_in[6] ,
    \sw_429_module_data_in[5] ,
    \sw_429_module_data_in[4] ,
    \sw_429_module_data_in[3] ,
    \sw_429_module_data_in[2] ,
    \sw_429_module_data_in[1] ,
    \sw_429_module_data_in[0] }),
    .io_out({\sw_429_module_data_out[7] ,
    \sw_429_module_data_out[6] ,
    \sw_429_module_data_out[5] ,
    \sw_429_module_data_out[4] ,
    \sw_429_module_data_out[3] ,
    \sw_429_module_data_out[2] ,
    \sw_429_module_data_out[1] ,
    \sw_429_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_43 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_043_module_data_in[7] ,
    \sw_043_module_data_in[6] ,
    \sw_043_module_data_in[5] ,
    \sw_043_module_data_in[4] ,
    \sw_043_module_data_in[3] ,
    \sw_043_module_data_in[2] ,
    \sw_043_module_data_in[1] ,
    \sw_043_module_data_in[0] }),
    .io_out({\sw_043_module_data_out[7] ,
    \sw_043_module_data_out[6] ,
    \sw_043_module_data_out[5] ,
    \sw_043_module_data_out[4] ,
    \sw_043_module_data_out[3] ,
    \sw_043_module_data_out[2] ,
    \sw_043_module_data_out[1] ,
    \sw_043_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_430 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_430_module_data_in[7] ,
    \sw_430_module_data_in[6] ,
    \sw_430_module_data_in[5] ,
    \sw_430_module_data_in[4] ,
    \sw_430_module_data_in[3] ,
    \sw_430_module_data_in[2] ,
    \sw_430_module_data_in[1] ,
    \sw_430_module_data_in[0] }),
    .io_out({\sw_430_module_data_out[7] ,
    \sw_430_module_data_out[6] ,
    \sw_430_module_data_out[5] ,
    \sw_430_module_data_out[4] ,
    \sw_430_module_data_out[3] ,
    \sw_430_module_data_out[2] ,
    \sw_430_module_data_out[1] ,
    \sw_430_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_431 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_431_module_data_in[7] ,
    \sw_431_module_data_in[6] ,
    \sw_431_module_data_in[5] ,
    \sw_431_module_data_in[4] ,
    \sw_431_module_data_in[3] ,
    \sw_431_module_data_in[2] ,
    \sw_431_module_data_in[1] ,
    \sw_431_module_data_in[0] }),
    .io_out({\sw_431_module_data_out[7] ,
    \sw_431_module_data_out[6] ,
    \sw_431_module_data_out[5] ,
    \sw_431_module_data_out[4] ,
    \sw_431_module_data_out[3] ,
    \sw_431_module_data_out[2] ,
    \sw_431_module_data_out[1] ,
    \sw_431_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_432 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_432_module_data_in[7] ,
    \sw_432_module_data_in[6] ,
    \sw_432_module_data_in[5] ,
    \sw_432_module_data_in[4] ,
    \sw_432_module_data_in[3] ,
    \sw_432_module_data_in[2] ,
    \sw_432_module_data_in[1] ,
    \sw_432_module_data_in[0] }),
    .io_out({\sw_432_module_data_out[7] ,
    \sw_432_module_data_out[6] ,
    \sw_432_module_data_out[5] ,
    \sw_432_module_data_out[4] ,
    \sw_432_module_data_out[3] ,
    \sw_432_module_data_out[2] ,
    \sw_432_module_data_out[1] ,
    \sw_432_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_433 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_433_module_data_in[7] ,
    \sw_433_module_data_in[6] ,
    \sw_433_module_data_in[5] ,
    \sw_433_module_data_in[4] ,
    \sw_433_module_data_in[3] ,
    \sw_433_module_data_in[2] ,
    \sw_433_module_data_in[1] ,
    \sw_433_module_data_in[0] }),
    .io_out({\sw_433_module_data_out[7] ,
    \sw_433_module_data_out[6] ,
    \sw_433_module_data_out[5] ,
    \sw_433_module_data_out[4] ,
    \sw_433_module_data_out[3] ,
    \sw_433_module_data_out[2] ,
    \sw_433_module_data_out[1] ,
    \sw_433_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_434 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_434_module_data_in[7] ,
    \sw_434_module_data_in[6] ,
    \sw_434_module_data_in[5] ,
    \sw_434_module_data_in[4] ,
    \sw_434_module_data_in[3] ,
    \sw_434_module_data_in[2] ,
    \sw_434_module_data_in[1] ,
    \sw_434_module_data_in[0] }),
    .io_out({\sw_434_module_data_out[7] ,
    \sw_434_module_data_out[6] ,
    \sw_434_module_data_out[5] ,
    \sw_434_module_data_out[4] ,
    \sw_434_module_data_out[3] ,
    \sw_434_module_data_out[2] ,
    \sw_434_module_data_out[1] ,
    \sw_434_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_435 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_435_module_data_in[7] ,
    \sw_435_module_data_in[6] ,
    \sw_435_module_data_in[5] ,
    \sw_435_module_data_in[4] ,
    \sw_435_module_data_in[3] ,
    \sw_435_module_data_in[2] ,
    \sw_435_module_data_in[1] ,
    \sw_435_module_data_in[0] }),
    .io_out({\sw_435_module_data_out[7] ,
    \sw_435_module_data_out[6] ,
    \sw_435_module_data_out[5] ,
    \sw_435_module_data_out[4] ,
    \sw_435_module_data_out[3] ,
    \sw_435_module_data_out[2] ,
    \sw_435_module_data_out[1] ,
    \sw_435_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_436 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_436_module_data_in[7] ,
    \sw_436_module_data_in[6] ,
    \sw_436_module_data_in[5] ,
    \sw_436_module_data_in[4] ,
    \sw_436_module_data_in[3] ,
    \sw_436_module_data_in[2] ,
    \sw_436_module_data_in[1] ,
    \sw_436_module_data_in[0] }),
    .io_out({\sw_436_module_data_out[7] ,
    \sw_436_module_data_out[6] ,
    \sw_436_module_data_out[5] ,
    \sw_436_module_data_out[4] ,
    \sw_436_module_data_out[3] ,
    \sw_436_module_data_out[2] ,
    \sw_436_module_data_out[1] ,
    \sw_436_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_437 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_437_module_data_in[7] ,
    \sw_437_module_data_in[6] ,
    \sw_437_module_data_in[5] ,
    \sw_437_module_data_in[4] ,
    \sw_437_module_data_in[3] ,
    \sw_437_module_data_in[2] ,
    \sw_437_module_data_in[1] ,
    \sw_437_module_data_in[0] }),
    .io_out({\sw_437_module_data_out[7] ,
    \sw_437_module_data_out[6] ,
    \sw_437_module_data_out[5] ,
    \sw_437_module_data_out[4] ,
    \sw_437_module_data_out[3] ,
    \sw_437_module_data_out[2] ,
    \sw_437_module_data_out[1] ,
    \sw_437_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_438 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_438_module_data_in[7] ,
    \sw_438_module_data_in[6] ,
    \sw_438_module_data_in[5] ,
    \sw_438_module_data_in[4] ,
    \sw_438_module_data_in[3] ,
    \sw_438_module_data_in[2] ,
    \sw_438_module_data_in[1] ,
    \sw_438_module_data_in[0] }),
    .io_out({\sw_438_module_data_out[7] ,
    \sw_438_module_data_out[6] ,
    \sw_438_module_data_out[5] ,
    \sw_438_module_data_out[4] ,
    \sw_438_module_data_out[3] ,
    \sw_438_module_data_out[2] ,
    \sw_438_module_data_out[1] ,
    \sw_438_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_439 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_439_module_data_in[7] ,
    \sw_439_module_data_in[6] ,
    \sw_439_module_data_in[5] ,
    \sw_439_module_data_in[4] ,
    \sw_439_module_data_in[3] ,
    \sw_439_module_data_in[2] ,
    \sw_439_module_data_in[1] ,
    \sw_439_module_data_in[0] }),
    .io_out({\sw_439_module_data_out[7] ,
    \sw_439_module_data_out[6] ,
    \sw_439_module_data_out[5] ,
    \sw_439_module_data_out[4] ,
    \sw_439_module_data_out[3] ,
    \sw_439_module_data_out[2] ,
    \sw_439_module_data_out[1] ,
    \sw_439_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_44 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_044_module_data_in[7] ,
    \sw_044_module_data_in[6] ,
    \sw_044_module_data_in[5] ,
    \sw_044_module_data_in[4] ,
    \sw_044_module_data_in[3] ,
    \sw_044_module_data_in[2] ,
    \sw_044_module_data_in[1] ,
    \sw_044_module_data_in[0] }),
    .io_out({\sw_044_module_data_out[7] ,
    \sw_044_module_data_out[6] ,
    \sw_044_module_data_out[5] ,
    \sw_044_module_data_out[4] ,
    \sw_044_module_data_out[3] ,
    \sw_044_module_data_out[2] ,
    \sw_044_module_data_out[1] ,
    \sw_044_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_440 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_440_module_data_in[7] ,
    \sw_440_module_data_in[6] ,
    \sw_440_module_data_in[5] ,
    \sw_440_module_data_in[4] ,
    \sw_440_module_data_in[3] ,
    \sw_440_module_data_in[2] ,
    \sw_440_module_data_in[1] ,
    \sw_440_module_data_in[0] }),
    .io_out({\sw_440_module_data_out[7] ,
    \sw_440_module_data_out[6] ,
    \sw_440_module_data_out[5] ,
    \sw_440_module_data_out[4] ,
    \sw_440_module_data_out[3] ,
    \sw_440_module_data_out[2] ,
    \sw_440_module_data_out[1] ,
    \sw_440_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_441 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_441_module_data_in[7] ,
    \sw_441_module_data_in[6] ,
    \sw_441_module_data_in[5] ,
    \sw_441_module_data_in[4] ,
    \sw_441_module_data_in[3] ,
    \sw_441_module_data_in[2] ,
    \sw_441_module_data_in[1] ,
    \sw_441_module_data_in[0] }),
    .io_out({\sw_441_module_data_out[7] ,
    \sw_441_module_data_out[6] ,
    \sw_441_module_data_out[5] ,
    \sw_441_module_data_out[4] ,
    \sw_441_module_data_out[3] ,
    \sw_441_module_data_out[2] ,
    \sw_441_module_data_out[1] ,
    \sw_441_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_442 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_442_module_data_in[7] ,
    \sw_442_module_data_in[6] ,
    \sw_442_module_data_in[5] ,
    \sw_442_module_data_in[4] ,
    \sw_442_module_data_in[3] ,
    \sw_442_module_data_in[2] ,
    \sw_442_module_data_in[1] ,
    \sw_442_module_data_in[0] }),
    .io_out({\sw_442_module_data_out[7] ,
    \sw_442_module_data_out[6] ,
    \sw_442_module_data_out[5] ,
    \sw_442_module_data_out[4] ,
    \sw_442_module_data_out[3] ,
    \sw_442_module_data_out[2] ,
    \sw_442_module_data_out[1] ,
    \sw_442_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_443 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_443_module_data_in[7] ,
    \sw_443_module_data_in[6] ,
    \sw_443_module_data_in[5] ,
    \sw_443_module_data_in[4] ,
    \sw_443_module_data_in[3] ,
    \sw_443_module_data_in[2] ,
    \sw_443_module_data_in[1] ,
    \sw_443_module_data_in[0] }),
    .io_out({\sw_443_module_data_out[7] ,
    \sw_443_module_data_out[6] ,
    \sw_443_module_data_out[5] ,
    \sw_443_module_data_out[4] ,
    \sw_443_module_data_out[3] ,
    \sw_443_module_data_out[2] ,
    \sw_443_module_data_out[1] ,
    \sw_443_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_444 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_444_module_data_in[7] ,
    \sw_444_module_data_in[6] ,
    \sw_444_module_data_in[5] ,
    \sw_444_module_data_in[4] ,
    \sw_444_module_data_in[3] ,
    \sw_444_module_data_in[2] ,
    \sw_444_module_data_in[1] ,
    \sw_444_module_data_in[0] }),
    .io_out({\sw_444_module_data_out[7] ,
    \sw_444_module_data_out[6] ,
    \sw_444_module_data_out[5] ,
    \sw_444_module_data_out[4] ,
    \sw_444_module_data_out[3] ,
    \sw_444_module_data_out[2] ,
    \sw_444_module_data_out[1] ,
    \sw_444_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_445 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_445_module_data_in[7] ,
    \sw_445_module_data_in[6] ,
    \sw_445_module_data_in[5] ,
    \sw_445_module_data_in[4] ,
    \sw_445_module_data_in[3] ,
    \sw_445_module_data_in[2] ,
    \sw_445_module_data_in[1] ,
    \sw_445_module_data_in[0] }),
    .io_out({\sw_445_module_data_out[7] ,
    \sw_445_module_data_out[6] ,
    \sw_445_module_data_out[5] ,
    \sw_445_module_data_out[4] ,
    \sw_445_module_data_out[3] ,
    \sw_445_module_data_out[2] ,
    \sw_445_module_data_out[1] ,
    \sw_445_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_446 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_446_module_data_in[7] ,
    \sw_446_module_data_in[6] ,
    \sw_446_module_data_in[5] ,
    \sw_446_module_data_in[4] ,
    \sw_446_module_data_in[3] ,
    \sw_446_module_data_in[2] ,
    \sw_446_module_data_in[1] ,
    \sw_446_module_data_in[0] }),
    .io_out({\sw_446_module_data_out[7] ,
    \sw_446_module_data_out[6] ,
    \sw_446_module_data_out[5] ,
    \sw_446_module_data_out[4] ,
    \sw_446_module_data_out[3] ,
    \sw_446_module_data_out[2] ,
    \sw_446_module_data_out[1] ,
    \sw_446_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_447 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_447_module_data_in[7] ,
    \sw_447_module_data_in[6] ,
    \sw_447_module_data_in[5] ,
    \sw_447_module_data_in[4] ,
    \sw_447_module_data_in[3] ,
    \sw_447_module_data_in[2] ,
    \sw_447_module_data_in[1] ,
    \sw_447_module_data_in[0] }),
    .io_out({\sw_447_module_data_out[7] ,
    \sw_447_module_data_out[6] ,
    \sw_447_module_data_out[5] ,
    \sw_447_module_data_out[4] ,
    \sw_447_module_data_out[3] ,
    \sw_447_module_data_out[2] ,
    \sw_447_module_data_out[1] ,
    \sw_447_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_448 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_448_module_data_in[7] ,
    \sw_448_module_data_in[6] ,
    \sw_448_module_data_in[5] ,
    \sw_448_module_data_in[4] ,
    \sw_448_module_data_in[3] ,
    \sw_448_module_data_in[2] ,
    \sw_448_module_data_in[1] ,
    \sw_448_module_data_in[0] }),
    .io_out({\sw_448_module_data_out[7] ,
    \sw_448_module_data_out[6] ,
    \sw_448_module_data_out[5] ,
    \sw_448_module_data_out[4] ,
    \sw_448_module_data_out[3] ,
    \sw_448_module_data_out[2] ,
    \sw_448_module_data_out[1] ,
    \sw_448_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_449 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_449_module_data_in[7] ,
    \sw_449_module_data_in[6] ,
    \sw_449_module_data_in[5] ,
    \sw_449_module_data_in[4] ,
    \sw_449_module_data_in[3] ,
    \sw_449_module_data_in[2] ,
    \sw_449_module_data_in[1] ,
    \sw_449_module_data_in[0] }),
    .io_out({\sw_449_module_data_out[7] ,
    \sw_449_module_data_out[6] ,
    \sw_449_module_data_out[5] ,
    \sw_449_module_data_out[4] ,
    \sw_449_module_data_out[3] ,
    \sw_449_module_data_out[2] ,
    \sw_449_module_data_out[1] ,
    \sw_449_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_45 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_045_module_data_in[7] ,
    \sw_045_module_data_in[6] ,
    \sw_045_module_data_in[5] ,
    \sw_045_module_data_in[4] ,
    \sw_045_module_data_in[3] ,
    \sw_045_module_data_in[2] ,
    \sw_045_module_data_in[1] ,
    \sw_045_module_data_in[0] }),
    .io_out({\sw_045_module_data_out[7] ,
    \sw_045_module_data_out[6] ,
    \sw_045_module_data_out[5] ,
    \sw_045_module_data_out[4] ,
    \sw_045_module_data_out[3] ,
    \sw_045_module_data_out[2] ,
    \sw_045_module_data_out[1] ,
    \sw_045_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_450 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_450_module_data_in[7] ,
    \sw_450_module_data_in[6] ,
    \sw_450_module_data_in[5] ,
    \sw_450_module_data_in[4] ,
    \sw_450_module_data_in[3] ,
    \sw_450_module_data_in[2] ,
    \sw_450_module_data_in[1] ,
    \sw_450_module_data_in[0] }),
    .io_out({\sw_450_module_data_out[7] ,
    \sw_450_module_data_out[6] ,
    \sw_450_module_data_out[5] ,
    \sw_450_module_data_out[4] ,
    \sw_450_module_data_out[3] ,
    \sw_450_module_data_out[2] ,
    \sw_450_module_data_out[1] ,
    \sw_450_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_451 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_451_module_data_in[7] ,
    \sw_451_module_data_in[6] ,
    \sw_451_module_data_in[5] ,
    \sw_451_module_data_in[4] ,
    \sw_451_module_data_in[3] ,
    \sw_451_module_data_in[2] ,
    \sw_451_module_data_in[1] ,
    \sw_451_module_data_in[0] }),
    .io_out({\sw_451_module_data_out[7] ,
    \sw_451_module_data_out[6] ,
    \sw_451_module_data_out[5] ,
    \sw_451_module_data_out[4] ,
    \sw_451_module_data_out[3] ,
    \sw_451_module_data_out[2] ,
    \sw_451_module_data_out[1] ,
    \sw_451_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_452 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_452_module_data_in[7] ,
    \sw_452_module_data_in[6] ,
    \sw_452_module_data_in[5] ,
    \sw_452_module_data_in[4] ,
    \sw_452_module_data_in[3] ,
    \sw_452_module_data_in[2] ,
    \sw_452_module_data_in[1] ,
    \sw_452_module_data_in[0] }),
    .io_out({\sw_452_module_data_out[7] ,
    \sw_452_module_data_out[6] ,
    \sw_452_module_data_out[5] ,
    \sw_452_module_data_out[4] ,
    \sw_452_module_data_out[3] ,
    \sw_452_module_data_out[2] ,
    \sw_452_module_data_out[1] ,
    \sw_452_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_453 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_453_module_data_in[7] ,
    \sw_453_module_data_in[6] ,
    \sw_453_module_data_in[5] ,
    \sw_453_module_data_in[4] ,
    \sw_453_module_data_in[3] ,
    \sw_453_module_data_in[2] ,
    \sw_453_module_data_in[1] ,
    \sw_453_module_data_in[0] }),
    .io_out({\sw_453_module_data_out[7] ,
    \sw_453_module_data_out[6] ,
    \sw_453_module_data_out[5] ,
    \sw_453_module_data_out[4] ,
    \sw_453_module_data_out[3] ,
    \sw_453_module_data_out[2] ,
    \sw_453_module_data_out[1] ,
    \sw_453_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_454 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_454_module_data_in[7] ,
    \sw_454_module_data_in[6] ,
    \sw_454_module_data_in[5] ,
    \sw_454_module_data_in[4] ,
    \sw_454_module_data_in[3] ,
    \sw_454_module_data_in[2] ,
    \sw_454_module_data_in[1] ,
    \sw_454_module_data_in[0] }),
    .io_out({\sw_454_module_data_out[7] ,
    \sw_454_module_data_out[6] ,
    \sw_454_module_data_out[5] ,
    \sw_454_module_data_out[4] ,
    \sw_454_module_data_out[3] ,
    \sw_454_module_data_out[2] ,
    \sw_454_module_data_out[1] ,
    \sw_454_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_455 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_455_module_data_in[7] ,
    \sw_455_module_data_in[6] ,
    \sw_455_module_data_in[5] ,
    \sw_455_module_data_in[4] ,
    \sw_455_module_data_in[3] ,
    \sw_455_module_data_in[2] ,
    \sw_455_module_data_in[1] ,
    \sw_455_module_data_in[0] }),
    .io_out({\sw_455_module_data_out[7] ,
    \sw_455_module_data_out[6] ,
    \sw_455_module_data_out[5] ,
    \sw_455_module_data_out[4] ,
    \sw_455_module_data_out[3] ,
    \sw_455_module_data_out[2] ,
    \sw_455_module_data_out[1] ,
    \sw_455_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_456 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_456_module_data_in[7] ,
    \sw_456_module_data_in[6] ,
    \sw_456_module_data_in[5] ,
    \sw_456_module_data_in[4] ,
    \sw_456_module_data_in[3] ,
    \sw_456_module_data_in[2] ,
    \sw_456_module_data_in[1] ,
    \sw_456_module_data_in[0] }),
    .io_out({\sw_456_module_data_out[7] ,
    \sw_456_module_data_out[6] ,
    \sw_456_module_data_out[5] ,
    \sw_456_module_data_out[4] ,
    \sw_456_module_data_out[3] ,
    \sw_456_module_data_out[2] ,
    \sw_456_module_data_out[1] ,
    \sw_456_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_457 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_457_module_data_in[7] ,
    \sw_457_module_data_in[6] ,
    \sw_457_module_data_in[5] ,
    \sw_457_module_data_in[4] ,
    \sw_457_module_data_in[3] ,
    \sw_457_module_data_in[2] ,
    \sw_457_module_data_in[1] ,
    \sw_457_module_data_in[0] }),
    .io_out({\sw_457_module_data_out[7] ,
    \sw_457_module_data_out[6] ,
    \sw_457_module_data_out[5] ,
    \sw_457_module_data_out[4] ,
    \sw_457_module_data_out[3] ,
    \sw_457_module_data_out[2] ,
    \sw_457_module_data_out[1] ,
    \sw_457_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_458 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_458_module_data_in[7] ,
    \sw_458_module_data_in[6] ,
    \sw_458_module_data_in[5] ,
    \sw_458_module_data_in[4] ,
    \sw_458_module_data_in[3] ,
    \sw_458_module_data_in[2] ,
    \sw_458_module_data_in[1] ,
    \sw_458_module_data_in[0] }),
    .io_out({\sw_458_module_data_out[7] ,
    \sw_458_module_data_out[6] ,
    \sw_458_module_data_out[5] ,
    \sw_458_module_data_out[4] ,
    \sw_458_module_data_out[3] ,
    \sw_458_module_data_out[2] ,
    \sw_458_module_data_out[1] ,
    \sw_458_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_459 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_459_module_data_in[7] ,
    \sw_459_module_data_in[6] ,
    \sw_459_module_data_in[5] ,
    \sw_459_module_data_in[4] ,
    \sw_459_module_data_in[3] ,
    \sw_459_module_data_in[2] ,
    \sw_459_module_data_in[1] ,
    \sw_459_module_data_in[0] }),
    .io_out({\sw_459_module_data_out[7] ,
    \sw_459_module_data_out[6] ,
    \sw_459_module_data_out[5] ,
    \sw_459_module_data_out[4] ,
    \sw_459_module_data_out[3] ,
    \sw_459_module_data_out[2] ,
    \sw_459_module_data_out[1] ,
    \sw_459_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_46 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_046_module_data_in[7] ,
    \sw_046_module_data_in[6] ,
    \sw_046_module_data_in[5] ,
    \sw_046_module_data_in[4] ,
    \sw_046_module_data_in[3] ,
    \sw_046_module_data_in[2] ,
    \sw_046_module_data_in[1] ,
    \sw_046_module_data_in[0] }),
    .io_out({\sw_046_module_data_out[7] ,
    \sw_046_module_data_out[6] ,
    \sw_046_module_data_out[5] ,
    \sw_046_module_data_out[4] ,
    \sw_046_module_data_out[3] ,
    \sw_046_module_data_out[2] ,
    \sw_046_module_data_out[1] ,
    \sw_046_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_460 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_460_module_data_in[7] ,
    \sw_460_module_data_in[6] ,
    \sw_460_module_data_in[5] ,
    \sw_460_module_data_in[4] ,
    \sw_460_module_data_in[3] ,
    \sw_460_module_data_in[2] ,
    \sw_460_module_data_in[1] ,
    \sw_460_module_data_in[0] }),
    .io_out({\sw_460_module_data_out[7] ,
    \sw_460_module_data_out[6] ,
    \sw_460_module_data_out[5] ,
    \sw_460_module_data_out[4] ,
    \sw_460_module_data_out[3] ,
    \sw_460_module_data_out[2] ,
    \sw_460_module_data_out[1] ,
    \sw_460_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_461 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_461_module_data_in[7] ,
    \sw_461_module_data_in[6] ,
    \sw_461_module_data_in[5] ,
    \sw_461_module_data_in[4] ,
    \sw_461_module_data_in[3] ,
    \sw_461_module_data_in[2] ,
    \sw_461_module_data_in[1] ,
    \sw_461_module_data_in[0] }),
    .io_out({\sw_461_module_data_out[7] ,
    \sw_461_module_data_out[6] ,
    \sw_461_module_data_out[5] ,
    \sw_461_module_data_out[4] ,
    \sw_461_module_data_out[3] ,
    \sw_461_module_data_out[2] ,
    \sw_461_module_data_out[1] ,
    \sw_461_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_462 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_462_module_data_in[7] ,
    \sw_462_module_data_in[6] ,
    \sw_462_module_data_in[5] ,
    \sw_462_module_data_in[4] ,
    \sw_462_module_data_in[3] ,
    \sw_462_module_data_in[2] ,
    \sw_462_module_data_in[1] ,
    \sw_462_module_data_in[0] }),
    .io_out({\sw_462_module_data_out[7] ,
    \sw_462_module_data_out[6] ,
    \sw_462_module_data_out[5] ,
    \sw_462_module_data_out[4] ,
    \sw_462_module_data_out[3] ,
    \sw_462_module_data_out[2] ,
    \sw_462_module_data_out[1] ,
    \sw_462_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_463 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_463_module_data_in[7] ,
    \sw_463_module_data_in[6] ,
    \sw_463_module_data_in[5] ,
    \sw_463_module_data_in[4] ,
    \sw_463_module_data_in[3] ,
    \sw_463_module_data_in[2] ,
    \sw_463_module_data_in[1] ,
    \sw_463_module_data_in[0] }),
    .io_out({\sw_463_module_data_out[7] ,
    \sw_463_module_data_out[6] ,
    \sw_463_module_data_out[5] ,
    \sw_463_module_data_out[4] ,
    \sw_463_module_data_out[3] ,
    \sw_463_module_data_out[2] ,
    \sw_463_module_data_out[1] ,
    \sw_463_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_464 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_464_module_data_in[7] ,
    \sw_464_module_data_in[6] ,
    \sw_464_module_data_in[5] ,
    \sw_464_module_data_in[4] ,
    \sw_464_module_data_in[3] ,
    \sw_464_module_data_in[2] ,
    \sw_464_module_data_in[1] ,
    \sw_464_module_data_in[0] }),
    .io_out({\sw_464_module_data_out[7] ,
    \sw_464_module_data_out[6] ,
    \sw_464_module_data_out[5] ,
    \sw_464_module_data_out[4] ,
    \sw_464_module_data_out[3] ,
    \sw_464_module_data_out[2] ,
    \sw_464_module_data_out[1] ,
    \sw_464_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_465 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_465_module_data_in[7] ,
    \sw_465_module_data_in[6] ,
    \sw_465_module_data_in[5] ,
    \sw_465_module_data_in[4] ,
    \sw_465_module_data_in[3] ,
    \sw_465_module_data_in[2] ,
    \sw_465_module_data_in[1] ,
    \sw_465_module_data_in[0] }),
    .io_out({\sw_465_module_data_out[7] ,
    \sw_465_module_data_out[6] ,
    \sw_465_module_data_out[5] ,
    \sw_465_module_data_out[4] ,
    \sw_465_module_data_out[3] ,
    \sw_465_module_data_out[2] ,
    \sw_465_module_data_out[1] ,
    \sw_465_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_466 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_466_module_data_in[7] ,
    \sw_466_module_data_in[6] ,
    \sw_466_module_data_in[5] ,
    \sw_466_module_data_in[4] ,
    \sw_466_module_data_in[3] ,
    \sw_466_module_data_in[2] ,
    \sw_466_module_data_in[1] ,
    \sw_466_module_data_in[0] }),
    .io_out({\sw_466_module_data_out[7] ,
    \sw_466_module_data_out[6] ,
    \sw_466_module_data_out[5] ,
    \sw_466_module_data_out[4] ,
    \sw_466_module_data_out[3] ,
    \sw_466_module_data_out[2] ,
    \sw_466_module_data_out[1] ,
    \sw_466_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_467 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_467_module_data_in[7] ,
    \sw_467_module_data_in[6] ,
    \sw_467_module_data_in[5] ,
    \sw_467_module_data_in[4] ,
    \sw_467_module_data_in[3] ,
    \sw_467_module_data_in[2] ,
    \sw_467_module_data_in[1] ,
    \sw_467_module_data_in[0] }),
    .io_out({\sw_467_module_data_out[7] ,
    \sw_467_module_data_out[6] ,
    \sw_467_module_data_out[5] ,
    \sw_467_module_data_out[4] ,
    \sw_467_module_data_out[3] ,
    \sw_467_module_data_out[2] ,
    \sw_467_module_data_out[1] ,
    \sw_467_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_468 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_468_module_data_in[7] ,
    \sw_468_module_data_in[6] ,
    \sw_468_module_data_in[5] ,
    \sw_468_module_data_in[4] ,
    \sw_468_module_data_in[3] ,
    \sw_468_module_data_in[2] ,
    \sw_468_module_data_in[1] ,
    \sw_468_module_data_in[0] }),
    .io_out({\sw_468_module_data_out[7] ,
    \sw_468_module_data_out[6] ,
    \sw_468_module_data_out[5] ,
    \sw_468_module_data_out[4] ,
    \sw_468_module_data_out[3] ,
    \sw_468_module_data_out[2] ,
    \sw_468_module_data_out[1] ,
    \sw_468_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_469 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_469_module_data_in[7] ,
    \sw_469_module_data_in[6] ,
    \sw_469_module_data_in[5] ,
    \sw_469_module_data_in[4] ,
    \sw_469_module_data_in[3] ,
    \sw_469_module_data_in[2] ,
    \sw_469_module_data_in[1] ,
    \sw_469_module_data_in[0] }),
    .io_out({\sw_469_module_data_out[7] ,
    \sw_469_module_data_out[6] ,
    \sw_469_module_data_out[5] ,
    \sw_469_module_data_out[4] ,
    \sw_469_module_data_out[3] ,
    \sw_469_module_data_out[2] ,
    \sw_469_module_data_out[1] ,
    \sw_469_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_47 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_047_module_data_in[7] ,
    \sw_047_module_data_in[6] ,
    \sw_047_module_data_in[5] ,
    \sw_047_module_data_in[4] ,
    \sw_047_module_data_in[3] ,
    \sw_047_module_data_in[2] ,
    \sw_047_module_data_in[1] ,
    \sw_047_module_data_in[0] }),
    .io_out({\sw_047_module_data_out[7] ,
    \sw_047_module_data_out[6] ,
    \sw_047_module_data_out[5] ,
    \sw_047_module_data_out[4] ,
    \sw_047_module_data_out[3] ,
    \sw_047_module_data_out[2] ,
    \sw_047_module_data_out[1] ,
    \sw_047_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_470 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_470_module_data_in[7] ,
    \sw_470_module_data_in[6] ,
    \sw_470_module_data_in[5] ,
    \sw_470_module_data_in[4] ,
    \sw_470_module_data_in[3] ,
    \sw_470_module_data_in[2] ,
    \sw_470_module_data_in[1] ,
    \sw_470_module_data_in[0] }),
    .io_out({\sw_470_module_data_out[7] ,
    \sw_470_module_data_out[6] ,
    \sw_470_module_data_out[5] ,
    \sw_470_module_data_out[4] ,
    \sw_470_module_data_out[3] ,
    \sw_470_module_data_out[2] ,
    \sw_470_module_data_out[1] ,
    \sw_470_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_471 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_471_module_data_in[7] ,
    \sw_471_module_data_in[6] ,
    \sw_471_module_data_in[5] ,
    \sw_471_module_data_in[4] ,
    \sw_471_module_data_in[3] ,
    \sw_471_module_data_in[2] ,
    \sw_471_module_data_in[1] ,
    \sw_471_module_data_in[0] }),
    .io_out({\sw_471_module_data_out[7] ,
    \sw_471_module_data_out[6] ,
    \sw_471_module_data_out[5] ,
    \sw_471_module_data_out[4] ,
    \sw_471_module_data_out[3] ,
    \sw_471_module_data_out[2] ,
    \sw_471_module_data_out[1] ,
    \sw_471_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_472 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_472_module_data_in[7] ,
    \sw_472_module_data_in[6] ,
    \sw_472_module_data_in[5] ,
    \sw_472_module_data_in[4] ,
    \sw_472_module_data_in[3] ,
    \sw_472_module_data_in[2] ,
    \sw_472_module_data_in[1] ,
    \sw_472_module_data_in[0] }),
    .io_out({\sw_472_module_data_out[7] ,
    \sw_472_module_data_out[6] ,
    \sw_472_module_data_out[5] ,
    \sw_472_module_data_out[4] ,
    \sw_472_module_data_out[3] ,
    \sw_472_module_data_out[2] ,
    \sw_472_module_data_out[1] ,
    \sw_472_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_48 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_048_module_data_in[7] ,
    \sw_048_module_data_in[6] ,
    \sw_048_module_data_in[5] ,
    \sw_048_module_data_in[4] ,
    \sw_048_module_data_in[3] ,
    \sw_048_module_data_in[2] ,
    \sw_048_module_data_in[1] ,
    \sw_048_module_data_in[0] }),
    .io_out({\sw_048_module_data_out[7] ,
    \sw_048_module_data_out[6] ,
    \sw_048_module_data_out[5] ,
    \sw_048_module_data_out[4] ,
    \sw_048_module_data_out[3] ,
    \sw_048_module_data_out[2] ,
    \sw_048_module_data_out[1] ,
    \sw_048_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_49 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_049_module_data_in[7] ,
    \sw_049_module_data_in[6] ,
    \sw_049_module_data_in[5] ,
    \sw_049_module_data_in[4] ,
    \sw_049_module_data_in[3] ,
    \sw_049_module_data_in[2] ,
    \sw_049_module_data_in[1] ,
    \sw_049_module_data_in[0] }),
    .io_out({\sw_049_module_data_out[7] ,
    \sw_049_module_data_out[6] ,
    \sw_049_module_data_out[5] ,
    \sw_049_module_data_out[4] ,
    \sw_049_module_data_out[3] ,
    \sw_049_module_data_out[2] ,
    \sw_049_module_data_out[1] ,
    \sw_049_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_50 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_050_module_data_in[7] ,
    \sw_050_module_data_in[6] ,
    \sw_050_module_data_in[5] ,
    \sw_050_module_data_in[4] ,
    \sw_050_module_data_in[3] ,
    \sw_050_module_data_in[2] ,
    \sw_050_module_data_in[1] ,
    \sw_050_module_data_in[0] }),
    .io_out({\sw_050_module_data_out[7] ,
    \sw_050_module_data_out[6] ,
    \sw_050_module_data_out[5] ,
    \sw_050_module_data_out[4] ,
    \sw_050_module_data_out[3] ,
    \sw_050_module_data_out[2] ,
    \sw_050_module_data_out[1] ,
    \sw_050_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_51 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_051_module_data_in[7] ,
    \sw_051_module_data_in[6] ,
    \sw_051_module_data_in[5] ,
    \sw_051_module_data_in[4] ,
    \sw_051_module_data_in[3] ,
    \sw_051_module_data_in[2] ,
    \sw_051_module_data_in[1] ,
    \sw_051_module_data_in[0] }),
    .io_out({\sw_051_module_data_out[7] ,
    \sw_051_module_data_out[6] ,
    \sw_051_module_data_out[5] ,
    \sw_051_module_data_out[4] ,
    \sw_051_module_data_out[3] ,
    \sw_051_module_data_out[2] ,
    \sw_051_module_data_out[1] ,
    \sw_051_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_52 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_052_module_data_in[7] ,
    \sw_052_module_data_in[6] ,
    \sw_052_module_data_in[5] ,
    \sw_052_module_data_in[4] ,
    \sw_052_module_data_in[3] ,
    \sw_052_module_data_in[2] ,
    \sw_052_module_data_in[1] ,
    \sw_052_module_data_in[0] }),
    .io_out({\sw_052_module_data_out[7] ,
    \sw_052_module_data_out[6] ,
    \sw_052_module_data_out[5] ,
    \sw_052_module_data_out[4] ,
    \sw_052_module_data_out[3] ,
    \sw_052_module_data_out[2] ,
    \sw_052_module_data_out[1] ,
    \sw_052_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_53 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_053_module_data_in[7] ,
    \sw_053_module_data_in[6] ,
    \sw_053_module_data_in[5] ,
    \sw_053_module_data_in[4] ,
    \sw_053_module_data_in[3] ,
    \sw_053_module_data_in[2] ,
    \sw_053_module_data_in[1] ,
    \sw_053_module_data_in[0] }),
    .io_out({\sw_053_module_data_out[7] ,
    \sw_053_module_data_out[6] ,
    \sw_053_module_data_out[5] ,
    \sw_053_module_data_out[4] ,
    \sw_053_module_data_out[3] ,
    \sw_053_module_data_out[2] ,
    \sw_053_module_data_out[1] ,
    \sw_053_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_54 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_054_module_data_in[7] ,
    \sw_054_module_data_in[6] ,
    \sw_054_module_data_in[5] ,
    \sw_054_module_data_in[4] ,
    \sw_054_module_data_in[3] ,
    \sw_054_module_data_in[2] ,
    \sw_054_module_data_in[1] ,
    \sw_054_module_data_in[0] }),
    .io_out({\sw_054_module_data_out[7] ,
    \sw_054_module_data_out[6] ,
    \sw_054_module_data_out[5] ,
    \sw_054_module_data_out[4] ,
    \sw_054_module_data_out[3] ,
    \sw_054_module_data_out[2] ,
    \sw_054_module_data_out[1] ,
    \sw_054_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_55 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_055_module_data_in[7] ,
    \sw_055_module_data_in[6] ,
    \sw_055_module_data_in[5] ,
    \sw_055_module_data_in[4] ,
    \sw_055_module_data_in[3] ,
    \sw_055_module_data_in[2] ,
    \sw_055_module_data_in[1] ,
    \sw_055_module_data_in[0] }),
    .io_out({\sw_055_module_data_out[7] ,
    \sw_055_module_data_out[6] ,
    \sw_055_module_data_out[5] ,
    \sw_055_module_data_out[4] ,
    \sw_055_module_data_out[3] ,
    \sw_055_module_data_out[2] ,
    \sw_055_module_data_out[1] ,
    \sw_055_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_56 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_056_module_data_in[7] ,
    \sw_056_module_data_in[6] ,
    \sw_056_module_data_in[5] ,
    \sw_056_module_data_in[4] ,
    \sw_056_module_data_in[3] ,
    \sw_056_module_data_in[2] ,
    \sw_056_module_data_in[1] ,
    \sw_056_module_data_in[0] }),
    .io_out({\sw_056_module_data_out[7] ,
    \sw_056_module_data_out[6] ,
    \sw_056_module_data_out[5] ,
    \sw_056_module_data_out[4] ,
    \sw_056_module_data_out[3] ,
    \sw_056_module_data_out[2] ,
    \sw_056_module_data_out[1] ,
    \sw_056_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_57 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_057_module_data_in[7] ,
    \sw_057_module_data_in[6] ,
    \sw_057_module_data_in[5] ,
    \sw_057_module_data_in[4] ,
    \sw_057_module_data_in[3] ,
    \sw_057_module_data_in[2] ,
    \sw_057_module_data_in[1] ,
    \sw_057_module_data_in[0] }),
    .io_out({\sw_057_module_data_out[7] ,
    \sw_057_module_data_out[6] ,
    \sw_057_module_data_out[5] ,
    \sw_057_module_data_out[4] ,
    \sw_057_module_data_out[3] ,
    \sw_057_module_data_out[2] ,
    \sw_057_module_data_out[1] ,
    \sw_057_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_58 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_058_module_data_in[7] ,
    \sw_058_module_data_in[6] ,
    \sw_058_module_data_in[5] ,
    \sw_058_module_data_in[4] ,
    \sw_058_module_data_in[3] ,
    \sw_058_module_data_in[2] ,
    \sw_058_module_data_in[1] ,
    \sw_058_module_data_in[0] }),
    .io_out({\sw_058_module_data_out[7] ,
    \sw_058_module_data_out[6] ,
    \sw_058_module_data_out[5] ,
    \sw_058_module_data_out[4] ,
    \sw_058_module_data_out[3] ,
    \sw_058_module_data_out[2] ,
    \sw_058_module_data_out[1] ,
    \sw_058_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_59 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_059_module_data_in[7] ,
    \sw_059_module_data_in[6] ,
    \sw_059_module_data_in[5] ,
    \sw_059_module_data_in[4] ,
    \sw_059_module_data_in[3] ,
    \sw_059_module_data_in[2] ,
    \sw_059_module_data_in[1] ,
    \sw_059_module_data_in[0] }),
    .io_out({\sw_059_module_data_out[7] ,
    \sw_059_module_data_out[6] ,
    \sw_059_module_data_out[5] ,
    \sw_059_module_data_out[4] ,
    \sw_059_module_data_out[3] ,
    \sw_059_module_data_out[2] ,
    \sw_059_module_data_out[1] ,
    \sw_059_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_60 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_060_module_data_in[7] ,
    \sw_060_module_data_in[6] ,
    \sw_060_module_data_in[5] ,
    \sw_060_module_data_in[4] ,
    \sw_060_module_data_in[3] ,
    \sw_060_module_data_in[2] ,
    \sw_060_module_data_in[1] ,
    \sw_060_module_data_in[0] }),
    .io_out({\sw_060_module_data_out[7] ,
    \sw_060_module_data_out[6] ,
    \sw_060_module_data_out[5] ,
    \sw_060_module_data_out[4] ,
    \sw_060_module_data_out[3] ,
    \sw_060_module_data_out[2] ,
    \sw_060_module_data_out[1] ,
    \sw_060_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_61 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_061_module_data_in[7] ,
    \sw_061_module_data_in[6] ,
    \sw_061_module_data_in[5] ,
    \sw_061_module_data_in[4] ,
    \sw_061_module_data_in[3] ,
    \sw_061_module_data_in[2] ,
    \sw_061_module_data_in[1] ,
    \sw_061_module_data_in[0] }),
    .io_out({\sw_061_module_data_out[7] ,
    \sw_061_module_data_out[6] ,
    \sw_061_module_data_out[5] ,
    \sw_061_module_data_out[4] ,
    \sw_061_module_data_out[3] ,
    \sw_061_module_data_out[2] ,
    \sw_061_module_data_out[1] ,
    \sw_061_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_62 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_062_module_data_in[7] ,
    \sw_062_module_data_in[6] ,
    \sw_062_module_data_in[5] ,
    \sw_062_module_data_in[4] ,
    \sw_062_module_data_in[3] ,
    \sw_062_module_data_in[2] ,
    \sw_062_module_data_in[1] ,
    \sw_062_module_data_in[0] }),
    .io_out({\sw_062_module_data_out[7] ,
    \sw_062_module_data_out[6] ,
    \sw_062_module_data_out[5] ,
    \sw_062_module_data_out[4] ,
    \sw_062_module_data_out[3] ,
    \sw_062_module_data_out[2] ,
    \sw_062_module_data_out[1] ,
    \sw_062_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_63 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_063_module_data_in[7] ,
    \sw_063_module_data_in[6] ,
    \sw_063_module_data_in[5] ,
    \sw_063_module_data_in[4] ,
    \sw_063_module_data_in[3] ,
    \sw_063_module_data_in[2] ,
    \sw_063_module_data_in[1] ,
    \sw_063_module_data_in[0] }),
    .io_out({\sw_063_module_data_out[7] ,
    \sw_063_module_data_out[6] ,
    \sw_063_module_data_out[5] ,
    \sw_063_module_data_out[4] ,
    \sw_063_module_data_out[3] ,
    \sw_063_module_data_out[2] ,
    \sw_063_module_data_out[1] ,
    \sw_063_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_64 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_064_module_data_in[7] ,
    \sw_064_module_data_in[6] ,
    \sw_064_module_data_in[5] ,
    \sw_064_module_data_in[4] ,
    \sw_064_module_data_in[3] ,
    \sw_064_module_data_in[2] ,
    \sw_064_module_data_in[1] ,
    \sw_064_module_data_in[0] }),
    .io_out({\sw_064_module_data_out[7] ,
    \sw_064_module_data_out[6] ,
    \sw_064_module_data_out[5] ,
    \sw_064_module_data_out[4] ,
    \sw_064_module_data_out[3] ,
    \sw_064_module_data_out[2] ,
    \sw_064_module_data_out[1] ,
    \sw_064_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_65 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_065_module_data_in[7] ,
    \sw_065_module_data_in[6] ,
    \sw_065_module_data_in[5] ,
    \sw_065_module_data_in[4] ,
    \sw_065_module_data_in[3] ,
    \sw_065_module_data_in[2] ,
    \sw_065_module_data_in[1] ,
    \sw_065_module_data_in[0] }),
    .io_out({\sw_065_module_data_out[7] ,
    \sw_065_module_data_out[6] ,
    \sw_065_module_data_out[5] ,
    \sw_065_module_data_out[4] ,
    \sw_065_module_data_out[3] ,
    \sw_065_module_data_out[2] ,
    \sw_065_module_data_out[1] ,
    \sw_065_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_66 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_066_module_data_in[7] ,
    \sw_066_module_data_in[6] ,
    \sw_066_module_data_in[5] ,
    \sw_066_module_data_in[4] ,
    \sw_066_module_data_in[3] ,
    \sw_066_module_data_in[2] ,
    \sw_066_module_data_in[1] ,
    \sw_066_module_data_in[0] }),
    .io_out({\sw_066_module_data_out[7] ,
    \sw_066_module_data_out[6] ,
    \sw_066_module_data_out[5] ,
    \sw_066_module_data_out[4] ,
    \sw_066_module_data_out[3] ,
    \sw_066_module_data_out[2] ,
    \sw_066_module_data_out[1] ,
    \sw_066_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_67 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_067_module_data_in[7] ,
    \sw_067_module_data_in[6] ,
    \sw_067_module_data_in[5] ,
    \sw_067_module_data_in[4] ,
    \sw_067_module_data_in[3] ,
    \sw_067_module_data_in[2] ,
    \sw_067_module_data_in[1] ,
    \sw_067_module_data_in[0] }),
    .io_out({\sw_067_module_data_out[7] ,
    \sw_067_module_data_out[6] ,
    \sw_067_module_data_out[5] ,
    \sw_067_module_data_out[4] ,
    \sw_067_module_data_out[3] ,
    \sw_067_module_data_out[2] ,
    \sw_067_module_data_out[1] ,
    \sw_067_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_68 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_068_module_data_in[7] ,
    \sw_068_module_data_in[6] ,
    \sw_068_module_data_in[5] ,
    \sw_068_module_data_in[4] ,
    \sw_068_module_data_in[3] ,
    \sw_068_module_data_in[2] ,
    \sw_068_module_data_in[1] ,
    \sw_068_module_data_in[0] }),
    .io_out({\sw_068_module_data_out[7] ,
    \sw_068_module_data_out[6] ,
    \sw_068_module_data_out[5] ,
    \sw_068_module_data_out[4] ,
    \sw_068_module_data_out[3] ,
    \sw_068_module_data_out[2] ,
    \sw_068_module_data_out[1] ,
    \sw_068_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_69 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_069_module_data_in[7] ,
    \sw_069_module_data_in[6] ,
    \sw_069_module_data_in[5] ,
    \sw_069_module_data_in[4] ,
    \sw_069_module_data_in[3] ,
    \sw_069_module_data_in[2] ,
    \sw_069_module_data_in[1] ,
    \sw_069_module_data_in[0] }),
    .io_out({\sw_069_module_data_out[7] ,
    \sw_069_module_data_out[6] ,
    \sw_069_module_data_out[5] ,
    \sw_069_module_data_out[4] ,
    \sw_069_module_data_out[3] ,
    \sw_069_module_data_out[2] ,
    \sw_069_module_data_out[1] ,
    \sw_069_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_70 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_070_module_data_in[7] ,
    \sw_070_module_data_in[6] ,
    \sw_070_module_data_in[5] ,
    \sw_070_module_data_in[4] ,
    \sw_070_module_data_in[3] ,
    \sw_070_module_data_in[2] ,
    \sw_070_module_data_in[1] ,
    \sw_070_module_data_in[0] }),
    .io_out({\sw_070_module_data_out[7] ,
    \sw_070_module_data_out[6] ,
    \sw_070_module_data_out[5] ,
    \sw_070_module_data_out[4] ,
    \sw_070_module_data_out[3] ,
    \sw_070_module_data_out[2] ,
    \sw_070_module_data_out[1] ,
    \sw_070_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_71 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_071_module_data_in[7] ,
    \sw_071_module_data_in[6] ,
    \sw_071_module_data_in[5] ,
    \sw_071_module_data_in[4] ,
    \sw_071_module_data_in[3] ,
    \sw_071_module_data_in[2] ,
    \sw_071_module_data_in[1] ,
    \sw_071_module_data_in[0] }),
    .io_out({\sw_071_module_data_out[7] ,
    \sw_071_module_data_out[6] ,
    \sw_071_module_data_out[5] ,
    \sw_071_module_data_out[4] ,
    \sw_071_module_data_out[3] ,
    \sw_071_module_data_out[2] ,
    \sw_071_module_data_out[1] ,
    \sw_071_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_72 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_072_module_data_in[7] ,
    \sw_072_module_data_in[6] ,
    \sw_072_module_data_in[5] ,
    \sw_072_module_data_in[4] ,
    \sw_072_module_data_in[3] ,
    \sw_072_module_data_in[2] ,
    \sw_072_module_data_in[1] ,
    \sw_072_module_data_in[0] }),
    .io_out({\sw_072_module_data_out[7] ,
    \sw_072_module_data_out[6] ,
    \sw_072_module_data_out[5] ,
    \sw_072_module_data_out[4] ,
    \sw_072_module_data_out[3] ,
    \sw_072_module_data_out[2] ,
    \sw_072_module_data_out[1] ,
    \sw_072_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_73 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_073_module_data_in[7] ,
    \sw_073_module_data_in[6] ,
    \sw_073_module_data_in[5] ,
    \sw_073_module_data_in[4] ,
    \sw_073_module_data_in[3] ,
    \sw_073_module_data_in[2] ,
    \sw_073_module_data_in[1] ,
    \sw_073_module_data_in[0] }),
    .io_out({\sw_073_module_data_out[7] ,
    \sw_073_module_data_out[6] ,
    \sw_073_module_data_out[5] ,
    \sw_073_module_data_out[4] ,
    \sw_073_module_data_out[3] ,
    \sw_073_module_data_out[2] ,
    \sw_073_module_data_out[1] ,
    \sw_073_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_74 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_074_module_data_in[7] ,
    \sw_074_module_data_in[6] ,
    \sw_074_module_data_in[5] ,
    \sw_074_module_data_in[4] ,
    \sw_074_module_data_in[3] ,
    \sw_074_module_data_in[2] ,
    \sw_074_module_data_in[1] ,
    \sw_074_module_data_in[0] }),
    .io_out({\sw_074_module_data_out[7] ,
    \sw_074_module_data_out[6] ,
    \sw_074_module_data_out[5] ,
    \sw_074_module_data_out[4] ,
    \sw_074_module_data_out[3] ,
    \sw_074_module_data_out[2] ,
    \sw_074_module_data_out[1] ,
    \sw_074_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_75 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_075_module_data_in[7] ,
    \sw_075_module_data_in[6] ,
    \sw_075_module_data_in[5] ,
    \sw_075_module_data_in[4] ,
    \sw_075_module_data_in[3] ,
    \sw_075_module_data_in[2] ,
    \sw_075_module_data_in[1] ,
    \sw_075_module_data_in[0] }),
    .io_out({\sw_075_module_data_out[7] ,
    \sw_075_module_data_out[6] ,
    \sw_075_module_data_out[5] ,
    \sw_075_module_data_out[4] ,
    \sw_075_module_data_out[3] ,
    \sw_075_module_data_out[2] ,
    \sw_075_module_data_out[1] ,
    \sw_075_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_76 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_076_module_data_in[7] ,
    \sw_076_module_data_in[6] ,
    \sw_076_module_data_in[5] ,
    \sw_076_module_data_in[4] ,
    \sw_076_module_data_in[3] ,
    \sw_076_module_data_in[2] ,
    \sw_076_module_data_in[1] ,
    \sw_076_module_data_in[0] }),
    .io_out({\sw_076_module_data_out[7] ,
    \sw_076_module_data_out[6] ,
    \sw_076_module_data_out[5] ,
    \sw_076_module_data_out[4] ,
    \sw_076_module_data_out[3] ,
    \sw_076_module_data_out[2] ,
    \sw_076_module_data_out[1] ,
    \sw_076_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_77 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_077_module_data_in[7] ,
    \sw_077_module_data_in[6] ,
    \sw_077_module_data_in[5] ,
    \sw_077_module_data_in[4] ,
    \sw_077_module_data_in[3] ,
    \sw_077_module_data_in[2] ,
    \sw_077_module_data_in[1] ,
    \sw_077_module_data_in[0] }),
    .io_out({\sw_077_module_data_out[7] ,
    \sw_077_module_data_out[6] ,
    \sw_077_module_data_out[5] ,
    \sw_077_module_data_out[4] ,
    \sw_077_module_data_out[3] ,
    \sw_077_module_data_out[2] ,
    \sw_077_module_data_out[1] ,
    \sw_077_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_78 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_078_module_data_in[7] ,
    \sw_078_module_data_in[6] ,
    \sw_078_module_data_in[5] ,
    \sw_078_module_data_in[4] ,
    \sw_078_module_data_in[3] ,
    \sw_078_module_data_in[2] ,
    \sw_078_module_data_in[1] ,
    \sw_078_module_data_in[0] }),
    .io_out({\sw_078_module_data_out[7] ,
    \sw_078_module_data_out[6] ,
    \sw_078_module_data_out[5] ,
    \sw_078_module_data_out[4] ,
    \sw_078_module_data_out[3] ,
    \sw_078_module_data_out[2] ,
    \sw_078_module_data_out[1] ,
    \sw_078_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_79 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_079_module_data_in[7] ,
    \sw_079_module_data_in[6] ,
    \sw_079_module_data_in[5] ,
    \sw_079_module_data_in[4] ,
    \sw_079_module_data_in[3] ,
    \sw_079_module_data_in[2] ,
    \sw_079_module_data_in[1] ,
    \sw_079_module_data_in[0] }),
    .io_out({\sw_079_module_data_out[7] ,
    \sw_079_module_data_out[6] ,
    \sw_079_module_data_out[5] ,
    \sw_079_module_data_out[4] ,
    \sw_079_module_data_out[3] ,
    \sw_079_module_data_out[2] ,
    \sw_079_module_data_out[1] ,
    \sw_079_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_80 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_080_module_data_in[7] ,
    \sw_080_module_data_in[6] ,
    \sw_080_module_data_in[5] ,
    \sw_080_module_data_in[4] ,
    \sw_080_module_data_in[3] ,
    \sw_080_module_data_in[2] ,
    \sw_080_module_data_in[1] ,
    \sw_080_module_data_in[0] }),
    .io_out({\sw_080_module_data_out[7] ,
    \sw_080_module_data_out[6] ,
    \sw_080_module_data_out[5] ,
    \sw_080_module_data_out[4] ,
    \sw_080_module_data_out[3] ,
    \sw_080_module_data_out[2] ,
    \sw_080_module_data_out[1] ,
    \sw_080_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_81 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_081_module_data_in[7] ,
    \sw_081_module_data_in[6] ,
    \sw_081_module_data_in[5] ,
    \sw_081_module_data_in[4] ,
    \sw_081_module_data_in[3] ,
    \sw_081_module_data_in[2] ,
    \sw_081_module_data_in[1] ,
    \sw_081_module_data_in[0] }),
    .io_out({\sw_081_module_data_out[7] ,
    \sw_081_module_data_out[6] ,
    \sw_081_module_data_out[5] ,
    \sw_081_module_data_out[4] ,
    \sw_081_module_data_out[3] ,
    \sw_081_module_data_out[2] ,
    \sw_081_module_data_out[1] ,
    \sw_081_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_82 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_082_module_data_in[7] ,
    \sw_082_module_data_in[6] ,
    \sw_082_module_data_in[5] ,
    \sw_082_module_data_in[4] ,
    \sw_082_module_data_in[3] ,
    \sw_082_module_data_in[2] ,
    \sw_082_module_data_in[1] ,
    \sw_082_module_data_in[0] }),
    .io_out({\sw_082_module_data_out[7] ,
    \sw_082_module_data_out[6] ,
    \sw_082_module_data_out[5] ,
    \sw_082_module_data_out[4] ,
    \sw_082_module_data_out[3] ,
    \sw_082_module_data_out[2] ,
    \sw_082_module_data_out[1] ,
    \sw_082_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_83 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_083_module_data_in[7] ,
    \sw_083_module_data_in[6] ,
    \sw_083_module_data_in[5] ,
    \sw_083_module_data_in[4] ,
    \sw_083_module_data_in[3] ,
    \sw_083_module_data_in[2] ,
    \sw_083_module_data_in[1] ,
    \sw_083_module_data_in[0] }),
    .io_out({\sw_083_module_data_out[7] ,
    \sw_083_module_data_out[6] ,
    \sw_083_module_data_out[5] ,
    \sw_083_module_data_out[4] ,
    \sw_083_module_data_out[3] ,
    \sw_083_module_data_out[2] ,
    \sw_083_module_data_out[1] ,
    \sw_083_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_84 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_084_module_data_in[7] ,
    \sw_084_module_data_in[6] ,
    \sw_084_module_data_in[5] ,
    \sw_084_module_data_in[4] ,
    \sw_084_module_data_in[3] ,
    \sw_084_module_data_in[2] ,
    \sw_084_module_data_in[1] ,
    \sw_084_module_data_in[0] }),
    .io_out({\sw_084_module_data_out[7] ,
    \sw_084_module_data_out[6] ,
    \sw_084_module_data_out[5] ,
    \sw_084_module_data_out[4] ,
    \sw_084_module_data_out[3] ,
    \sw_084_module_data_out[2] ,
    \sw_084_module_data_out[1] ,
    \sw_084_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_85 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_085_module_data_in[7] ,
    \sw_085_module_data_in[6] ,
    \sw_085_module_data_in[5] ,
    \sw_085_module_data_in[4] ,
    \sw_085_module_data_in[3] ,
    \sw_085_module_data_in[2] ,
    \sw_085_module_data_in[1] ,
    \sw_085_module_data_in[0] }),
    .io_out({\sw_085_module_data_out[7] ,
    \sw_085_module_data_out[6] ,
    \sw_085_module_data_out[5] ,
    \sw_085_module_data_out[4] ,
    \sw_085_module_data_out[3] ,
    \sw_085_module_data_out[2] ,
    \sw_085_module_data_out[1] ,
    \sw_085_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_86 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_086_module_data_in[7] ,
    \sw_086_module_data_in[6] ,
    \sw_086_module_data_in[5] ,
    \sw_086_module_data_in[4] ,
    \sw_086_module_data_in[3] ,
    \sw_086_module_data_in[2] ,
    \sw_086_module_data_in[1] ,
    \sw_086_module_data_in[0] }),
    .io_out({\sw_086_module_data_out[7] ,
    \sw_086_module_data_out[6] ,
    \sw_086_module_data_out[5] ,
    \sw_086_module_data_out[4] ,
    \sw_086_module_data_out[3] ,
    \sw_086_module_data_out[2] ,
    \sw_086_module_data_out[1] ,
    \sw_086_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_87 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_087_module_data_in[7] ,
    \sw_087_module_data_in[6] ,
    \sw_087_module_data_in[5] ,
    \sw_087_module_data_in[4] ,
    \sw_087_module_data_in[3] ,
    \sw_087_module_data_in[2] ,
    \sw_087_module_data_in[1] ,
    \sw_087_module_data_in[0] }),
    .io_out({\sw_087_module_data_out[7] ,
    \sw_087_module_data_out[6] ,
    \sw_087_module_data_out[5] ,
    \sw_087_module_data_out[4] ,
    \sw_087_module_data_out[3] ,
    \sw_087_module_data_out[2] ,
    \sw_087_module_data_out[1] ,
    \sw_087_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_88 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_088_module_data_in[7] ,
    \sw_088_module_data_in[6] ,
    \sw_088_module_data_in[5] ,
    \sw_088_module_data_in[4] ,
    \sw_088_module_data_in[3] ,
    \sw_088_module_data_in[2] ,
    \sw_088_module_data_in[1] ,
    \sw_088_module_data_in[0] }),
    .io_out({\sw_088_module_data_out[7] ,
    \sw_088_module_data_out[6] ,
    \sw_088_module_data_out[5] ,
    \sw_088_module_data_out[4] ,
    \sw_088_module_data_out[3] ,
    \sw_088_module_data_out[2] ,
    \sw_088_module_data_out[1] ,
    \sw_088_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_89 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_089_module_data_in[7] ,
    \sw_089_module_data_in[6] ,
    \sw_089_module_data_in[5] ,
    \sw_089_module_data_in[4] ,
    \sw_089_module_data_in[3] ,
    \sw_089_module_data_in[2] ,
    \sw_089_module_data_in[1] ,
    \sw_089_module_data_in[0] }),
    .io_out({\sw_089_module_data_out[7] ,
    \sw_089_module_data_out[6] ,
    \sw_089_module_data_out[5] ,
    \sw_089_module_data_out[4] ,
    \sw_089_module_data_out[3] ,
    \sw_089_module_data_out[2] ,
    \sw_089_module_data_out[1] ,
    \sw_089_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_90 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_090_module_data_in[7] ,
    \sw_090_module_data_in[6] ,
    \sw_090_module_data_in[5] ,
    \sw_090_module_data_in[4] ,
    \sw_090_module_data_in[3] ,
    \sw_090_module_data_in[2] ,
    \sw_090_module_data_in[1] ,
    \sw_090_module_data_in[0] }),
    .io_out({\sw_090_module_data_out[7] ,
    \sw_090_module_data_out[6] ,
    \sw_090_module_data_out[5] ,
    \sw_090_module_data_out[4] ,
    \sw_090_module_data_out[3] ,
    \sw_090_module_data_out[2] ,
    \sw_090_module_data_out[1] ,
    \sw_090_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_91 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_091_module_data_in[7] ,
    \sw_091_module_data_in[6] ,
    \sw_091_module_data_in[5] ,
    \sw_091_module_data_in[4] ,
    \sw_091_module_data_in[3] ,
    \sw_091_module_data_in[2] ,
    \sw_091_module_data_in[1] ,
    \sw_091_module_data_in[0] }),
    .io_out({\sw_091_module_data_out[7] ,
    \sw_091_module_data_out[6] ,
    \sw_091_module_data_out[5] ,
    \sw_091_module_data_out[4] ,
    \sw_091_module_data_out[3] ,
    \sw_091_module_data_out[2] ,
    \sw_091_module_data_out[1] ,
    \sw_091_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_92 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_092_module_data_in[7] ,
    \sw_092_module_data_in[6] ,
    \sw_092_module_data_in[5] ,
    \sw_092_module_data_in[4] ,
    \sw_092_module_data_in[3] ,
    \sw_092_module_data_in[2] ,
    \sw_092_module_data_in[1] ,
    \sw_092_module_data_in[0] }),
    .io_out({\sw_092_module_data_out[7] ,
    \sw_092_module_data_out[6] ,
    \sw_092_module_data_out[5] ,
    \sw_092_module_data_out[4] ,
    \sw_092_module_data_out[3] ,
    \sw_092_module_data_out[2] ,
    \sw_092_module_data_out[1] ,
    \sw_092_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_93 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_093_module_data_in[7] ,
    \sw_093_module_data_in[6] ,
    \sw_093_module_data_in[5] ,
    \sw_093_module_data_in[4] ,
    \sw_093_module_data_in[3] ,
    \sw_093_module_data_in[2] ,
    \sw_093_module_data_in[1] ,
    \sw_093_module_data_in[0] }),
    .io_out({\sw_093_module_data_out[7] ,
    \sw_093_module_data_out[6] ,
    \sw_093_module_data_out[5] ,
    \sw_093_module_data_out[4] ,
    \sw_093_module_data_out[3] ,
    \sw_093_module_data_out[2] ,
    \sw_093_module_data_out[1] ,
    \sw_093_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_94 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_094_module_data_in[7] ,
    \sw_094_module_data_in[6] ,
    \sw_094_module_data_in[5] ,
    \sw_094_module_data_in[4] ,
    \sw_094_module_data_in[3] ,
    \sw_094_module_data_in[2] ,
    \sw_094_module_data_in[1] ,
    \sw_094_module_data_in[0] }),
    .io_out({\sw_094_module_data_out[7] ,
    \sw_094_module_data_out[6] ,
    \sw_094_module_data_out[5] ,
    \sw_094_module_data_out[4] ,
    \sw_094_module_data_out[3] ,
    \sw_094_module_data_out[2] ,
    \sw_094_module_data_out[1] ,
    \sw_094_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_95 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_095_module_data_in[7] ,
    \sw_095_module_data_in[6] ,
    \sw_095_module_data_in[5] ,
    \sw_095_module_data_in[4] ,
    \sw_095_module_data_in[3] ,
    \sw_095_module_data_in[2] ,
    \sw_095_module_data_in[1] ,
    \sw_095_module_data_in[0] }),
    .io_out({\sw_095_module_data_out[7] ,
    \sw_095_module_data_out[6] ,
    \sw_095_module_data_out[5] ,
    \sw_095_module_data_out[4] ,
    \sw_095_module_data_out[3] ,
    \sw_095_module_data_out[2] ,
    \sw_095_module_data_out[1] ,
    \sw_095_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_96 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_096_module_data_in[7] ,
    \sw_096_module_data_in[6] ,
    \sw_096_module_data_in[5] ,
    \sw_096_module_data_in[4] ,
    \sw_096_module_data_in[3] ,
    \sw_096_module_data_in[2] ,
    \sw_096_module_data_in[1] ,
    \sw_096_module_data_in[0] }),
    .io_out({\sw_096_module_data_out[7] ,
    \sw_096_module_data_out[6] ,
    \sw_096_module_data_out[5] ,
    \sw_096_module_data_out[4] ,
    \sw_096_module_data_out[3] ,
    \sw_096_module_data_out[2] ,
    \sw_096_module_data_out[1] ,
    \sw_096_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_97 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_097_module_data_in[7] ,
    \sw_097_module_data_in[6] ,
    \sw_097_module_data_in[5] ,
    \sw_097_module_data_in[4] ,
    \sw_097_module_data_in[3] ,
    \sw_097_module_data_in[2] ,
    \sw_097_module_data_in[1] ,
    \sw_097_module_data_in[0] }),
    .io_out({\sw_097_module_data_out[7] ,
    \sw_097_module_data_out[6] ,
    \sw_097_module_data_out[5] ,
    \sw_097_module_data_out[4] ,
    \sw_097_module_data_out[3] ,
    \sw_097_module_data_out[2] ,
    \sw_097_module_data_out[1] ,
    \sw_097_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_98 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_098_module_data_in[7] ,
    \sw_098_module_data_in[6] ,
    \sw_098_module_data_in[5] ,
    \sw_098_module_data_in[4] ,
    \sw_098_module_data_in[3] ,
    \sw_098_module_data_in[2] ,
    \sw_098_module_data_in[1] ,
    \sw_098_module_data_in[0] }),
    .io_out({\sw_098_module_data_out[7] ,
    \sw_098_module_data_out[6] ,
    \sw_098_module_data_out[5] ,
    \sw_098_module_data_out[4] ,
    \sw_098_module_data_out[3] ,
    \sw_098_module_data_out[2] ,
    \sw_098_module_data_out[1] ,
    \sw_098_module_data_out[0] }));
 user_module_339501025136214612 user_module_339501025136214612_99 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_099_module_data_in[7] ,
    \sw_099_module_data_in[6] ,
    \sw_099_module_data_in[5] ,
    \sw_099_module_data_in[4] ,
    \sw_099_module_data_in[3] ,
    \sw_099_module_data_in[2] ,
    \sw_099_module_data_in[1] ,
    \sw_099_module_data_in[0] }),
    .io_out({\sw_099_module_data_out[7] ,
    \sw_099_module_data_out[6] ,
    \sw_099_module_data_out[5] ,
    \sw_099_module_data_out[4] ,
    \sw_099_module_data_out[3] ,
    \sw_099_module_data_out[2] ,
    \sw_099_module_data_out[1] ,
    \sw_099_module_data_out[0] }));
 user_module_342981109408072274 user_module_342981109408072274_22 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_022_module_data_in[7] ,
    \sw_022_module_data_in[6] ,
    \sw_022_module_data_in[5] ,
    \sw_022_module_data_in[4] ,
    \sw_022_module_data_in[3] ,
    \sw_022_module_data_in[2] ,
    \sw_022_module_data_in[1] ,
    \sw_022_module_data_in[0] }),
    .io_out({\sw_022_module_data_out[7] ,
    \sw_022_module_data_out[6] ,
    \sw_022_module_data_out[5] ,
    \sw_022_module_data_out[4] ,
    \sw_022_module_data_out[3] ,
    \sw_022_module_data_out[2] ,
    \sw_022_module_data_out[1] ,
    \sw_022_module_data_out[0] }));
 user_module_346553315158393428 user_module_346553315158393428_16 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_016_module_data_in[7] ,
    \sw_016_module_data_in[6] ,
    \sw_016_module_data_in[5] ,
    \sw_016_module_data_in[4] ,
    \sw_016_module_data_in[3] ,
    \sw_016_module_data_in[2] ,
    \sw_016_module_data_in[1] ,
    \sw_016_module_data_in[0] }),
    .io_out({\sw_016_module_data_out[7] ,
    \sw_016_module_data_out[6] ,
    \sw_016_module_data_out[5] ,
    \sw_016_module_data_out[4] ,
    \sw_016_module_data_out[3] ,
    \sw_016_module_data_out[2] ,
    \sw_016_module_data_out[1] ,
    \sw_016_module_data_out[0] }));
 user_module_346916357828248146 user_module_346916357828248146_18 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_018_module_data_in[7] ,
    \sw_018_module_data_in[6] ,
    \sw_018_module_data_in[5] ,
    \sw_018_module_data_in[4] ,
    \sw_018_module_data_in[3] ,
    \sw_018_module_data_in[2] ,
    \sw_018_module_data_in[1] ,
    \sw_018_module_data_in[0] }),
    .io_out({\sw_018_module_data_out[7] ,
    \sw_018_module_data_out[6] ,
    \sw_018_module_data_out[5] ,
    \sw_018_module_data_out[4] ,
    \sw_018_module_data_out[3] ,
    \sw_018_module_data_out[2] ,
    \sw_018_module_data_out[1] ,
    \sw_018_module_data_out[0] }));
 user_module_347592305412145748 user_module_347592305412145748_13 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_013_module_data_in[7] ,
    \sw_013_module_data_in[6] ,
    \sw_013_module_data_in[5] ,
    \sw_013_module_data_in[4] ,
    \sw_013_module_data_in[3] ,
    \sw_013_module_data_in[2] ,
    \sw_013_module_data_in[1] ,
    \sw_013_module_data_in[0] }),
    .io_out({\sw_013_module_data_out[7] ,
    \sw_013_module_data_out[6] ,
    \sw_013_module_data_out[5] ,
    \sw_013_module_data_out[4] ,
    \sw_013_module_data_out[3] ,
    \sw_013_module_data_out[2] ,
    \sw_013_module_data_out[1] ,
    \sw_013_module_data_out[0] }));
 user_module_347594509754827347 user_module_347594509754827347_19 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_019_module_data_in[7] ,
    \sw_019_module_data_in[6] ,
    \sw_019_module_data_in[5] ,
    \sw_019_module_data_in[4] ,
    \sw_019_module_data_in[3] ,
    \sw_019_module_data_in[2] ,
    \sw_019_module_data_in[1] ,
    \sw_019_module_data_in[0] }),
    .io_out({\sw_019_module_data_out[7] ,
    \sw_019_module_data_out[6] ,
    \sw_019_module_data_out[5] ,
    \sw_019_module_data_out[4] ,
    \sw_019_module_data_out[3] ,
    \sw_019_module_data_out[2] ,
    \sw_019_module_data_out[1] ,
    \sw_019_module_data_out[0] }));
 user_module_347688030570545747 user_module_347688030570545747_21 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_021_module_data_in[7] ,
    \sw_021_module_data_in[6] ,
    \sw_021_module_data_in[5] ,
    \sw_021_module_data_in[4] ,
    \sw_021_module_data_in[3] ,
    \sw_021_module_data_in[2] ,
    \sw_021_module_data_in[1] ,
    \sw_021_module_data_in[0] }),
    .io_out({\sw_021_module_data_out[7] ,
    \sw_021_module_data_out[6] ,
    \sw_021_module_data_out[5] ,
    \sw_021_module_data_out[4] ,
    \sw_021_module_data_out[3] ,
    \sw_021_module_data_out[2] ,
    \sw_021_module_data_out[1] ,
    \sw_021_module_data_out[0] }));
 user_module_347690870424732244 user_module_347690870424732244_12 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_012_module_data_in[7] ,
    \sw_012_module_data_in[6] ,
    \sw_012_module_data_in[5] ,
    \sw_012_module_data_in[4] ,
    \sw_012_module_data_in[3] ,
    \sw_012_module_data_in[2] ,
    \sw_012_module_data_in[1] ,
    \sw_012_module_data_in[0] }),
    .io_out({\sw_012_module_data_out[7] ,
    \sw_012_module_data_out[6] ,
    \sw_012_module_data_out[5] ,
    \sw_012_module_data_out[4] ,
    \sw_012_module_data_out[3] ,
    \sw_012_module_data_out[2] ,
    \sw_012_module_data_out[1] ,
    \sw_012_module_data_out[0] }));
 user_module_347787021138264660 user_module_347787021138264660_10 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_010_module_data_in[7] ,
    \sw_010_module_data_in[6] ,
    \sw_010_module_data_in[5] ,
    \sw_010_module_data_in[4] ,
    \sw_010_module_data_in[3] ,
    \sw_010_module_data_in[2] ,
    \sw_010_module_data_in[1] ,
    \sw_010_module_data_in[0] }),
    .io_out({\sw_010_module_data_out[7] ,
    \sw_010_module_data_out[6] ,
    \sw_010_module_data_out[5] ,
    \sw_010_module_data_out[4] ,
    \sw_010_module_data_out[3] ,
    \sw_010_module_data_out[2] ,
    \sw_010_module_data_out[1] ,
    \sw_010_module_data_out[0] }));
 user_module_347894637149553236 user_module_347894637149553236_17 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_017_module_data_in[7] ,
    \sw_017_module_data_in[6] ,
    \sw_017_module_data_in[5] ,
    \sw_017_module_data_in[4] ,
    \sw_017_module_data_in[3] ,
    \sw_017_module_data_in[2] ,
    \sw_017_module_data_in[1] ,
    \sw_017_module_data_in[0] }),
    .io_out({\sw_017_module_data_out[7] ,
    \sw_017_module_data_out[6] ,
    \sw_017_module_data_out[5] ,
    \sw_017_module_data_out[4] ,
    \sw_017_module_data_out[3] ,
    \sw_017_module_data_out[2] ,
    \sw_017_module_data_out[1] ,
    \sw_017_module_data_out[0] }));
 user_module_348121131386929746 user_module_348121131386929746_28 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_028_module_data_in[7] ,
    \sw_028_module_data_in[6] ,
    \sw_028_module_data_in[5] ,
    \sw_028_module_data_in[4] ,
    \sw_028_module_data_in[3] ,
    \sw_028_module_data_in[2] ,
    \sw_028_module_data_in[1] ,
    \sw_028_module_data_in[0] }),
    .io_out({\sw_028_module_data_out[7] ,
    \sw_028_module_data_out[6] ,
    \sw_028_module_data_out[5] ,
    \sw_028_module_data_out[4] ,
    \sw_028_module_data_out[3] ,
    \sw_028_module_data_out[2] ,
    \sw_028_module_data_out[1] ,
    \sw_028_module_data_out[0] }));
 user_module_348195845106041428 user_module_348195845106041428_27 (.vccd1(vccd1),
    .vssd1(vssd1),
    .io_in({\sw_027_module_data_in[7] ,
    \sw_027_module_data_in[6] ,
    \sw_027_module_data_in[5] ,
    \sw_027_module_data_in[4] ,
    \sw_027_module_data_in[3] ,
    \sw_027_module_data_in[2] ,
    \sw_027_module_data_in[1] ,
    \sw_027_module_data_in[0] }),
    .io_out({\sw_027_module_data_out[7] ,
    \sw_027_module_data_out[6] ,
    \sw_027_module_data_out[5] ,
    \sw_027_module_data_out[4] ,
    \sw_027_module_data_out[3] ,
    \sw_027_module_data_out[2] ,
    \sw_027_module_data_out[1] ,
    \sw_027_module_data_out[0] }));
endmodule
