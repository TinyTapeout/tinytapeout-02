/* Automatically generated from https://wokwi.com/projects/347594509754827347 */

`default_nettype none

module user_module_347594509754827347(
  input [7:0] io_in,
  output [7:0] io_out
);
  wire net1 = io_in[0];
  wire net2 = io_in[1];
  wire net3 = io_in[2];
  wire net4 = io_in[4];
  wire net5 = io_in[5];
  wire net6 = io_in[6];
  wire net7 = io_in[7];
  wire net8;
  wire net9;
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16 = 1'b0;
  wire net17 = 1'b1;
  wire net18 = 1'b1;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37 = 1'b0;
  wire net38 = 1'b0;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45 = 1'b0;
  wire net46 = 1'b0;
  wire net47;
  wire net48;
  wire net49;
  wire net50 = 1'b0;
  wire net51;
  wire net52 = 1'b0;
  wire net53;
  wire net54;
  wire net55;
  wire net56 = 1'b0;
  wire net57;
  wire net58 = 1'b0;
  wire net59;
  wire net60;
  wire net61;
  wire net62 = 1'b0;
  wire net63;
  wire net64 = 1'b0;
  wire net65;
  wire net66;
  wire net67;
  wire net68 = 1'b0;
  wire net69;
  wire net70 = 1'b0;
  wire net71;
  wire net72;
  wire net73;
  wire net74 = 1'b0;
  wire net75;
  wire net76 = 1'b0;
  wire net77;
  wire net78;
  wire net79;
  wire net80 = 1'b0;
  wire net81;
  wire net82 = 1'b0;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90 = 1'b0;
  wire net91 = 1'b0;
  wire net92;
  wire net93;
  wire net94 = 1'b0;
  wire net95;
  wire net96 = 1'b0;
  wire net97;
  wire net98;
  wire net99 = 1'b1;
  wire net100;
  wire net101;
  wire net102 = 1'b1;
  wire net103;
  wire net104;
  wire net105;
  wire net106 = 1'b0;
  wire net107 = 1'b0;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125 = 1'b0;
  wire net126;
  wire net127;
  wire net128 = 1'b0;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150 = 1'b0;
  wire net151;
  wire net152;
  wire net153 = 1'b0;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174 = 1'b0;
  wire net175;
  wire net176;
  wire net177 = 1'b0;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199 = 1'b0;
  wire net200;
  wire net201;
  wire net202 = 1'b0;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224 = 1'b0;
  wire net225;
  wire net226;
  wire net227 = 1'b0;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249 = 1'b0;
  wire net250;
  wire net251;
  wire net252 = 1'b0;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273 = 1'b0;
  wire net274;
  wire net275;
  wire net276 = 1'b0;
  wire net277;
  wire net278;
  wire net279;
  wire net280 = 1'b0;
  wire net281 = 1'b0;
  wire net282;
  wire net283 = 1'b0;
  wire net284 = 1'b1;
  wire net285;
  wire net286 = 1'b0;
  wire net287 = 1'b1;
  wire net288;
  wire net289 = 1'b0;
  wire net290 = 1'b1;
  wire net291;
  wire net292 = 1'b0;
  wire net293 = 1'b1;
  wire net294;
  wire net295 = 1'b0;
  wire net296 = 1'b1;
  wire net297;
  wire net298 = 1'b0;
  wire net299 = 1'b0;
  wire net300;
  wire net301;
  wire net302 = 1'b0;
  wire net303 = 1'b0;
  wire net304 = 1'b1;
  wire net305 = 1'b1;
  wire net306;
  wire net307 = 1'b1;
  wire net308 = 1'b0;
  wire net309;
  wire net310 = 1'b1;
  wire net311 = 1'b0;
  wire net312;
  wire net313 = 1'b1;
  wire net314 = 1'b0;
  wire net315;
  wire net316 = 1'b1;
  wire net317 = 1'b0;
  wire net318;
  wire net319 = 1'b1;
  wire net320 = 1'b0;
  wire net321;
  wire net322 = 1'b1;
  wire net323 = 1'b0;
  wire net324;
  wire net325 = 1'b0;
  wire net326 = 1'b0;
  wire net327;
  wire net328 = 1'b0;
  wire net329 = 1'b0;
  wire net330;
  wire net331 = 1'b0;
  wire net332 = 1'b0;
  wire net333;
  wire net334 = 1'b0;
  wire net335 = 1'b1;
  wire net336;
  wire net337 = 1'b0;
  wire net338 = 1'b1;
  wire net339;
  wire net340 = 1'b0;
  wire net341 = 1'b1;
  wire net342;
  wire net343 = 1'b0;
  wire net344 = 1'b0;
  wire net345;
  wire net346;
  wire net347 = 1'b0;
  wire net348 = 1'b0;
  wire net349 = 1'b1;
  wire net350 = 1'b1;
  wire net351;
  wire net352 = 1'b0;
  wire net353 = 1'b0;
  wire net354;
  wire net355 = 1'b0;
  wire net356 = 1'b1;
  wire net357;
  wire net358 = 1'b0;
  wire net359 = 1'b0;
  wire net360;
  wire net361 = 1'b0;
  wire net362 = 1'b0;
  wire net363;
  wire net364 = 1'b0;
  wire net365 = 1'b0;
  wire net366;
  wire net367 = 1'b0;
  wire net368 = 1'b1;
  wire net369;
  wire net370 = 1'b0;
  wire net371 = 1'b0;
  wire net372;
  wire net373;
  wire net374 = 1'b0;
  wire net375 = 1'b0;
  wire net376 = 1'b1;
  wire net377 = 1'b0;
  wire net378;
  wire net379 = 1'b0;
  wire net380 = 1'b0;
  wire net381;
  wire net382 = 1'b0;
  wire net383 = 1'b1;
  wire net384;
  wire net385 = 1'b0;
  wire net386 = 1'b1;
  wire net387;
  wire net388 = 1'b0;
  wire net389 = 1'b0;
  wire net390;
  wire net391 = 1'b0;
  wire net392 = 1'b1;
  wire net393;
  wire net394 = 1'b0;
  wire net395 = 1'b1;
  wire net396;
  wire net397 = 1'b0;
  wire net398 = 1'b0;
  wire net399;
  wire net400;
  wire net401 = 1'b0;
  wire net402 = 1'b0;
  wire net403 = 1'b1;
  wire net404 = 1'b1;
  wire net405;
  wire net406 = 1'b0;
  wire net407 = 1'b1;
  wire net408;
  wire net409 = 1'b0;
  wire net410 = 1'b0;
  wire net411;
  wire net412 = 1'b0;
  wire net413 = 1'b1;
  wire net414;
  wire net415 = 1'b0;
  wire net416 = 1'b1;
  wire net417;
  wire net418 = 1'b0;
  wire net419 = 1'b1;
  wire net420;
  wire net421 = 1'b0;
  wire net422 = 1'b1;
  wire net423;
  wire net424 = 1'b0;
  wire net425 = 1'b1;
  wire net426;
  wire net427;
  wire net428 = 1'b0;
  wire net429 = 1'b0;
  wire net430 = 1'b1;
  wire net431 = 1'b1;
  wire net432;
  wire net433 = 1'b0;
  wire net434 = 1'b1;
  wire net435;
  wire net436 = 1'b0;
  wire net437 = 1'b1;
  wire net438;
  wire net439 = 1'b0;
  wire net440 = 1'b1;
  wire net441;
  wire net442 = 1'b0;
  wire net443 = 1'b1;
  wire net444;
  wire net445 = 1'b0;
  wire net446 = 1'b0;
  wire net447;
  wire net448 = 1'b0;
  wire net449 = 1'b0;
  wire net450;
  wire net451 = 1'b0;
  wire net452 = 1'b1;
  wire net453;
  wire net454;
  wire net455 = 1'b0;
  wire net456 = 1'b0;
  wire net457 = 1'b1;
  wire net458 = 1'b1;
  wire net459;
  wire net460 = 1'b0;
  wire net461 = 1'b0;
  wire net462;
  wire net463 = 1'b0;
  wire net464 = 1'b1;
  wire net465;
  wire net466 = 1'b0;
  wire net467 = 1'b1;
  wire net468;
  wire net469 = 1'b0;
  wire net470 = 1'b0;
  wire net471;
  wire net472 = 1'b0;
  wire net473 = 1'b1;
  wire net474;
  wire net475 = 1'b0;
  wire net476 = 1'b1;
  wire net477;
  wire net478 = 1'b0;
  wire net479 = 1'b1;
  wire net480;
  wire net481;
  wire net482 = 1'b0;
  wire net483 = 1'b0;
  wire net484 = 1'b1;
  wire net485 = 1'b1;
  wire net486 = 1'b0;

  assign io_out[0] = net8;
  assign io_out[1] = net9;
  assign io_out[2] = net10;
  assign io_out[3] = net11;
  assign io_out[4] = net12;
  assign io_out[5] = net13;
  assign io_out[6] = net14;
  assign io_out[7] = net15;

  and_cell gate1 (

  );
  or_cell gate2 (

  );
  xor_cell gate3 (

  );
  nand_cell gate4 (

  );
  not_cell gate5 (

  );
  buffer_cell gate6 (

  );
  mux_cell mux1 (

  );
  dff_cell flipflop1 (

  );
  mux_cell mux2 (
    .a (net19),
    .b (net20),
    .sel (net21),
    .out (net22)
  );
  mux_cell mux7 (
    .a (net23),
    .b (net24),
    .sel (net25),
    .out (net20)
  );
  mux_cell mux12 (
    .a (net26),
    .b (net27),
    .sel (net25),
    .out (net19)
  );
  mux_cell mux5 (
    .a (net28),
    .b (net29),
    .sel (net30),
    .out (net27)
  );
  mux_cell mux6 (
    .a (net31),
    .b (net32),
    .sel (net30),
    .out (net26)
  );
  dff_cell flipflop2 (
    .d (net33),
    .clk (net34),
    .q (net31)
  );
  dff_cell flipflop10 (
    .d (net35),
    .clk (net36),
    .q (net32)
  );
  mux_cell mux18 (
    .a (net39),
    .b (net40),
    .sel (net30),
    .out (net24)
  );
  mux_cell mux19 (
    .a (net41),
    .b (net42),
    .sel (net30),
    .out (net23)
  );
  buffer_cell gate7 (
    .in (net1),
    .out (net34)
  );
  not_cell gate8 (
    .in (net3),
    .out (net43)
  );
  buffer_cell gate9 (
    .in (net1),
    .out (net36)
  );
  not_cell gate10 (
    .in (net3),
    .out (net44)
  );
  buffer_cell gate11 (
    .in (net7),
    .out (net30)
  );
  buffer_cell gate12 (
    .in (net6),
    .out (net25)
  );
  buffer_cell gate13 (
    .in (net5),
    .out (net21)
  );
  mux_cell mux3 (
    .a (net45),
    .b (net2),
    .sel (net43),
    .out (net33)
  );
  mux_cell mux4 (
    .a (net46),
    .b (net47),
    .sel (net44),
    .out (net35)
  );
  dff_cell flipflop8 (
    .d (net48),
    .clk (net49),
    .q (net28)
  );
  buffer_cell gate14 (
    .in (net1),
    .out (net49)
  );
  not_cell gate15 (
    .in (net3),
    .out (net51)
  );
  mux_cell mux11 (
    .a (net52),
    .b (net53),
    .sel (net51),
    .out (net48)
  );
  dff_cell flipflop3 (
    .d (net54),
    .clk (net55),
    .q (net29)
  );
  buffer_cell gate16 (
    .in (net1),
    .out (net55)
  );
  not_cell gate17 (
    .in (net3),
    .out (net57)
  );
  mux_cell mux16 (
    .a (net58),
    .b (net59),
    .sel (net57),
    .out (net54)
  );
  dff_cell flipflop4 (
    .d (net60),
    .clk (net61),
    .q (net41)
  );
  buffer_cell gate18 (
    .in (net1),
    .out (net61)
  );
  not_cell gate19 (
    .in (net3),
    .out (net63)
  );
  mux_cell mux17 (
    .a (net64),
    .b (net65),
    .sel (net63),
    .out (net60)
  );
  dff_cell flipflop5 (
    .d (net66),
    .clk (net67),
    .q (net42)
  );
  buffer_cell gate20 (
    .in (net1),
    .out (net67)
  );
  not_cell gate21 (
    .in (net3),
    .out (net69)
  );
  mux_cell mux24 (
    .a (net70),
    .b (net71),
    .sel (net69),
    .out (net66)
  );
  dff_cell flipflop6 (
    .d (net72),
    .clk (net73),
    .q (net39)
  );
  buffer_cell gate22 (
    .in (net1),
    .out (net73)
  );
  not_cell gate23 (
    .in (net3),
    .out (net75)
  );
  mux_cell mux25 (
    .a (net76),
    .b (net77),
    .sel (net75),
    .out (net72)
  );
  dff_cell flipflop7 (
    .d (net78),
    .clk (net79),
    .q (net40)
  );
  buffer_cell gate24 (
    .in (net1),
    .out (net79)
  );
  not_cell gate25 (
    .in (net3),
    .out (net81)
  );
  mux_cell mux30 (
    .a (net82),
    .b (net83),
    .sel (net81),
    .out (net78)
  );
  dff_cell flipflop9 (
    .d (net84),
    .clk (net85),
    .q (net86)
  );
  dff_cell flipflop11 (
    .d (net87),
    .clk (net88),
    .q (net89)
  );
  buffer_cell gate26 (
    .in (net1),
    .out (net85)
  );
  not_cell gate27 (
    .in (net3),
    .out (net92)
  );
  buffer_cell gate28 (
    .in (net1),
    .out (net88)
  );
  not_cell gate29 (
    .in (net3),
    .out (net93)
  );
  mux_cell mux33 (
    .a (net94),
    .b (net95),
    .sel (net92),
    .out (net84)
  );
  mux_cell mux34 (
    .a (net96),
    .b (net97),
    .sel (net93),
    .out (net87)
  );
  mux_cell mux43 (
    .a (net98),
    .b (net99),
    .sel (net21),
    .out (net100)
  );
  mux_cell mux45 (
    .a (net101),
    .b (net102),
    .sel (net25),
    .out (net98)
  );
  mux_cell mux47 (
    .a (net86),
    .b (net89),
    .sel (net30),
    .out (net101)
  );
  mux_cell mux50 (
    .a (net22),
    .b (net100),
    .sel (net103),
    .out (net15)
  );
  buffer_cell gate42 (
    .in (net4),
    .out (net103)
  );
  dff_cell flipflop18 (
    .d (net104),
    .clk (net34),
    .q (net105)
  );
  mux_cell mux8 (
    .a (net107),
    .b (net31),
    .sel (net43),
    .out (net104)
  );
  mux_cell mux9 (
    .a (net108),
    .b (net109),
    .sel (net21),
    .out (net110)
  );
  mux_cell mux10 (
    .a (net111),
    .b (net112),
    .sel (net113),
    .out (net109)
  );
  mux_cell mux13 (
    .a (net114),
    .b (net115),
    .sel (net113),
    .out (net108)
  );
  mux_cell mux14 (
    .a (net116),
    .b (net117),
    .sel (net118),
    .out (net115)
  );
  mux_cell mux15 (
    .a (net105),
    .b (net119),
    .sel (net118),
    .out (net114)
  );
  mux_cell mux20 (
    .a (net120),
    .b (net121),
    .sel (net118),
    .out (net112)
  );
  mux_cell mux21 (
    .a (net122),
    .b (net123),
    .sel (net118),
    .out (net111)
  );
  mux_cell mux22 (
    .a (net124),
    .b (net125),
    .sel (net21),
    .out (net126)
  );
  mux_cell mux26 (
    .a (net127),
    .b (net128),
    .sel (net113),
    .out (net124)
  );
  mux_cell mux28 (
    .a (net129),
    .b (net130),
    .sel (net118),
    .out (net127)
  );
  mux_cell mux32 (
    .a (net110),
    .b (net126),
    .sel (net103),
    .out (net14)
  );
  mux_cell mux42 (
    .a (net131),
    .b (net132),
    .sel (net133),
    .out (net134)
  );
  mux_cell mux51 (
    .a (net135),
    .b (net136),
    .sel (net137),
    .out (net132)
  );
  mux_cell mux52 (
    .a (net138),
    .b (net139),
    .sel (net137),
    .out (net131)
  );
  mux_cell mux53 (
    .a (net140),
    .b (net141),
    .sel (net142),
    .out (net139)
  );
  mux_cell mux54 (
    .a (net143),
    .b (net144),
    .sel (net142),
    .out (net138)
  );
  mux_cell mux55 (
    .a (net145),
    .b (net146),
    .sel (net142),
    .out (net136)
  );
  mux_cell mux56 (
    .a (net147),
    .b (net148),
    .sel (net142),
    .out (net135)
  );
  mux_cell mux57 (
    .a (net149),
    .b (net150),
    .sel (net133),
    .out (net151)
  );
  mux_cell mux59 (
    .a (net152),
    .b (net153),
    .sel (net137),
    .out (net149)
  );
  mux_cell mux61 (
    .a (net154),
    .b (net155),
    .sel (net142),
    .out (net152)
  );
  mux_cell mux64 (
    .a (net134),
    .b (net151),
    .sel (net103),
    .out (net13)
  );
  mux_cell mux66 (
    .a (net156),
    .b (net157),
    .sel (net133),
    .out (net158)
  );
  mux_cell mux67 (
    .a (net159),
    .b (net160),
    .sel (net161),
    .out (net157)
  );
  mux_cell mux68 (
    .a (net162),
    .b (net163),
    .sel (net161),
    .out (net156)
  );
  mux_cell mux69 (
    .a (net164),
    .b (net165),
    .sel (net166),
    .out (net163)
  );
  mux_cell mux70 (
    .a (net167),
    .b (net168),
    .sel (net166),
    .out (net162)
  );
  mux_cell mux71 (
    .a (net169),
    .b (net170),
    .sel (net166),
    .out (net160)
  );
  mux_cell mux72 (
    .a (net171),
    .b (net172),
    .sel (net166),
    .out (net159)
  );
  mux_cell mux73 (
    .a (net173),
    .b (net174),
    .sel (net133),
    .out (net175)
  );
  mux_cell mux75 (
    .a (net176),
    .b (net177),
    .sel (net161),
    .out (net173)
  );
  mux_cell mux77 (
    .a (net178),
    .b (net179),
    .sel (net166),
    .out (net176)
  );
  mux_cell mux80 (
    .a (net158),
    .b (net175),
    .sel (net103),
    .out (net12)
  );
  mux_cell mux82 (
    .a (net180),
    .b (net181),
    .sel (net182),
    .out (net183)
  );
  mux_cell mux83 (
    .a (net184),
    .b (net185),
    .sel (net186),
    .out (net181)
  );
  mux_cell mux84 (
    .a (net187),
    .b (net188),
    .sel (net186),
    .out (net180)
  );
  mux_cell mux85 (
    .a (net189),
    .b (net190),
    .sel (net191),
    .out (net188)
  );
  mux_cell mux86 (
    .a (net192),
    .b (net193),
    .sel (net191),
    .out (net187)
  );
  mux_cell mux87 (
    .a (net194),
    .b (net195),
    .sel (net191),
    .out (net185)
  );
  mux_cell mux88 (
    .a (net196),
    .b (net197),
    .sel (net191),
    .out (net184)
  );
  mux_cell mux89 (
    .a (net198),
    .b (net199),
    .sel (net182),
    .out (net200)
  );
  mux_cell mux91 (
    .a (net201),
    .b (net202),
    .sel (net186),
    .out (net198)
  );
  mux_cell mux93 (
    .a (net203),
    .b (net204),
    .sel (net191),
    .out (net201)
  );
  mux_cell mux96 (
    .a (net183),
    .b (net200),
    .sel (net205),
    .out (net11)
  );
  mux_cell mux98 (
    .a (net206),
    .b (net207),
    .sel (net182),
    .out (net208)
  );
  mux_cell mux99 (
    .a (net209),
    .b (net210),
    .sel (net211),
    .out (net207)
  );
  mux_cell mux100 (
    .a (net212),
    .b (net213),
    .sel (net211),
    .out (net206)
  );
  mux_cell mux101 (
    .a (net214),
    .b (net215),
    .sel (net216),
    .out (net213)
  );
  mux_cell mux102 (
    .a (net217),
    .b (net218),
    .sel (net216),
    .out (net212)
  );
  mux_cell mux103 (
    .a (net219),
    .b (net220),
    .sel (net216),
    .out (net210)
  );
  mux_cell mux104 (
    .a (net221),
    .b (net222),
    .sel (net216),
    .out (net209)
  );
  mux_cell mux105 (
    .a (net223),
    .b (net224),
    .sel (net182),
    .out (net225)
  );
  mux_cell mux107 (
    .a (net226),
    .b (net227),
    .sel (net211),
    .out (net223)
  );
  mux_cell mux109 (
    .a (net228),
    .b (net229),
    .sel (net216),
    .out (net226)
  );
  mux_cell mux112 (
    .a (net208),
    .b (net225),
    .sel (net205),
    .out (net10)
  );
  mux_cell mux114 (
    .a (net230),
    .b (net231),
    .sel (net232),
    .out (net233)
  );
  mux_cell mux115 (
    .a (net234),
    .b (net235),
    .sel (net236),
    .out (net231)
  );
  mux_cell mux116 (
    .a (net237),
    .b (net238),
    .sel (net236),
    .out (net230)
  );
  mux_cell mux117 (
    .a (net239),
    .b (net240),
    .sel (net241),
    .out (net238)
  );
  mux_cell mux118 (
    .a (net242),
    .b (net243),
    .sel (net241),
    .out (net237)
  );
  mux_cell mux119 (
    .a (net244),
    .b (net245),
    .sel (net241),
    .out (net235)
  );
  mux_cell mux120 (
    .a (net246),
    .b (net247),
    .sel (net241),
    .out (net234)
  );
  mux_cell mux121 (
    .a (net248),
    .b (net249),
    .sel (net232),
    .out (net250)
  );
  mux_cell mux123 (
    .a (net251),
    .b (net252),
    .sel (net236),
    .out (net248)
  );
  mux_cell mux125 (
    .a (net253),
    .b (net254),
    .sel (net241),
    .out (net251)
  );
  mux_cell mux128 (
    .a (net233),
    .b (net250),
    .sel (net205),
    .out (net9)
  );
  mux_cell mux130 (
    .a (net255),
    .b (net256),
    .sel (net232),
    .out (net257)
  );
  mux_cell mux131 (
    .a (net258),
    .b (net259),
    .sel (net260),
    .out (net256)
  );
  mux_cell mux132 (
    .a (net261),
    .b (net262),
    .sel (net260),
    .out (net255)
  );
  mux_cell mux133 (
    .a (net263),
    .b (net264),
    .sel (net265),
    .out (net262)
  );
  mux_cell mux134 (
    .a (net266),
    .b (net267),
    .sel (net265),
    .out (net261)
  );
  mux_cell mux135 (
    .a (net268),
    .b (net269),
    .sel (net265),
    .out (net259)
  );
  mux_cell mux136 (
    .a (net270),
    .b (net271),
    .sel (net265),
    .out (net258)
  );
  mux_cell mux137 (
    .a (net272),
    .b (net273),
    .sel (net232),
    .out (net274)
  );
  mux_cell mux139 (
    .a (net275),
    .b (net276),
    .sel (net260),
    .out (net272)
  );
  mux_cell mux141 (
    .a (net277),
    .b (net278),
    .sel (net265),
    .out (net275)
  );
  mux_cell mux144 (
    .a (net257),
    .b (net274),
    .sel (net205),
    .out (net8)
  );
  dff_cell flipflop20 (
    .d (net279),
    .clk (net36),
    .q (net119)
  );
  mux_cell mux41 (
    .a (net281),
    .b (net32),
    .sel (net44),
    .out (net279)
  );
  dff_cell flipflop21 (
    .d (net282),
    .clk (net49),
    .q (net116)
  );
  mux_cell mux65 (
    .a (net284),
    .b (net28),
    .sel (net51),
    .out (net282)
  );
  dff_cell flipflop22 (
    .d (net285),
    .clk (net55),
    .q (net117)
  );
  mux_cell mux81 (
    .a (net287),
    .b (net29),
    .sel (net57),
    .out (net285)
  );
  dff_cell flipflop23 (
    .d (net288),
    .clk (net61),
    .q (net122)
  );
  mux_cell mux97 (
    .a (net290),
    .b (net41),
    .sel (net63),
    .out (net288)
  );
  dff_cell flipflop24 (
    .d (net291),
    .clk (net67),
    .q (net123)
  );
  mux_cell mux113 (
    .a (net293),
    .b (net42),
    .sel (net69),
    .out (net291)
  );
  dff_cell flipflop25 (
    .d (net294),
    .clk (net73),
    .q (net120)
  );
  mux_cell mux129 (
    .a (net296),
    .b (net39),
    .sel (net75),
    .out (net294)
  );
  dff_cell flipflop26 (
    .d (net297),
    .clk (net79),
    .q (net121)
  );
  mux_cell mux145 (
    .a (net299),
    .b (net40),
    .sel (net81),
    .out (net297)
  );
  dff_cell flipflop27 (
    .d (net300),
    .clk (net85),
    .q (net129)
  );
  dff_cell flipflop28 (
    .d (net301),
    .clk (net88),
    .q (net130)
  );
  mux_cell mux146 (
    .a (net304),
    .b (net86),
    .sel (net92),
    .out (net300)
  );
  mux_cell mux147 (
    .a (net305),
    .b (net89),
    .sel (net93),
    .out (net301)
  );
  dff_cell flipflop19 (
    .d (net306),
    .clk (net34),
    .q (net143)
  );
  mux_cell mux154 (
    .a (net307),
    .b (net105),
    .sel (net43),
    .out (net306)
  );
  dff_cell flipflop35 (
    .d (net309),
    .clk (net34),
    .q (net167)
  );
  mux_cell mux155 (
    .a (net310),
    .b (net143),
    .sel (net43),
    .out (net309)
  );
  dff_cell flipflop36 (
    .d (net312),
    .clk (net34),
    .q (net192)
  );
  mux_cell mux156 (
    .a (net313),
    .b (net167),
    .sel (net43),
    .out (net312)
  );
  dff_cell flipflop37 (
    .d (net315),
    .clk (net34),
    .q (net217)
  );
  mux_cell mux157 (
    .a (net316),
    .b (net192),
    .sel (net43),
    .out (net315)
  );
  dff_cell flipflop38 (
    .d (net318),
    .clk (net34),
    .q (net242)
  );
  mux_cell mux158 (
    .a (net319),
    .b (net217),
    .sel (net43),
    .out (net318)
  );
  dff_cell flipflop39 (
    .d (net321),
    .clk (net34),
    .q (net266)
  );
  mux_cell mux159 (
    .a (net322),
    .b (net242),
    .sel (net43),
    .out (net321)
  );
  dff_cell flipflop41 (
    .d (net324),
    .clk (net36),
    .q (net144)
  );
  mux_cell mux160 (
    .a (net326),
    .b (net119),
    .sel (net44),
    .out (net324)
  );
  dff_cell flipflop42 (
    .d (net327),
    .clk (net49),
    .q (net140)
  );
  mux_cell mux161 (
    .a (net329),
    .b (net116),
    .sel (net51),
    .out (net327)
  );
  dff_cell flipflop43 (
    .d (net330),
    .clk (net55),
    .q (net141)
  );
  mux_cell mux162 (
    .a (net332),
    .b (net117),
    .sel (net57),
    .out (net330)
  );
  dff_cell flipflop44 (
    .d (net333),
    .clk (net61),
    .q (net147)
  );
  mux_cell mux163 (
    .a (net335),
    .b (net122),
    .sel (net63),
    .out (net333)
  );
  dff_cell flipflop45 (
    .d (net336),
    .clk (net67),
    .q (net148)
  );
  mux_cell mux164 (
    .a (net338),
    .b (net123),
    .sel (net69),
    .out (net336)
  );
  dff_cell flipflop46 (
    .d (net339),
    .clk (net73),
    .q (net145)
  );
  mux_cell mux165 (
    .a (net341),
    .b (net120),
    .sel (net75),
    .out (net339)
  );
  dff_cell flipflop47 (
    .d (net342),
    .clk (net79),
    .q (net146)
  );
  mux_cell mux166 (
    .a (net344),
    .b (net121),
    .sel (net81),
    .out (net342)
  );
  dff_cell flipflop48 (
    .d (net345),
    .clk (net85),
    .q (net154)
  );
  dff_cell flipflop49 (
    .d (net346),
    .clk (net88),
    .q (net155)
  );
  mux_cell mux167 (
    .a (net349),
    .b (net129),
    .sel (net92),
    .out (net345)
  );
  mux_cell mux168 (
    .a (net350),
    .b (net130),
    .sel (net93),
    .out (net346)
  );
  dff_cell flipflop56 (
    .d (net351),
    .clk (net36),
    .q (net168)
  );
  mux_cell mux175 (
    .a (net353),
    .b (net144),
    .sel (net44),
    .out (net351)
  );
  dff_cell flipflop57 (
    .d (net354),
    .clk (net49),
    .q (net164)
  );
  mux_cell mux176 (
    .a (net356),
    .b (net140),
    .sel (net51),
    .out (net354)
  );
  dff_cell flipflop58 (
    .d (net357),
    .clk (net55),
    .q (net165)
  );
  mux_cell mux177 (
    .a (net359),
    .b (net141),
    .sel (net57),
    .out (net357)
  );
  dff_cell flipflop59 (
    .d (net360),
    .clk (net61),
    .q (net171)
  );
  mux_cell mux178 (
    .a (net362),
    .b (net147),
    .sel (net63),
    .out (net360)
  );
  dff_cell flipflop60 (
    .d (net363),
    .clk (net67),
    .q (net172)
  );
  mux_cell mux179 (
    .a (net365),
    .b (net148),
    .sel (net69),
    .out (net363)
  );
  dff_cell flipflop61 (
    .d (net366),
    .clk (net73),
    .q (net169)
  );
  mux_cell mux180 (
    .a (net368),
    .b (net145),
    .sel (net75),
    .out (net366)
  );
  dff_cell flipflop62 (
    .d (net369),
    .clk (net79),
    .q (net170)
  );
  mux_cell mux181 (
    .a (net371),
    .b (net146),
    .sel (net81),
    .out (net369)
  );
  dff_cell flipflop63 (
    .d (net372),
    .clk (net85),
    .q (net178)
  );
  dff_cell flipflop64 (
    .d (net373),
    .clk (net88),
    .q (net179)
  );
  mux_cell mux182 (
    .a (net376),
    .b (net154),
    .sel (net92),
    .out (net372)
  );
  mux_cell mux183 (
    .a (net377),
    .b (net155),
    .sel (net93),
    .out (net373)
  );
  dff_cell flipflop72 (
    .d (net378),
    .clk (net36),
    .q (net193)
  );
  mux_cell mux190 (
    .a (net380),
    .b (net168),
    .sel (net44),
    .out (net378)
  );
  dff_cell flipflop73 (
    .d (net381),
    .clk (net49),
    .q (net189)
  );
  mux_cell mux191 (
    .a (net383),
    .b (net164),
    .sel (net51),
    .out (net381)
  );
  dff_cell flipflop74 (
    .d (net384),
    .clk (net55),
    .q (net190)
  );
  mux_cell mux192 (
    .a (net386),
    .b (net165),
    .sel (net57),
    .out (net384)
  );
  dff_cell flipflop75 (
    .d (net387),
    .clk (net61),
    .q (net196)
  );
  mux_cell mux193 (
    .a (net389),
    .b (net171),
    .sel (net63),
    .out (net387)
  );
  dff_cell flipflop76 (
    .d (net390),
    .clk (net67),
    .q (net197)
  );
  mux_cell mux194 (
    .a (net392),
    .b (net172),
    .sel (net69),
    .out (net390)
  );
  dff_cell flipflop77 (
    .d (net393),
    .clk (net73),
    .q (net194)
  );
  mux_cell mux195 (
    .a (net395),
    .b (net169),
    .sel (net75),
    .out (net393)
  );
  dff_cell flipflop78 (
    .d (net396),
    .clk (net79),
    .q (net195)
  );
  mux_cell mux196 (
    .a (net398),
    .b (net170),
    .sel (net81),
    .out (net396)
  );
  dff_cell flipflop79 (
    .d (net399),
    .clk (net85),
    .q (net203)
  );
  dff_cell flipflop80 (
    .d (net400),
    .clk (net88),
    .q (net204)
  );
  mux_cell mux197 (
    .a (net403),
    .b (net178),
    .sel (net92),
    .out (net399)
  );
  mux_cell mux198 (
    .a (net404),
    .b (net179),
    .sel (net93),
    .out (net400)
  );
  dff_cell flipflop87 (
    .d (net405),
    .clk (net36),
    .q (net218)
  );
  mux_cell mux205 (
    .a (net407),
    .b (net193),
    .sel (net44),
    .out (net405)
  );
  dff_cell flipflop88 (
    .d (net408),
    .clk (net49),
    .q (net214)
  );
  mux_cell mux206 (
    .a (net410),
    .b (net189),
    .sel (net51),
    .out (net408)
  );
  dff_cell flipflop89 (
    .d (net411),
    .clk (net55),
    .q (net215)
  );
  mux_cell mux207 (
    .a (net413),
    .b (net190),
    .sel (net57),
    .out (net411)
  );
  dff_cell flipflop90 (
    .d (net414),
    .clk (net61),
    .q (net221)
  );
  mux_cell mux208 (
    .a (net416),
    .b (net196),
    .sel (net63),
    .out (net414)
  );
  dff_cell flipflop91 (
    .d (net417),
    .clk (net67),
    .q (net222)
  );
  mux_cell mux209 (
    .a (net419),
    .b (net197),
    .sel (net69),
    .out (net417)
  );
  dff_cell flipflop92 (
    .d (net420),
    .clk (net73),
    .q (net219)
  );
  mux_cell mux210 (
    .a (net422),
    .b (net194),
    .sel (net75),
    .out (net420)
  );
  dff_cell flipflop93 (
    .d (net423),
    .clk (net79),
    .q (net220)
  );
  mux_cell mux211 (
    .a (net425),
    .b (net195),
    .sel (net81),
    .out (net423)
  );
  dff_cell flipflop94 (
    .d (net426),
    .clk (net85),
    .q (net228)
  );
  dff_cell flipflop95 (
    .d (net427),
    .clk (net88),
    .q (net229)
  );
  mux_cell mux212 (
    .a (net430),
    .b (net203),
    .sel (net92),
    .out (net426)
  );
  mux_cell mux213 (
    .a (net431),
    .b (net204),
    .sel (net93),
    .out (net427)
  );
  dff_cell flipflop103 (
    .d (net432),
    .clk (net36),
    .q (net243)
  );
  mux_cell mux220 (
    .a (net434),
    .b (net218),
    .sel (net44),
    .out (net432)
  );
  dff_cell flipflop104 (
    .d (net435),
    .clk (net49),
    .q (net239)
  );
  mux_cell mux221 (
    .a (net437),
    .b (net214),
    .sel (net51),
    .out (net435)
  );
  dff_cell flipflop105 (
    .d (net438),
    .clk (net55),
    .q (net240)
  );
  mux_cell mux222 (
    .a (net440),
    .b (net215),
    .sel (net57),
    .out (net438)
  );
  dff_cell flipflop106 (
    .d (net441),
    .clk (net61),
    .q (net246)
  );
  mux_cell mux223 (
    .a (net443),
    .b (net221),
    .sel (net63),
    .out (net441)
  );
  dff_cell flipflop107 (
    .d (net444),
    .clk (net67),
    .q (net247)
  );
  mux_cell mux224 (
    .a (net446),
    .b (net222),
    .sel (net69),
    .out (net444)
  );
  dff_cell flipflop108 (
    .d (net447),
    .clk (net73),
    .q (net244)
  );
  mux_cell mux225 (
    .a (net449),
    .b (net219),
    .sel (net75),
    .out (net447)
  );
  dff_cell flipflop109 (
    .d (net450),
    .clk (net79),
    .q (net245)
  );
  mux_cell mux226 (
    .a (net452),
    .b (net220),
    .sel (net81),
    .out (net450)
  );
  dff_cell flipflop110 (
    .d (net453),
    .clk (net85),
    .q (net253)
  );
  dff_cell flipflop111 (
    .d (net454),
    .clk (net88),
    .q (net254)
  );
  mux_cell mux227 (
    .a (net457),
    .b (net228),
    .sel (net92),
    .out (net453)
  );
  mux_cell mux228 (
    .a (net458),
    .b (net229),
    .sel (net93),
    .out (net454)
  );
  dff_cell flipflop118 (
    .d (net459),
    .clk (net36),
    .q (net267)
  );
  mux_cell mux235 (
    .a (net461),
    .b (net243),
    .sel (net44),
    .out (net459)
  );
  dff_cell flipflop119 (
    .d (net462),
    .clk (net49),
    .q (net263)
  );
  mux_cell mux236 (
    .a (net464),
    .b (net239),
    .sel (net51),
    .out (net462)
  );
  dff_cell flipflop120 (
    .d (net465),
    .clk (net55),
    .q (net264)
  );
  mux_cell mux237 (
    .a (net467),
    .b (net240),
    .sel (net57),
    .out (net465)
  );
  dff_cell flipflop121 (
    .d (net468),
    .clk (net61),
    .q (net270)
  );
  mux_cell mux238 (
    .a (net470),
    .b (net246),
    .sel (net63),
    .out (net468)
  );
  dff_cell flipflop122 (
    .d (net471),
    .clk (net67),
    .q (net271)
  );
  mux_cell mux239 (
    .a (net473),
    .b (net247),
    .sel (net69),
    .out (net471)
  );
  dff_cell flipflop123 (
    .d (net474),
    .clk (net73),
    .q (net268)
  );
  mux_cell mux240 (
    .a (net476),
    .b (net244),
    .sel (net75),
    .out (net474)
  );
  dff_cell flipflop124 (
    .d (net477),
    .clk (net79),
    .q (net269)
  );
  mux_cell mux241 (
    .a (net479),
    .b (net245),
    .sel (net81),
    .out (net477)
  );
  dff_cell flipflop125 (
    .d (net480),
    .clk (net85),
    .q (net277)
  );
  dff_cell flipflop126 (
    .d (net481),
    .clk (net88),
    .q (net278)
  );
  mux_cell mux242 (
    .a (net484),
    .b (net253),
    .sel (net92),
    .out (net480)
  );
  mux_cell mux243 (
    .a (net485),
    .b (net254),
    .sel (net93),
    .out (net481)
  );
  buffer_cell gate43 (
    .in (net7),
    .out (net118)
  );
  buffer_cell gate44 (
    .in (net6),
    .out (net113)
  );
  buffer_cell gate45 (
    .in (net7),
    .out (net142)
  );
  buffer_cell gate46 (
    .in (net6),
    .out (net137)
  );
  buffer_cell gate47 (
    .in (net5),
    .out (net133)
  );
  buffer_cell gate48 (
    .in (net7),
    .out (net166)
  );
  buffer_cell gate49 (
    .in (net6),
    .out (net161)
  );
  buffer_cell gate50 (
    .in (net7),
    .out (net191)
  );
  buffer_cell gate51 (
    .in (net6),
    .out (net186)
  );
  buffer_cell gate52 (
    .in (net5),
    .out (net182)
  );
  buffer_cell gate53 (
    .in (net7),
    .out (net216)
  );
  buffer_cell gate54 (
    .in (net6),
    .out (net211)
  );
  buffer_cell gate55 (
    .in (net7),
    .out (net241)
  );
  buffer_cell gate56 (
    .in (net6),
    .out (net236)
  );
  buffer_cell gate57 (
    .in (net5),
    .out (net232)
  );
  buffer_cell gate58 (
    .in (net7),
    .out (net265)
  );
  buffer_cell gate59 (
    .in (net6),
    .out (net260)
  );
  buffer_cell gate60 (
    .in (net4),
    .out (net205)
  );
  buffer_cell gate61 (
    .in (net266),
    .out (net47)
  );
  buffer_cell gate62 (
    .in (net267),
    .out (net53)
  );
  buffer_cell gate63 (
    .in (net263),
    .out (net59)
  );
  buffer_cell gate64 (
    .in (net264),
    .out (net65)
  );
  buffer_cell gate65 (
    .in (net270),
    .out (net71)
  );
  buffer_cell gate66 (
    .in (net271),
    .out (net77)
  );
  buffer_cell gate67 (
    .in (net268),
    .out (net83)
  );
  buffer_cell gate68 (
    .in (net269),
    .out (net95)
  );
  buffer_cell gate69 (
    .in (net277),
    .out (net97)
  );
endmodule
