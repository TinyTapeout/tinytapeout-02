VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO s4ga
  CLASS BLOCK ;
  FOREIGN s4ga ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 170.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.000 8.800 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.000 19.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.000 29.200 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.000 39.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.000 49.600 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.000 59.800 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.000 70.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.000 80.200 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.000 90.400 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.000 100.600 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.000 110.800 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 2.000 121.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.000 131.200 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 2.000 141.400 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 2.000 151.600 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 2.000 161.800 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.090 5.200 23.690 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.830 5.200 58.430 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.570 5.200 93.170 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.310 5.200 127.910 163.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.460 5.200 41.060 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.200 5.200 75.800 163.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.940 5.200 110.540 163.440 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 144.440 163.285 ;
      LAYER met1 ;
        RECT 5.130 1.800 144.440 166.900 ;
      LAYER met2 ;
        RECT 5.160 2.390 142.040 166.930 ;
      LAYER met3 ;
        RECT 2.000 162.200 140.695 163.365 ;
        RECT 2.400 160.800 140.695 162.200 ;
        RECT 2.000 152.000 140.695 160.800 ;
        RECT 2.400 150.600 140.695 152.000 ;
        RECT 2.000 141.800 140.695 150.600 ;
        RECT 2.400 140.400 140.695 141.800 ;
        RECT 2.000 131.600 140.695 140.400 ;
        RECT 2.400 130.200 140.695 131.600 ;
        RECT 2.000 121.400 140.695 130.200 ;
        RECT 2.400 120.000 140.695 121.400 ;
        RECT 2.000 111.200 140.695 120.000 ;
        RECT 2.400 109.800 140.695 111.200 ;
        RECT 2.000 101.000 140.695 109.800 ;
        RECT 2.400 99.600 140.695 101.000 ;
        RECT 2.000 90.800 140.695 99.600 ;
        RECT 2.400 89.400 140.695 90.800 ;
        RECT 2.000 80.600 140.695 89.400 ;
        RECT 2.400 79.200 140.695 80.600 ;
        RECT 2.000 70.400 140.695 79.200 ;
        RECT 2.400 69.000 140.695 70.400 ;
        RECT 2.000 60.200 140.695 69.000 ;
        RECT 2.400 58.800 140.695 60.200 ;
        RECT 2.000 50.000 140.695 58.800 ;
        RECT 2.400 48.600 140.695 50.000 ;
        RECT 2.000 39.800 140.695 48.600 ;
        RECT 2.400 38.400 140.695 39.800 ;
        RECT 2.000 29.600 140.695 38.400 ;
        RECT 2.400 28.200 140.695 29.600 ;
        RECT 2.000 19.400 140.695 28.200 ;
        RECT 2.400 18.000 140.695 19.400 ;
        RECT 2.000 9.200 140.695 18.000 ;
        RECT 2.400 7.800 140.695 9.200 ;
        RECT 2.000 5.275 140.695 7.800 ;
      LAYER met4 ;
        RECT 11.335 6.295 21.690 156.225 ;
        RECT 24.090 6.295 39.060 156.225 ;
        RECT 41.460 6.295 56.430 156.225 ;
        RECT 58.830 6.295 73.800 156.225 ;
        RECT 76.200 6.295 91.170 156.225 ;
        RECT 93.570 6.295 96.305 156.225 ;
  END
END s4ga
END LIBRARY

