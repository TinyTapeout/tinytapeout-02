magic
tech sky130B
magscale 1 2
timestamp 1669906243
<< viali >>
rect 4169 22593 4203 22627
rect 3985 22389 4019 22423
rect 4169 21981 4203 22015
rect 3985 21845 4019 21879
rect 4169 20417 4203 20451
rect 3985 20213 4019 20247
rect 4169 18717 4203 18751
rect 3985 18581 4019 18615
rect 1685 17697 1719 17731
rect 1869 17629 1903 17663
rect 4169 17629 4203 17663
rect 3985 17493 4019 17527
rect 1869 17221 1903 17255
rect 2145 17153 2179 17187
rect 3617 16065 3651 16099
rect 3341 15997 3375 16031
rect 4169 15453 4203 15487
rect 3985 15317 4019 15351
rect 1593 15045 1627 15079
rect 1869 14977 1903 15011
rect 2652 14977 2686 15011
rect 3065 14977 3099 15011
rect 2329 14909 2363 14943
rect 2792 14909 2826 14943
rect 4169 14773 4203 14807
rect 1732 14433 1766 14467
rect 1872 14433 1906 14467
rect 1409 14365 1443 14399
rect 2145 14365 2179 14399
rect 4169 14365 4203 14399
rect 3249 14229 3283 14263
rect 3985 14229 4019 14263
rect 2329 14025 2363 14059
rect 3846 13889 3880 13923
rect 4169 13889 4203 13923
rect 3433 13821 3467 13855
rect 3706 13823 3740 13857
rect 3893 13413 3927 13447
rect 2743 13345 2777 13379
rect 2926 13345 2960 13379
rect 2513 13277 2547 13311
rect 3249 13277 3283 13311
rect 4077 13209 4111 13243
rect 1409 13141 1443 13175
rect 2795 12937 2829 12971
rect 4169 12937 4203 12971
rect 1593 12869 1627 12903
rect 1869 12801 1903 12835
rect 3065 12801 3099 12835
rect 2329 12733 2363 12767
rect 2792 12733 2826 12767
rect 2513 12257 2547 12291
rect 2786 12257 2820 12291
rect 3249 12189 3283 12223
rect 4169 12189 4203 12223
rect 1409 12053 1443 12087
rect 2782 12053 2816 12087
rect 3985 12053 4019 12087
rect 3702 11849 3736 11883
rect 4169 11713 4203 11747
rect 3433 11645 3467 11679
rect 3706 11645 3740 11679
rect 2329 11577 2363 11611
rect 3249 11237 3283 11271
rect 2237 11101 2271 11135
rect 2513 11101 2547 11135
rect 3985 11033 4019 11067
rect 1593 10761 1627 10795
rect 4169 10761 4203 10795
rect 2697 10693 2731 10727
rect 1409 10625 1443 10659
rect 2421 10557 2455 10591
rect 2237 10081 2271 10115
rect 2513 10013 2547 10047
rect 3801 10013 3835 10047
rect 3249 9877 3283 9911
rect 3985 9877 4019 9911
rect 2703 9673 2737 9707
rect 2973 9537 3007 9571
rect 2237 9469 2271 9503
rect 2700 9469 2734 9503
rect 4077 9333 4111 9367
rect 3801 9061 3835 9095
rect 2237 8993 2271 9027
rect 2513 8925 2547 8959
rect 3985 8925 4019 8959
rect 3249 8789 3283 8823
rect 2697 8585 2731 8619
rect 1685 8449 1719 8483
rect 1961 8449 1995 8483
rect 3157 8449 3191 8483
rect 3433 8449 3467 8483
rect 4169 8313 4203 8347
rect 1593 8041 1627 8075
rect 2237 7905 2271 7939
rect 1409 7837 1443 7871
rect 2513 7837 2547 7871
rect 3249 7701 3283 7735
rect 3157 7361 3191 7395
rect 3433 7361 3467 7395
rect 4169 7157 4203 7191
rect 2053 6341 2087 6375
rect 1869 6273 1903 6307
rect 3157 6273 3191 6307
rect 3433 6273 3467 6307
rect 4169 6069 4203 6103
rect 1593 4777 1627 4811
rect 1409 4573 1443 4607
<< metal1 >>
rect 1104 22874 4876 22896
rect 1104 22822 1898 22874
rect 1950 22822 1962 22874
rect 2014 22822 2026 22874
rect 2078 22822 2090 22874
rect 2142 22822 2154 22874
rect 2206 22822 2846 22874
rect 2898 22822 2910 22874
rect 2962 22822 2974 22874
rect 3026 22822 3038 22874
rect 3090 22822 3102 22874
rect 3154 22822 3794 22874
rect 3846 22822 3858 22874
rect 3910 22822 3922 22874
rect 3974 22822 3986 22874
rect 4038 22822 4050 22874
rect 4102 22822 4876 22874
rect 1104 22800 4876 22822
rect 4154 22624 4160 22636
rect 4115 22596 4160 22624
rect 4154 22584 4160 22596
rect 4212 22584 4218 22636
rect 2774 22380 2780 22432
rect 2832 22420 2838 22432
rect 3973 22423 4031 22429
rect 3973 22420 3985 22423
rect 2832 22392 3985 22420
rect 2832 22380 2838 22392
rect 3973 22389 3985 22392
rect 4019 22389 4031 22423
rect 3973 22383 4031 22389
rect 1104 22330 4876 22352
rect 1104 22278 1424 22330
rect 1476 22278 1488 22330
rect 1540 22278 1552 22330
rect 1604 22278 1616 22330
rect 1668 22278 1680 22330
rect 1732 22278 2372 22330
rect 2424 22278 2436 22330
rect 2488 22278 2500 22330
rect 2552 22278 2564 22330
rect 2616 22278 2628 22330
rect 2680 22278 3320 22330
rect 3372 22278 3384 22330
rect 3436 22278 3448 22330
rect 3500 22278 3512 22330
rect 3564 22278 3576 22330
rect 3628 22278 4268 22330
rect 4320 22278 4332 22330
rect 4384 22278 4396 22330
rect 4448 22278 4460 22330
rect 4512 22278 4524 22330
rect 4576 22278 4876 22330
rect 1104 22256 4876 22278
rect 4157 22015 4215 22021
rect 4157 21981 4169 22015
rect 4203 22012 4215 22015
rect 4246 22012 4252 22024
rect 4203 21984 4252 22012
rect 4203 21981 4215 21984
rect 4157 21975 4215 21981
rect 4246 21972 4252 21984
rect 4304 21972 4310 22024
rect 3694 21836 3700 21888
rect 3752 21876 3758 21888
rect 3973 21879 4031 21885
rect 3973 21876 3985 21879
rect 3752 21848 3985 21876
rect 3752 21836 3758 21848
rect 3973 21845 3985 21848
rect 4019 21845 4031 21879
rect 3973 21839 4031 21845
rect 1104 21786 4876 21808
rect 1104 21734 1898 21786
rect 1950 21734 1962 21786
rect 2014 21734 2026 21786
rect 2078 21734 2090 21786
rect 2142 21734 2154 21786
rect 2206 21734 2846 21786
rect 2898 21734 2910 21786
rect 2962 21734 2974 21786
rect 3026 21734 3038 21786
rect 3090 21734 3102 21786
rect 3154 21734 3794 21786
rect 3846 21734 3858 21786
rect 3910 21734 3922 21786
rect 3974 21734 3986 21786
rect 4038 21734 4050 21786
rect 4102 21734 4876 21786
rect 1104 21712 4876 21734
rect 1104 21242 4876 21264
rect 1104 21190 1424 21242
rect 1476 21190 1488 21242
rect 1540 21190 1552 21242
rect 1604 21190 1616 21242
rect 1668 21190 1680 21242
rect 1732 21190 2372 21242
rect 2424 21190 2436 21242
rect 2488 21190 2500 21242
rect 2552 21190 2564 21242
rect 2616 21190 2628 21242
rect 2680 21190 3320 21242
rect 3372 21190 3384 21242
rect 3436 21190 3448 21242
rect 3500 21190 3512 21242
rect 3564 21190 3576 21242
rect 3628 21190 4268 21242
rect 4320 21190 4332 21242
rect 4384 21190 4396 21242
rect 4448 21190 4460 21242
rect 4512 21190 4524 21242
rect 4576 21190 4876 21242
rect 1104 21168 4876 21190
rect 1104 20698 4876 20720
rect 1104 20646 1898 20698
rect 1950 20646 1962 20698
rect 2014 20646 2026 20698
rect 2078 20646 2090 20698
rect 2142 20646 2154 20698
rect 2206 20646 2846 20698
rect 2898 20646 2910 20698
rect 2962 20646 2974 20698
rect 3026 20646 3038 20698
rect 3090 20646 3102 20698
rect 3154 20646 3794 20698
rect 3846 20646 3858 20698
rect 3910 20646 3922 20698
rect 3974 20646 3986 20698
rect 4038 20646 4050 20698
rect 4102 20646 4876 20698
rect 1104 20624 4876 20646
rect 4157 20451 4215 20457
rect 4157 20417 4169 20451
rect 4203 20448 4215 20451
rect 4706 20448 4712 20460
rect 4203 20420 4712 20448
rect 4203 20417 4215 20420
rect 4157 20411 4215 20417
rect 4706 20408 4712 20420
rect 4764 20408 4770 20460
rect 3694 20204 3700 20256
rect 3752 20244 3758 20256
rect 3973 20247 4031 20253
rect 3973 20244 3985 20247
rect 3752 20216 3985 20244
rect 3752 20204 3758 20216
rect 3973 20213 3985 20216
rect 4019 20213 4031 20247
rect 3973 20207 4031 20213
rect 1104 20154 4876 20176
rect 1104 20102 1424 20154
rect 1476 20102 1488 20154
rect 1540 20102 1552 20154
rect 1604 20102 1616 20154
rect 1668 20102 1680 20154
rect 1732 20102 2372 20154
rect 2424 20102 2436 20154
rect 2488 20102 2500 20154
rect 2552 20102 2564 20154
rect 2616 20102 2628 20154
rect 2680 20102 3320 20154
rect 3372 20102 3384 20154
rect 3436 20102 3448 20154
rect 3500 20102 3512 20154
rect 3564 20102 3576 20154
rect 3628 20102 4268 20154
rect 4320 20102 4332 20154
rect 4384 20102 4396 20154
rect 4448 20102 4460 20154
rect 4512 20102 4524 20154
rect 4576 20102 4876 20154
rect 1104 20080 4876 20102
rect 3786 19660 3792 19712
rect 3844 19700 3850 19712
rect 4890 19700 4896 19712
rect 3844 19672 4896 19700
rect 3844 19660 3850 19672
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 1104 19610 4876 19632
rect 1104 19558 1898 19610
rect 1950 19558 1962 19610
rect 2014 19558 2026 19610
rect 2078 19558 2090 19610
rect 2142 19558 2154 19610
rect 2206 19558 2846 19610
rect 2898 19558 2910 19610
rect 2962 19558 2974 19610
rect 3026 19558 3038 19610
rect 3090 19558 3102 19610
rect 3154 19558 3794 19610
rect 3846 19558 3858 19610
rect 3910 19558 3922 19610
rect 3974 19558 3986 19610
rect 4038 19558 4050 19610
rect 4102 19558 4876 19610
rect 1104 19536 4876 19558
rect 1104 19066 4876 19088
rect 1104 19014 1424 19066
rect 1476 19014 1488 19066
rect 1540 19014 1552 19066
rect 1604 19014 1616 19066
rect 1668 19014 1680 19066
rect 1732 19014 2372 19066
rect 2424 19014 2436 19066
rect 2488 19014 2500 19066
rect 2552 19014 2564 19066
rect 2616 19014 2628 19066
rect 2680 19014 3320 19066
rect 3372 19014 3384 19066
rect 3436 19014 3448 19066
rect 3500 19014 3512 19066
rect 3564 19014 3576 19066
rect 3628 19014 4268 19066
rect 4320 19014 4332 19066
rect 4384 19014 4396 19066
rect 4448 19014 4460 19066
rect 4512 19014 4524 19066
rect 4576 19014 4876 19066
rect 1104 18992 4876 19014
rect 4154 18748 4160 18760
rect 4115 18720 4160 18748
rect 4154 18708 4160 18720
rect 4212 18708 4218 18760
rect 3326 18572 3332 18624
rect 3384 18612 3390 18624
rect 3973 18615 4031 18621
rect 3973 18612 3985 18615
rect 3384 18584 3985 18612
rect 3384 18572 3390 18584
rect 3973 18581 3985 18584
rect 4019 18581 4031 18615
rect 3973 18575 4031 18581
rect 1104 18522 4876 18544
rect 1104 18470 1898 18522
rect 1950 18470 1962 18522
rect 2014 18470 2026 18522
rect 2078 18470 2090 18522
rect 2142 18470 2154 18522
rect 2206 18470 2846 18522
rect 2898 18470 2910 18522
rect 2962 18470 2974 18522
rect 3026 18470 3038 18522
rect 3090 18470 3102 18522
rect 3154 18470 3794 18522
rect 3846 18470 3858 18522
rect 3910 18470 3922 18522
rect 3974 18470 3986 18522
rect 4038 18470 4050 18522
rect 4102 18470 4876 18522
rect 1104 18448 4876 18470
rect 3142 18028 3148 18080
rect 3200 18068 3206 18080
rect 3326 18068 3332 18080
rect 3200 18040 3332 18068
rect 3200 18028 3206 18040
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 1104 17978 4876 18000
rect 1104 17926 1424 17978
rect 1476 17926 1488 17978
rect 1540 17926 1552 17978
rect 1604 17926 1616 17978
rect 1668 17926 1680 17978
rect 1732 17926 2372 17978
rect 2424 17926 2436 17978
rect 2488 17926 2500 17978
rect 2552 17926 2564 17978
rect 2616 17926 2628 17978
rect 2680 17926 3320 17978
rect 3372 17926 3384 17978
rect 3436 17926 3448 17978
rect 3500 17926 3512 17978
rect 3564 17926 3576 17978
rect 3628 17926 4268 17978
rect 4320 17926 4332 17978
rect 4384 17926 4396 17978
rect 4448 17926 4460 17978
rect 4512 17926 4524 17978
rect 4576 17926 4876 17978
rect 1104 17904 4876 17926
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17728 1731 17731
rect 1762 17728 1768 17740
rect 1719 17700 1768 17728
rect 1719 17697 1731 17700
rect 1673 17691 1731 17697
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 1857 17663 1915 17669
rect 1857 17629 1869 17663
rect 1903 17660 1915 17663
rect 2222 17660 2228 17672
rect 1903 17632 2228 17660
rect 1903 17629 1915 17632
rect 1857 17623 1915 17629
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 4154 17660 4160 17672
rect 4115 17632 4160 17660
rect 4154 17620 4160 17632
rect 4212 17620 4218 17672
rect 3510 17484 3516 17536
rect 3568 17524 3574 17536
rect 3973 17527 4031 17533
rect 3973 17524 3985 17527
rect 3568 17496 3985 17524
rect 3568 17484 3574 17496
rect 3973 17493 3985 17496
rect 4019 17493 4031 17527
rect 3973 17487 4031 17493
rect 1104 17434 4876 17456
rect 1104 17382 1898 17434
rect 1950 17382 1962 17434
rect 2014 17382 2026 17434
rect 2078 17382 2090 17434
rect 2142 17382 2154 17434
rect 2206 17382 2846 17434
rect 2898 17382 2910 17434
rect 2962 17382 2974 17434
rect 3026 17382 3038 17434
rect 3090 17382 3102 17434
rect 3154 17382 3794 17434
rect 3846 17382 3858 17434
rect 3910 17382 3922 17434
rect 3974 17382 3986 17434
rect 4038 17382 4050 17434
rect 4102 17382 4876 17434
rect 1104 17360 4876 17382
rect 1857 17255 1915 17261
rect 1857 17221 1869 17255
rect 1903 17252 1915 17255
rect 3418 17252 3424 17264
rect 1903 17224 3424 17252
rect 1903 17221 1915 17224
rect 1857 17215 1915 17221
rect 3418 17212 3424 17224
rect 3476 17212 3482 17264
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17184 2191 17187
rect 2179 17156 2774 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 2746 17116 2774 17156
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 4062 17184 4068 17196
rect 3568 17156 4068 17184
rect 3568 17144 3574 17156
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 4798 17116 4804 17128
rect 2746 17088 4804 17116
rect 4798 17076 4804 17088
rect 4856 17076 4862 17128
rect 1104 16890 4876 16912
rect 1104 16838 1424 16890
rect 1476 16838 1488 16890
rect 1540 16838 1552 16890
rect 1604 16838 1616 16890
rect 1668 16838 1680 16890
rect 1732 16838 2372 16890
rect 2424 16838 2436 16890
rect 2488 16838 2500 16890
rect 2552 16838 2564 16890
rect 2616 16838 2628 16890
rect 2680 16838 3320 16890
rect 3372 16838 3384 16890
rect 3436 16838 3448 16890
rect 3500 16838 3512 16890
rect 3564 16838 3576 16890
rect 3628 16838 4268 16890
rect 4320 16838 4332 16890
rect 4384 16838 4396 16890
rect 4448 16838 4460 16890
rect 4512 16838 4524 16890
rect 4576 16838 4876 16890
rect 1104 16816 4876 16838
rect 1104 16346 4876 16368
rect 1104 16294 1898 16346
rect 1950 16294 1962 16346
rect 2014 16294 2026 16346
rect 2078 16294 2090 16346
rect 2142 16294 2154 16346
rect 2206 16294 2846 16346
rect 2898 16294 2910 16346
rect 2962 16294 2974 16346
rect 3026 16294 3038 16346
rect 3090 16294 3102 16346
rect 3154 16294 3794 16346
rect 3846 16294 3858 16346
rect 3910 16294 3922 16346
rect 3974 16294 3986 16346
rect 4038 16294 4050 16346
rect 4102 16294 4876 16346
rect 1104 16272 4876 16294
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 3786 16096 3792 16108
rect 3651 16068 3792 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 3786 16056 3792 16068
rect 3844 16056 3850 16108
rect 3329 16031 3387 16037
rect 3329 15997 3341 16031
rect 3375 16028 3387 16031
rect 4614 16028 4620 16040
rect 3375 16000 4620 16028
rect 3375 15997 3387 16000
rect 3329 15991 3387 15997
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 1104 15802 4876 15824
rect 1104 15750 1424 15802
rect 1476 15750 1488 15802
rect 1540 15750 1552 15802
rect 1604 15750 1616 15802
rect 1668 15750 1680 15802
rect 1732 15750 2372 15802
rect 2424 15750 2436 15802
rect 2488 15750 2500 15802
rect 2552 15750 2564 15802
rect 2616 15750 2628 15802
rect 2680 15750 3320 15802
rect 3372 15750 3384 15802
rect 3436 15750 3448 15802
rect 3500 15750 3512 15802
rect 3564 15750 3576 15802
rect 3628 15750 4268 15802
rect 4320 15750 4332 15802
rect 4384 15750 4396 15802
rect 4448 15750 4460 15802
rect 4512 15750 4524 15802
rect 4576 15750 4876 15802
rect 1104 15728 4876 15750
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4706 15484 4712 15496
rect 4203 15456 4712 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 3510 15376 3516 15428
rect 3568 15416 3574 15428
rect 3786 15416 3792 15428
rect 3568 15388 3792 15416
rect 3568 15376 3574 15388
rect 3786 15376 3792 15388
rect 3844 15376 3850 15428
rect 3602 15308 3608 15360
rect 3660 15348 3666 15360
rect 3973 15351 4031 15357
rect 3973 15348 3985 15351
rect 3660 15320 3985 15348
rect 3660 15308 3666 15320
rect 3973 15317 3985 15320
rect 4019 15317 4031 15351
rect 3973 15311 4031 15317
rect 1104 15258 4876 15280
rect 1104 15206 1898 15258
rect 1950 15206 1962 15258
rect 2014 15206 2026 15258
rect 2078 15206 2090 15258
rect 2142 15206 2154 15258
rect 2206 15206 2846 15258
rect 2898 15206 2910 15258
rect 2962 15206 2974 15258
rect 3026 15206 3038 15258
rect 3090 15206 3102 15258
rect 3154 15206 3794 15258
rect 3846 15206 3858 15258
rect 3910 15206 3922 15258
rect 3974 15206 3986 15258
rect 4038 15206 4050 15258
rect 4102 15206 4876 15258
rect 1104 15184 4876 15206
rect 1394 15036 1400 15088
rect 1452 15076 1458 15088
rect 1581 15079 1639 15085
rect 1581 15076 1593 15079
rect 1452 15048 1593 15076
rect 1452 15036 1458 15048
rect 1581 15045 1593 15048
rect 1627 15045 1639 15079
rect 1581 15039 1639 15045
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 15008 1915 15011
rect 2640 15011 2698 15017
rect 2640 15008 2652 15011
rect 1903 14980 2652 15008
rect 1903 14977 1915 14980
rect 1857 14971 1915 14977
rect 2640 14977 2652 14980
rect 2686 15008 2698 15011
rect 2866 15008 2872 15020
rect 2686 14980 2872 15008
rect 2686 14977 2698 14980
rect 2640 14971 2698 14977
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 3053 15011 3111 15017
rect 3053 14977 3065 15011
rect 3099 15008 3111 15011
rect 3694 15008 3700 15020
rect 3099 14980 3700 15008
rect 3099 14977 3111 14980
rect 3053 14971 3111 14977
rect 3694 14968 3700 14980
rect 3752 14968 3758 15020
rect 2222 14900 2228 14952
rect 2280 14940 2286 14952
rect 2317 14943 2375 14949
rect 2317 14940 2329 14943
rect 2280 14912 2329 14940
rect 2280 14900 2286 14912
rect 2317 14909 2329 14912
rect 2363 14909 2375 14943
rect 2317 14903 2375 14909
rect 2498 14900 2504 14952
rect 2556 14940 2562 14952
rect 2780 14943 2838 14949
rect 2780 14940 2792 14943
rect 2556 14912 2792 14940
rect 2556 14900 2562 14912
rect 2780 14909 2792 14912
rect 2826 14909 2838 14943
rect 2780 14903 2838 14909
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 2498 14804 2504 14816
rect 1820 14776 2504 14804
rect 1820 14764 1826 14776
rect 2498 14764 2504 14776
rect 2556 14764 2562 14816
rect 3510 14764 3516 14816
rect 3568 14804 3574 14816
rect 3786 14804 3792 14816
rect 3568 14776 3792 14804
rect 3568 14764 3574 14776
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 4157 14807 4215 14813
rect 4157 14773 4169 14807
rect 4203 14804 4215 14807
rect 4706 14804 4712 14816
rect 4203 14776 4712 14804
rect 4203 14773 4215 14776
rect 4157 14767 4215 14773
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 1104 14714 4876 14736
rect 1104 14662 1424 14714
rect 1476 14662 1488 14714
rect 1540 14662 1552 14714
rect 1604 14662 1616 14714
rect 1668 14662 1680 14714
rect 1732 14662 2372 14714
rect 2424 14662 2436 14714
rect 2488 14662 2500 14714
rect 2552 14662 2564 14714
rect 2616 14662 2628 14714
rect 2680 14662 3320 14714
rect 3372 14662 3384 14714
rect 3436 14662 3448 14714
rect 3500 14662 3512 14714
rect 3564 14662 3576 14714
rect 3628 14662 4268 14714
rect 4320 14662 4332 14714
rect 4384 14662 4396 14714
rect 4448 14662 4460 14714
rect 4512 14662 4524 14714
rect 4576 14662 4876 14714
rect 1104 14640 4876 14662
rect 2866 14600 2872 14612
rect 1412 14572 2872 14600
rect 1412 14464 1440 14572
rect 2866 14560 2872 14572
rect 2924 14600 2930 14612
rect 3326 14600 3332 14612
rect 2924 14572 3332 14600
rect 2924 14560 2930 14572
rect 3326 14560 3332 14572
rect 3384 14560 3390 14612
rect 1720 14467 1778 14473
rect 1720 14464 1732 14467
rect 1412 14436 1732 14464
rect 1720 14433 1732 14436
rect 1766 14433 1778 14467
rect 1720 14427 1778 14433
rect 1854 14424 1860 14476
rect 1912 14464 1918 14476
rect 2222 14464 2228 14476
rect 1912 14436 1957 14464
rect 2056 14436 2228 14464
rect 1912 14424 1918 14436
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 2056 14396 2084 14436
rect 2222 14424 2228 14436
rect 2280 14424 2286 14476
rect 1443 14368 2084 14396
rect 2133 14399 2191 14405
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2774 14396 2780 14408
rect 2179 14368 2780 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2774 14356 2780 14368
rect 2832 14356 2838 14408
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4246 14396 4252 14408
rect 4203 14368 4252 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 4246 14356 4252 14368
rect 4304 14356 4310 14408
rect 3786 14328 3792 14340
rect 3620 14300 3792 14328
rect 3620 14272 3648 14300
rect 3786 14288 3792 14300
rect 3844 14288 3850 14340
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 3237 14263 3295 14269
rect 3237 14260 3249 14263
rect 2832 14232 3249 14260
rect 2832 14220 2838 14232
rect 3237 14229 3249 14232
rect 3283 14229 3295 14263
rect 3237 14223 3295 14229
rect 3602 14220 3608 14272
rect 3660 14220 3666 14272
rect 3694 14220 3700 14272
rect 3752 14260 3758 14272
rect 3973 14263 4031 14269
rect 3973 14260 3985 14263
rect 3752 14232 3985 14260
rect 3752 14220 3758 14232
rect 3973 14229 3985 14232
rect 4019 14229 4031 14263
rect 3973 14223 4031 14229
rect 1104 14170 4876 14192
rect 1104 14118 1898 14170
rect 1950 14118 1962 14170
rect 2014 14118 2026 14170
rect 2078 14118 2090 14170
rect 2142 14118 2154 14170
rect 2206 14118 2846 14170
rect 2898 14118 2910 14170
rect 2962 14118 2974 14170
rect 3026 14118 3038 14170
rect 3090 14118 3102 14170
rect 3154 14118 3794 14170
rect 3846 14118 3858 14170
rect 3910 14118 3922 14170
rect 3974 14118 3986 14170
rect 4038 14118 4050 14170
rect 4102 14118 4876 14170
rect 1104 14096 4876 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 1670 14056 1676 14068
rect 1452 14028 1676 14056
rect 1452 14016 1458 14028
rect 1670 14016 1676 14028
rect 1728 14056 1734 14068
rect 2317 14059 2375 14065
rect 2317 14056 2329 14059
rect 1728 14028 2329 14056
rect 1728 14016 1734 14028
rect 2317 14025 2329 14028
rect 2363 14025 2375 14059
rect 2317 14019 2375 14025
rect 3050 14016 3056 14068
rect 3108 14056 3114 14068
rect 3326 14056 3332 14068
rect 3108 14028 3332 14056
rect 3108 14016 3114 14028
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 3476 14028 4200 14056
rect 3476 14016 3482 14028
rect 2222 13880 2228 13932
rect 2280 13920 2286 13932
rect 3326 13920 3332 13932
rect 2280 13892 3332 13920
rect 2280 13880 2286 13892
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 4172 13929 4200 14028
rect 3834 13923 3892 13929
rect 3834 13920 3846 13923
rect 3620 13892 3846 13920
rect 3620 13864 3648 13892
rect 3834 13889 3846 13892
rect 3880 13889 3892 13923
rect 3834 13883 3892 13889
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13889 4215 13923
rect 4157 13883 4215 13889
rect 3234 13812 3240 13864
rect 3292 13852 3298 13864
rect 3421 13855 3479 13861
rect 3421 13852 3433 13855
rect 3292 13824 3433 13852
rect 3292 13812 3298 13824
rect 3421 13821 3433 13824
rect 3467 13821 3479 13855
rect 3421 13815 3479 13821
rect 3602 13812 3608 13864
rect 3660 13812 3666 13864
rect 3694 13857 3752 13863
rect 3694 13823 3706 13857
rect 3740 13854 3752 13857
rect 3740 13852 3924 13854
rect 3740 13826 4200 13852
rect 3740 13823 3752 13826
rect 3896 13824 4200 13826
rect 3694 13817 3752 13823
rect 4172 13796 4200 13824
rect 4154 13744 4160 13796
rect 4212 13744 4218 13796
rect 3234 13676 3240 13728
rect 3292 13716 3298 13728
rect 3510 13716 3516 13728
rect 3292 13688 3516 13716
rect 3292 13676 3298 13688
rect 3510 13676 3516 13688
rect 3568 13676 3574 13728
rect 3602 13676 3608 13728
rect 3660 13716 3666 13728
rect 3970 13716 3976 13728
rect 3660 13688 3976 13716
rect 3660 13676 3666 13688
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 1104 13626 4876 13648
rect 1104 13574 1424 13626
rect 1476 13574 1488 13626
rect 1540 13574 1552 13626
rect 1604 13574 1616 13626
rect 1668 13574 1680 13626
rect 1732 13574 2372 13626
rect 2424 13574 2436 13626
rect 2488 13574 2500 13626
rect 2552 13574 2564 13626
rect 2616 13574 2628 13626
rect 2680 13574 3320 13626
rect 3372 13574 3384 13626
rect 3436 13574 3448 13626
rect 3500 13574 3512 13626
rect 3564 13574 3576 13626
rect 3628 13574 4268 13626
rect 4320 13574 4332 13626
rect 4384 13574 4396 13626
rect 4448 13574 4460 13626
rect 4512 13574 4524 13626
rect 4576 13574 4876 13626
rect 1104 13552 4876 13574
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 4890 13512 4896 13524
rect 2556 13484 4896 13512
rect 2556 13472 2562 13484
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 3881 13447 3939 13453
rect 3881 13444 3893 13447
rect 3252 13416 3893 13444
rect 2240 13348 2636 13376
rect 2240 13320 2268 13348
rect 2222 13268 2228 13320
rect 2280 13268 2286 13320
rect 2498 13308 2504 13320
rect 2459 13280 2504 13308
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 2608 13308 2636 13348
rect 2682 13336 2688 13388
rect 2740 13385 2746 13388
rect 2740 13379 2789 13385
rect 2740 13345 2743 13379
rect 2777 13376 2789 13379
rect 2914 13379 2972 13385
rect 2777 13348 2833 13376
rect 2777 13345 2789 13348
rect 2740 13339 2789 13345
rect 2914 13345 2926 13379
rect 2960 13376 2972 13379
rect 3050 13376 3056 13388
rect 2960 13348 3056 13376
rect 2960 13345 2972 13348
rect 2914 13339 2972 13345
rect 2740 13336 2746 13339
rect 3050 13336 3056 13348
rect 3108 13376 3114 13388
rect 3252 13376 3280 13416
rect 3881 13413 3893 13416
rect 3927 13413 3939 13447
rect 3881 13407 3939 13413
rect 3108 13348 3280 13376
rect 3108 13336 3114 13348
rect 3326 13336 3332 13388
rect 3384 13376 3390 13388
rect 4062 13376 4068 13388
rect 3384 13348 4068 13376
rect 3384 13336 3390 13348
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 2608 13280 3249 13308
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 3237 13271 3295 13277
rect 3510 13200 3516 13252
rect 3568 13240 3574 13252
rect 3970 13240 3976 13252
rect 3568 13212 3976 13240
rect 3568 13200 3574 13212
rect 3970 13200 3976 13212
rect 4028 13240 4034 13252
rect 4065 13243 4123 13249
rect 4065 13240 4077 13243
rect 4028 13212 4077 13240
rect 4028 13200 4034 13212
rect 4065 13209 4077 13212
rect 4111 13209 4123 13243
rect 4065 13203 4123 13209
rect 1394 13172 1400 13184
rect 1355 13144 1400 13172
rect 1394 13132 1400 13144
rect 1452 13172 1458 13184
rect 1762 13172 1768 13184
rect 1452 13144 1768 13172
rect 1452 13132 1458 13144
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 2590 13132 2596 13184
rect 2648 13172 2654 13184
rect 4522 13172 4528 13184
rect 2648 13144 4528 13172
rect 2648 13132 2654 13144
rect 4522 13132 4528 13144
rect 4580 13172 4586 13184
rect 4706 13172 4712 13184
rect 4580 13144 4712 13172
rect 4580 13132 4586 13144
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 1104 13082 4876 13104
rect 1104 13030 1898 13082
rect 1950 13030 1962 13082
rect 2014 13030 2026 13082
rect 2078 13030 2090 13082
rect 2142 13030 2154 13082
rect 2206 13030 2846 13082
rect 2898 13030 2910 13082
rect 2962 13030 2974 13082
rect 3026 13030 3038 13082
rect 3090 13030 3102 13082
rect 3154 13030 3794 13082
rect 3846 13030 3858 13082
rect 3910 13030 3922 13082
rect 3974 13030 3986 13082
rect 4038 13030 4050 13082
rect 4102 13030 4876 13082
rect 1104 13008 4876 13030
rect 2783 12971 2841 12977
rect 2783 12937 2795 12971
rect 2829 12968 2841 12971
rect 3510 12968 3516 12980
rect 2829 12940 3516 12968
rect 2829 12937 2841 12940
rect 2783 12931 2841 12937
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 4154 12968 4160 12980
rect 4115 12940 4160 12968
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 1578 12900 1584 12912
rect 1539 12872 1584 12900
rect 1578 12860 1584 12872
rect 1636 12860 1642 12912
rect 1118 12792 1124 12844
rect 1176 12832 1182 12844
rect 1857 12835 1915 12841
rect 1857 12832 1869 12835
rect 1176 12804 1869 12832
rect 1176 12792 1182 12804
rect 1857 12801 1869 12804
rect 1903 12801 1915 12835
rect 1857 12795 1915 12801
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 3326 12832 3332 12844
rect 3099 12804 3332 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 2222 12724 2228 12776
rect 2280 12764 2286 12776
rect 2317 12767 2375 12773
rect 2317 12764 2329 12767
rect 2280 12736 2329 12764
rect 2280 12724 2286 12736
rect 2317 12733 2329 12736
rect 2363 12733 2375 12767
rect 2317 12727 2375 12733
rect 2780 12767 2838 12773
rect 2780 12733 2792 12767
rect 2826 12764 2838 12767
rect 2866 12764 2872 12776
rect 2826 12736 2872 12764
rect 2826 12733 2838 12736
rect 2780 12727 2838 12733
rect 2866 12724 2872 12736
rect 2924 12724 2930 12776
rect 3510 12588 3516 12640
rect 3568 12628 3574 12640
rect 3786 12628 3792 12640
rect 3568 12600 3792 12628
rect 3568 12588 3574 12600
rect 3786 12588 3792 12600
rect 3844 12588 3850 12640
rect 1104 12538 4876 12560
rect 1104 12486 1424 12538
rect 1476 12486 1488 12538
rect 1540 12486 1552 12538
rect 1604 12486 1616 12538
rect 1668 12486 1680 12538
rect 1732 12486 2372 12538
rect 2424 12486 2436 12538
rect 2488 12486 2500 12538
rect 2552 12486 2564 12538
rect 2616 12486 2628 12538
rect 2680 12486 3320 12538
rect 3372 12486 3384 12538
rect 3436 12486 3448 12538
rect 3500 12486 3512 12538
rect 3564 12486 3576 12538
rect 3628 12486 4268 12538
rect 4320 12486 4332 12538
rect 4384 12486 4396 12538
rect 4448 12486 4460 12538
rect 4512 12486 4524 12538
rect 4576 12486 4876 12538
rect 1104 12464 4876 12486
rect 2498 12384 2504 12436
rect 2556 12424 2562 12436
rect 3694 12424 3700 12436
rect 2556 12396 3700 12424
rect 2556 12384 2562 12396
rect 3694 12384 3700 12396
rect 3752 12384 3758 12436
rect 2498 12288 2504 12300
rect 2459 12260 2504 12288
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 2774 12291 2832 12297
rect 2774 12257 2786 12291
rect 2820 12288 2832 12291
rect 3602 12288 3608 12300
rect 2820 12260 3608 12288
rect 2820 12257 2832 12260
rect 2774 12251 2832 12257
rect 3602 12248 3608 12260
rect 3660 12248 3666 12300
rect 2590 12180 2596 12232
rect 2648 12220 2654 12232
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 2648 12192 3249 12220
rect 2648 12180 2654 12192
rect 3237 12189 3249 12192
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4157 12223 4215 12229
rect 4157 12220 4169 12223
rect 4120 12192 4169 12220
rect 4120 12180 4126 12192
rect 4157 12189 4169 12192
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 4706 12152 4712 12164
rect 3160 12124 4712 12152
rect 1394 12084 1400 12096
rect 1355 12056 1400 12084
rect 1394 12044 1400 12056
rect 1452 12044 1458 12096
rect 2770 12087 2828 12093
rect 2770 12053 2782 12087
rect 2816 12084 2828 12087
rect 3160 12084 3188 12124
rect 4706 12112 4712 12124
rect 4764 12112 4770 12164
rect 2816 12056 3188 12084
rect 2816 12053 2828 12056
rect 2770 12047 2828 12053
rect 3326 12044 3332 12096
rect 3384 12084 3390 12096
rect 3973 12087 4031 12093
rect 3973 12084 3985 12087
rect 3384 12056 3985 12084
rect 3384 12044 3390 12056
rect 3973 12053 3985 12056
rect 4019 12053 4031 12087
rect 3973 12047 4031 12053
rect 1104 11994 4876 12016
rect 1104 11942 1898 11994
rect 1950 11942 1962 11994
rect 2014 11942 2026 11994
rect 2078 11942 2090 11994
rect 2142 11942 2154 11994
rect 2206 11942 2846 11994
rect 2898 11942 2910 11994
rect 2962 11942 2974 11994
rect 3026 11942 3038 11994
rect 3090 11942 3102 11994
rect 3154 11942 3794 11994
rect 3846 11942 3858 11994
rect 3910 11942 3922 11994
rect 3974 11942 3986 11994
rect 4038 11942 4050 11994
rect 4102 11942 4876 11994
rect 1104 11920 4876 11942
rect 3142 11840 3148 11892
rect 3200 11880 3206 11892
rect 3326 11880 3332 11892
rect 3200 11852 3332 11880
rect 3200 11840 3206 11852
rect 3326 11840 3332 11852
rect 3384 11840 3390 11892
rect 3694 11889 3700 11892
rect 3690 11843 3700 11889
rect 3752 11880 3758 11892
rect 3752 11852 3790 11880
rect 3694 11840 3700 11843
rect 3752 11840 3758 11852
rect 2222 11704 2228 11756
rect 2280 11744 2286 11756
rect 2590 11744 2596 11756
rect 2280 11716 2596 11744
rect 2280 11704 2286 11716
rect 2590 11704 2596 11716
rect 2648 11744 2654 11756
rect 4157 11747 4215 11753
rect 4157 11744 4169 11747
rect 2648 11716 4169 11744
rect 2648 11704 2654 11716
rect 4157 11713 4169 11716
rect 4203 11713 4215 11747
rect 4157 11707 4215 11713
rect 3234 11636 3240 11688
rect 3292 11676 3298 11688
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 3292 11648 3433 11676
rect 3292 11636 3298 11648
rect 3421 11645 3433 11648
rect 3467 11645 3479 11679
rect 3421 11639 3479 11645
rect 3602 11636 3608 11688
rect 3660 11676 3666 11688
rect 3694 11679 3752 11685
rect 3694 11676 3706 11679
rect 3660 11648 3706 11676
rect 3660 11636 3666 11648
rect 3694 11645 3706 11648
rect 3740 11645 3752 11679
rect 3694 11639 3752 11645
rect 1302 11568 1308 11620
rect 1360 11608 1366 11620
rect 2314 11608 2320 11620
rect 1360 11580 2320 11608
rect 1360 11568 1366 11580
rect 2314 11568 2320 11580
rect 2372 11568 2378 11620
rect 1394 11500 1400 11552
rect 1452 11540 1458 11552
rect 3234 11540 3240 11552
rect 1452 11512 3240 11540
rect 1452 11500 1458 11512
rect 3234 11500 3240 11512
rect 3292 11540 3298 11552
rect 3602 11540 3608 11552
rect 3292 11512 3608 11540
rect 3292 11500 3298 11512
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 1104 11450 4876 11472
rect 1104 11398 1424 11450
rect 1476 11398 1488 11450
rect 1540 11398 1552 11450
rect 1604 11398 1616 11450
rect 1668 11398 1680 11450
rect 1732 11398 2372 11450
rect 2424 11398 2436 11450
rect 2488 11398 2500 11450
rect 2552 11398 2564 11450
rect 2616 11398 2628 11450
rect 2680 11398 3320 11450
rect 3372 11398 3384 11450
rect 3436 11398 3448 11450
rect 3500 11398 3512 11450
rect 3564 11398 3576 11450
rect 3628 11398 4268 11450
rect 4320 11398 4332 11450
rect 4384 11398 4396 11450
rect 4448 11398 4460 11450
rect 4512 11398 4524 11450
rect 4576 11398 4876 11450
rect 1104 11376 4876 11398
rect 3237 11271 3295 11277
rect 3237 11237 3249 11271
rect 3283 11268 3295 11271
rect 3418 11268 3424 11280
rect 3283 11240 3424 11268
rect 3283 11237 3295 11240
rect 3237 11231 3295 11237
rect 3418 11228 3424 11240
rect 3476 11228 3482 11280
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11101 2283 11135
rect 2225 11095 2283 11101
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11132 2559 11135
rect 2774 11132 2780 11144
rect 2547 11104 2780 11132
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 2240 11064 2268 11095
rect 2774 11092 2780 11104
rect 2832 11092 2838 11144
rect 3602 11064 3608 11076
rect 2240 11036 3608 11064
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 3694 11024 3700 11076
rect 3752 11064 3758 11076
rect 3973 11067 4031 11073
rect 3973 11064 3985 11067
rect 3752 11036 3985 11064
rect 3752 11024 3758 11036
rect 3973 11033 3985 11036
rect 4019 11033 4031 11067
rect 3973 11027 4031 11033
rect 1104 10906 4876 10928
rect 1104 10854 1898 10906
rect 1950 10854 1962 10906
rect 2014 10854 2026 10906
rect 2078 10854 2090 10906
rect 2142 10854 2154 10906
rect 2206 10854 2846 10906
rect 2898 10854 2910 10906
rect 2962 10854 2974 10906
rect 3026 10854 3038 10906
rect 3090 10854 3102 10906
rect 3154 10854 3794 10906
rect 3846 10854 3858 10906
rect 3910 10854 3922 10906
rect 3974 10854 3986 10906
rect 4038 10854 4050 10906
rect 4102 10854 4876 10906
rect 1104 10832 4876 10854
rect 1118 10752 1124 10804
rect 1176 10792 1182 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1176 10764 1593 10792
rect 1176 10752 1182 10764
rect 1581 10761 1593 10764
rect 1627 10792 1639 10795
rect 2130 10792 2136 10804
rect 1627 10764 2136 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3326 10792 3332 10804
rect 2832 10764 3332 10792
rect 2832 10752 2838 10764
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 4157 10795 4215 10801
rect 4157 10761 4169 10795
rect 4203 10792 4215 10795
rect 4798 10792 4804 10804
rect 4203 10764 4804 10792
rect 4203 10761 4215 10764
rect 4157 10755 4215 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 2682 10724 2688 10736
rect 2643 10696 2688 10724
rect 2682 10684 2688 10696
rect 2740 10684 2746 10736
rect 3694 10684 3700 10736
rect 3752 10684 3758 10736
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 2222 10548 2228 10600
rect 2280 10588 2286 10600
rect 2409 10591 2467 10597
rect 2409 10588 2421 10591
rect 2280 10560 2421 10588
rect 2280 10548 2286 10560
rect 2409 10557 2421 10560
rect 2455 10557 2467 10591
rect 2409 10551 2467 10557
rect 1104 10362 4876 10384
rect 1104 10310 1424 10362
rect 1476 10310 1488 10362
rect 1540 10310 1552 10362
rect 1604 10310 1616 10362
rect 1668 10310 1680 10362
rect 1732 10310 2372 10362
rect 2424 10310 2436 10362
rect 2488 10310 2500 10362
rect 2552 10310 2564 10362
rect 2616 10310 2628 10362
rect 2680 10310 3320 10362
rect 3372 10310 3384 10362
rect 3436 10310 3448 10362
rect 3500 10310 3512 10362
rect 3564 10310 3576 10362
rect 3628 10310 4268 10362
rect 4320 10310 4332 10362
rect 4384 10310 4396 10362
rect 4448 10310 4460 10362
rect 4512 10310 4524 10362
rect 4576 10310 4876 10362
rect 1104 10288 4876 10310
rect 1302 10208 1308 10260
rect 1360 10248 1366 10260
rect 1670 10248 1676 10260
rect 1360 10220 1676 10248
rect 1360 10208 1366 10220
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 1762 10140 1768 10192
rect 1820 10140 1826 10192
rect 1780 10044 1808 10140
rect 2130 10072 2136 10124
rect 2188 10112 2194 10124
rect 2225 10115 2283 10121
rect 2225 10112 2237 10115
rect 2188 10084 2237 10112
rect 2188 10072 2194 10084
rect 2225 10081 2237 10084
rect 2271 10081 2283 10115
rect 4706 10112 4712 10124
rect 2225 10075 2283 10081
rect 2792 10084 4712 10112
rect 2792 10056 2820 10084
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 2501 10047 2559 10053
rect 2501 10044 2513 10047
rect 1780 10016 2513 10044
rect 2501 10013 2513 10016
rect 2547 10013 2559 10047
rect 2501 10007 2559 10013
rect 2590 10004 2596 10056
rect 2648 10044 2654 10056
rect 2774 10044 2780 10056
rect 2648 10016 2780 10044
rect 2648 10004 2654 10016
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 2130 9936 2136 9988
rect 2188 9976 2194 9988
rect 3804 9976 3832 10007
rect 2188 9948 3832 9976
rect 2188 9936 2194 9948
rect 3234 9908 3240 9920
rect 3195 9880 3240 9908
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 3694 9868 3700 9920
rect 3752 9908 3758 9920
rect 3973 9911 4031 9917
rect 3973 9908 3985 9911
rect 3752 9880 3985 9908
rect 3752 9868 3758 9880
rect 3973 9877 3985 9880
rect 4019 9877 4031 9911
rect 3973 9871 4031 9877
rect 1104 9818 4876 9840
rect 1104 9766 1898 9818
rect 1950 9766 1962 9818
rect 2014 9766 2026 9818
rect 2078 9766 2090 9818
rect 2142 9766 2154 9818
rect 2206 9766 2846 9818
rect 2898 9766 2910 9818
rect 2962 9766 2974 9818
rect 3026 9766 3038 9818
rect 3090 9766 3102 9818
rect 3154 9766 3794 9818
rect 3846 9766 3858 9818
rect 3910 9766 3922 9818
rect 3974 9766 3986 9818
rect 4038 9766 4050 9818
rect 4102 9766 4876 9818
rect 1104 9744 4876 9766
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 2691 9707 2749 9713
rect 2691 9704 2703 9707
rect 2556 9676 2703 9704
rect 2556 9664 2562 9676
rect 2691 9673 2703 9676
rect 2737 9673 2749 9707
rect 2691 9667 2749 9673
rect 1394 9596 1400 9648
rect 1452 9636 1458 9648
rect 1854 9636 1860 9648
rect 1452 9608 1860 9636
rect 1452 9596 1458 9608
rect 1854 9596 1860 9608
rect 1912 9596 1918 9648
rect 1946 9528 1952 9580
rect 2004 9568 2010 9580
rect 2961 9571 3019 9577
rect 2004 9540 2360 9568
rect 2004 9528 2010 9540
rect 2222 9500 2228 9512
rect 2183 9472 2228 9500
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 2332 9500 2360 9540
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 3326 9568 3332 9580
rect 3007 9540 3332 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 2688 9503 2746 9509
rect 2688 9500 2700 9503
rect 2332 9472 2700 9500
rect 2688 9469 2700 9472
rect 2734 9469 2746 9503
rect 2688 9463 2746 9469
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 4065 9367 4123 9373
rect 4065 9364 4077 9367
rect 3660 9336 4077 9364
rect 3660 9324 3666 9336
rect 4065 9333 4077 9336
rect 4111 9364 4123 9367
rect 4798 9364 4804 9376
rect 4111 9336 4804 9364
rect 4111 9333 4123 9336
rect 4065 9327 4123 9333
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 1104 9274 4876 9296
rect 1104 9222 1424 9274
rect 1476 9222 1488 9274
rect 1540 9222 1552 9274
rect 1604 9222 1616 9274
rect 1668 9222 1680 9274
rect 1732 9222 2372 9274
rect 2424 9222 2436 9274
rect 2488 9222 2500 9274
rect 2552 9222 2564 9274
rect 2616 9222 2628 9274
rect 2680 9222 3320 9274
rect 3372 9222 3384 9274
rect 3436 9222 3448 9274
rect 3500 9222 3512 9274
rect 3564 9222 3576 9274
rect 3628 9222 4268 9274
rect 4320 9222 4332 9274
rect 4384 9222 4396 9274
rect 4448 9222 4460 9274
rect 4512 9222 4524 9274
rect 4576 9222 4876 9274
rect 1104 9200 4876 9222
rect 3326 9160 3332 9172
rect 2240 9132 3332 9160
rect 2240 9033 2268 9132
rect 3326 9120 3332 9132
rect 3384 9160 3390 9172
rect 3694 9160 3700 9172
rect 3384 9132 3700 9160
rect 3384 9120 3390 9132
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 3234 9052 3240 9104
rect 3292 9092 3298 9104
rect 3789 9095 3847 9101
rect 3789 9092 3801 9095
rect 3292 9064 3801 9092
rect 3292 9052 3298 9064
rect 3789 9061 3801 9064
rect 3835 9061 3847 9095
rect 3789 9055 3847 9061
rect 2225 9027 2283 9033
rect 2225 8993 2237 9027
rect 2271 8993 2283 9027
rect 2225 8987 2283 8993
rect 1854 8916 1860 8968
rect 1912 8956 1918 8968
rect 2501 8959 2559 8965
rect 2501 8956 2513 8959
rect 1912 8928 2513 8956
rect 1912 8916 1918 8928
rect 2501 8925 2513 8928
rect 2547 8925 2559 8959
rect 2501 8919 2559 8925
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3752 8928 3985 8956
rect 3752 8916 3758 8928
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 1394 8780 1400 8832
rect 1452 8820 1458 8832
rect 1946 8820 1952 8832
rect 1452 8792 1952 8820
rect 1452 8780 1458 8792
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 3237 8823 3295 8829
rect 3237 8789 3249 8823
rect 3283 8820 3295 8823
rect 3694 8820 3700 8832
rect 3283 8792 3700 8820
rect 3283 8789 3295 8792
rect 3237 8783 3295 8789
rect 3694 8780 3700 8792
rect 3752 8780 3758 8832
rect 1104 8730 4876 8752
rect 1104 8678 1898 8730
rect 1950 8678 1962 8730
rect 2014 8678 2026 8730
rect 2078 8678 2090 8730
rect 2142 8678 2154 8730
rect 2206 8678 2846 8730
rect 2898 8678 2910 8730
rect 2962 8678 2974 8730
rect 3026 8678 3038 8730
rect 3090 8678 3102 8730
rect 3154 8678 3794 8730
rect 3846 8678 3858 8730
rect 3910 8678 3922 8730
rect 3974 8678 3986 8730
rect 4038 8678 4050 8730
rect 4102 8678 4876 8730
rect 1104 8656 4876 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 1728 8588 2697 8616
rect 1728 8576 1734 8588
rect 2685 8585 2697 8588
rect 2731 8585 2743 8619
rect 2685 8579 2743 8585
rect 3234 8548 3240 8560
rect 1688 8520 3240 8548
rect 1688 8489 1716 8520
rect 3234 8508 3240 8520
rect 3292 8508 3298 8560
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 2682 8480 2688 8492
rect 1995 8452 2688 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 3326 8480 3332 8492
rect 3191 8452 3332 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8480 3479 8483
rect 4614 8480 4620 8492
rect 3467 8452 4620 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 4157 8347 4215 8353
rect 4157 8313 4169 8347
rect 4203 8344 4215 8347
rect 4706 8344 4712 8356
rect 4203 8316 4712 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 1104 8186 4876 8208
rect 1104 8134 1424 8186
rect 1476 8134 1488 8186
rect 1540 8134 1552 8186
rect 1604 8134 1616 8186
rect 1668 8134 1680 8186
rect 1732 8134 2372 8186
rect 2424 8134 2436 8186
rect 2488 8134 2500 8186
rect 2552 8134 2564 8186
rect 2616 8134 2628 8186
rect 2680 8134 3320 8186
rect 3372 8134 3384 8186
rect 3436 8134 3448 8186
rect 3500 8134 3512 8186
rect 3564 8134 3576 8186
rect 3628 8134 4268 8186
rect 4320 8134 4332 8186
rect 4384 8134 4396 8186
rect 4448 8134 4460 8186
rect 4512 8134 4524 8186
rect 4576 8134 4876 8186
rect 1104 8112 4876 8134
rect 1210 8032 1216 8084
rect 1268 8072 1274 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 1268 8044 1593 8072
rect 1268 8032 1274 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 3234 8072 3240 8084
rect 1581 8035 1639 8041
rect 2240 8044 3240 8072
rect 2240 7945 2268 8044
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7905 2283 7939
rect 2225 7899 2283 7905
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 2501 7871 2559 7877
rect 2501 7868 2513 7871
rect 1912 7840 2513 7868
rect 1912 7828 1918 7840
rect 2501 7837 2513 7840
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 3234 7732 3240 7744
rect 3195 7704 3240 7732
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 1104 7642 4876 7664
rect 1104 7590 1898 7642
rect 1950 7590 1962 7642
rect 2014 7590 2026 7642
rect 2078 7590 2090 7642
rect 2142 7590 2154 7642
rect 2206 7590 2846 7642
rect 2898 7590 2910 7642
rect 2962 7590 2974 7642
rect 3026 7590 3038 7642
rect 3090 7590 3102 7642
rect 3154 7590 3794 7642
rect 3846 7590 3858 7642
rect 3910 7590 3922 7642
rect 3974 7590 3986 7642
rect 4038 7590 4050 7642
rect 4102 7590 4876 7642
rect 1104 7568 4876 7590
rect 3142 7392 3148 7404
rect 3055 7364 3148 7392
rect 3142 7352 3148 7364
rect 3200 7392 3206 7404
rect 3326 7392 3332 7404
rect 3200 7364 3332 7392
rect 3200 7352 3206 7364
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7392 3479 7395
rect 4154 7392 4160 7404
rect 3467 7364 4160 7392
rect 3467 7361 3479 7364
rect 3421 7355 3479 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4154 7188 4160 7200
rect 4115 7160 4160 7188
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 1104 7098 4876 7120
rect 1104 7046 1424 7098
rect 1476 7046 1488 7098
rect 1540 7046 1552 7098
rect 1604 7046 1616 7098
rect 1668 7046 1680 7098
rect 1732 7046 2372 7098
rect 2424 7046 2436 7098
rect 2488 7046 2500 7098
rect 2552 7046 2564 7098
rect 2616 7046 2628 7098
rect 2680 7046 3320 7098
rect 3372 7046 3384 7098
rect 3436 7046 3448 7098
rect 3500 7046 3512 7098
rect 3564 7046 3576 7098
rect 3628 7046 4268 7098
rect 4320 7046 4332 7098
rect 4384 7046 4396 7098
rect 4448 7046 4460 7098
rect 4512 7046 4524 7098
rect 4576 7046 4876 7098
rect 1104 7024 4876 7046
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 3326 6644 3332 6656
rect 3200 6616 3332 6644
rect 3200 6604 3206 6616
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 1104 6554 4876 6576
rect 1104 6502 1898 6554
rect 1950 6502 1962 6554
rect 2014 6502 2026 6554
rect 2078 6502 2090 6554
rect 2142 6502 2154 6554
rect 2206 6502 2846 6554
rect 2898 6502 2910 6554
rect 2962 6502 2974 6554
rect 3026 6502 3038 6554
rect 3090 6502 3102 6554
rect 3154 6502 3794 6554
rect 3846 6502 3858 6554
rect 3910 6502 3922 6554
rect 3974 6502 3986 6554
rect 4038 6502 4050 6554
rect 4102 6502 4876 6554
rect 1104 6480 4876 6502
rect 1762 6400 1768 6452
rect 1820 6440 1826 6452
rect 2130 6440 2136 6452
rect 1820 6412 2136 6440
rect 1820 6400 1826 6412
rect 2130 6400 2136 6412
rect 2188 6400 2194 6452
rect 2041 6375 2099 6381
rect 2041 6341 2053 6375
rect 2087 6372 2099 6375
rect 2222 6372 2228 6384
rect 2087 6344 2228 6372
rect 2087 6341 2099 6344
rect 2041 6335 2099 6341
rect 2222 6332 2228 6344
rect 2280 6332 2286 6384
rect 1762 6264 1768 6316
rect 1820 6304 1826 6316
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1820 6276 1869 6304
rect 1820 6264 1826 6276
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6304 3203 6307
rect 3326 6304 3332 6316
rect 3191 6276 3332 6304
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 4798 6304 4804 6316
rect 3467 6276 4804 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 4798 6264 4804 6276
rect 4856 6264 4862 6316
rect 4157 6103 4215 6109
rect 4157 6069 4169 6103
rect 4203 6100 4215 6103
rect 4706 6100 4712 6112
rect 4203 6072 4712 6100
rect 4203 6069 4215 6072
rect 4157 6063 4215 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 1104 6010 4876 6032
rect 1104 5958 1424 6010
rect 1476 5958 1488 6010
rect 1540 5958 1552 6010
rect 1604 5958 1616 6010
rect 1668 5958 1680 6010
rect 1732 5958 2372 6010
rect 2424 5958 2436 6010
rect 2488 5958 2500 6010
rect 2552 5958 2564 6010
rect 2616 5958 2628 6010
rect 2680 5958 3320 6010
rect 3372 5958 3384 6010
rect 3436 5958 3448 6010
rect 3500 5958 3512 6010
rect 3564 5958 3576 6010
rect 3628 5958 4268 6010
rect 4320 5958 4332 6010
rect 4384 5958 4396 6010
rect 4448 5958 4460 6010
rect 4512 5958 4524 6010
rect 4576 5958 4876 6010
rect 1104 5936 4876 5958
rect 1104 5466 4876 5488
rect 1104 5414 1898 5466
rect 1950 5414 1962 5466
rect 2014 5414 2026 5466
rect 2078 5414 2090 5466
rect 2142 5414 2154 5466
rect 2206 5414 2846 5466
rect 2898 5414 2910 5466
rect 2962 5414 2974 5466
rect 3026 5414 3038 5466
rect 3090 5414 3102 5466
rect 3154 5414 3794 5466
rect 3846 5414 3858 5466
rect 3910 5414 3922 5466
rect 3974 5414 3986 5466
rect 4038 5414 4050 5466
rect 4102 5414 4876 5466
rect 1104 5392 4876 5414
rect 1104 4922 4876 4944
rect 1104 4870 1424 4922
rect 1476 4870 1488 4922
rect 1540 4870 1552 4922
rect 1604 4870 1616 4922
rect 1668 4870 1680 4922
rect 1732 4870 2372 4922
rect 2424 4870 2436 4922
rect 2488 4870 2500 4922
rect 2552 4870 2564 4922
rect 2616 4870 2628 4922
rect 2680 4870 3320 4922
rect 3372 4870 3384 4922
rect 3436 4870 3448 4922
rect 3500 4870 3512 4922
rect 3564 4870 3576 4922
rect 3628 4870 4268 4922
rect 4320 4870 4332 4922
rect 4384 4870 4396 4922
rect 4448 4870 4460 4922
rect 4512 4870 4524 4922
rect 4576 4870 4876 4922
rect 1104 4848 4876 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1360 4780 1593 4808
rect 1360 4768 1366 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1581 4771 1639 4777
rect 1394 4604 1400 4616
rect 1355 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 1104 4378 4876 4400
rect 1104 4326 1898 4378
rect 1950 4326 1962 4378
rect 2014 4326 2026 4378
rect 2078 4326 2090 4378
rect 2142 4326 2154 4378
rect 2206 4326 2846 4378
rect 2898 4326 2910 4378
rect 2962 4326 2974 4378
rect 3026 4326 3038 4378
rect 3090 4326 3102 4378
rect 3154 4326 3794 4378
rect 3846 4326 3858 4378
rect 3910 4326 3922 4378
rect 3974 4326 3986 4378
rect 4038 4326 4050 4378
rect 4102 4326 4876 4378
rect 1104 4304 4876 4326
rect 1104 3834 4876 3856
rect 1104 3782 1424 3834
rect 1476 3782 1488 3834
rect 1540 3782 1552 3834
rect 1604 3782 1616 3834
rect 1668 3782 1680 3834
rect 1732 3782 2372 3834
rect 2424 3782 2436 3834
rect 2488 3782 2500 3834
rect 2552 3782 2564 3834
rect 2616 3782 2628 3834
rect 2680 3782 3320 3834
rect 3372 3782 3384 3834
rect 3436 3782 3448 3834
rect 3500 3782 3512 3834
rect 3564 3782 3576 3834
rect 3628 3782 4268 3834
rect 4320 3782 4332 3834
rect 4384 3782 4396 3834
rect 4448 3782 4460 3834
rect 4512 3782 4524 3834
rect 4576 3782 4876 3834
rect 1104 3760 4876 3782
rect 1104 3290 4876 3312
rect 1104 3238 1898 3290
rect 1950 3238 1962 3290
rect 2014 3238 2026 3290
rect 2078 3238 2090 3290
rect 2142 3238 2154 3290
rect 2206 3238 2846 3290
rect 2898 3238 2910 3290
rect 2962 3238 2974 3290
rect 3026 3238 3038 3290
rect 3090 3238 3102 3290
rect 3154 3238 3794 3290
rect 3846 3238 3858 3290
rect 3910 3238 3922 3290
rect 3974 3238 3986 3290
rect 4038 3238 4050 3290
rect 4102 3238 4876 3290
rect 1104 3216 4876 3238
rect 1104 2746 4876 2768
rect 1104 2694 1424 2746
rect 1476 2694 1488 2746
rect 1540 2694 1552 2746
rect 1604 2694 1616 2746
rect 1668 2694 1680 2746
rect 1732 2694 2372 2746
rect 2424 2694 2436 2746
rect 2488 2694 2500 2746
rect 2552 2694 2564 2746
rect 2616 2694 2628 2746
rect 2680 2694 3320 2746
rect 3372 2694 3384 2746
rect 3436 2694 3448 2746
rect 3500 2694 3512 2746
rect 3564 2694 3576 2746
rect 3628 2694 4268 2746
rect 4320 2694 4332 2746
rect 4384 2694 4396 2746
rect 4448 2694 4460 2746
rect 4512 2694 4524 2746
rect 4576 2694 4876 2746
rect 1104 2672 4876 2694
rect 1104 2202 4876 2224
rect 1104 2150 1898 2202
rect 1950 2150 1962 2202
rect 2014 2150 2026 2202
rect 2078 2150 2090 2202
rect 2142 2150 2154 2202
rect 2206 2150 2846 2202
rect 2898 2150 2910 2202
rect 2962 2150 2974 2202
rect 3026 2150 3038 2202
rect 3090 2150 3102 2202
rect 3154 2150 3794 2202
rect 3846 2150 3858 2202
rect 3910 2150 3922 2202
rect 3974 2150 3986 2202
rect 4038 2150 4050 2202
rect 4102 2150 4876 2202
rect 1104 2128 4876 2150
rect 1104 1658 4876 1680
rect 1104 1606 1424 1658
rect 1476 1606 1488 1658
rect 1540 1606 1552 1658
rect 1604 1606 1616 1658
rect 1668 1606 1680 1658
rect 1732 1606 2372 1658
rect 2424 1606 2436 1658
rect 2488 1606 2500 1658
rect 2552 1606 2564 1658
rect 2616 1606 2628 1658
rect 2680 1606 3320 1658
rect 3372 1606 3384 1658
rect 3436 1606 3448 1658
rect 3500 1606 3512 1658
rect 3564 1606 3576 1658
rect 3628 1606 4268 1658
rect 4320 1606 4332 1658
rect 4384 1606 4396 1658
rect 4448 1606 4460 1658
rect 4512 1606 4524 1658
rect 4576 1606 4876 1658
rect 1104 1584 4876 1606
rect 1104 1114 4876 1136
rect 1104 1062 1898 1114
rect 1950 1062 1962 1114
rect 2014 1062 2026 1114
rect 2078 1062 2090 1114
rect 2142 1062 2154 1114
rect 2206 1062 2846 1114
rect 2898 1062 2910 1114
rect 2962 1062 2974 1114
rect 3026 1062 3038 1114
rect 3090 1062 3102 1114
rect 3154 1062 3794 1114
rect 3846 1062 3858 1114
rect 3910 1062 3922 1114
rect 3974 1062 3986 1114
rect 4038 1062 4050 1114
rect 4102 1062 4876 1114
rect 1104 1040 4876 1062
<< via1 >>
rect 1898 22822 1950 22874
rect 1962 22822 2014 22874
rect 2026 22822 2078 22874
rect 2090 22822 2142 22874
rect 2154 22822 2206 22874
rect 2846 22822 2898 22874
rect 2910 22822 2962 22874
rect 2974 22822 3026 22874
rect 3038 22822 3090 22874
rect 3102 22822 3154 22874
rect 3794 22822 3846 22874
rect 3858 22822 3910 22874
rect 3922 22822 3974 22874
rect 3986 22822 4038 22874
rect 4050 22822 4102 22874
rect 4160 22627 4212 22636
rect 4160 22593 4169 22627
rect 4169 22593 4203 22627
rect 4203 22593 4212 22627
rect 4160 22584 4212 22593
rect 2780 22380 2832 22432
rect 1424 22278 1476 22330
rect 1488 22278 1540 22330
rect 1552 22278 1604 22330
rect 1616 22278 1668 22330
rect 1680 22278 1732 22330
rect 2372 22278 2424 22330
rect 2436 22278 2488 22330
rect 2500 22278 2552 22330
rect 2564 22278 2616 22330
rect 2628 22278 2680 22330
rect 3320 22278 3372 22330
rect 3384 22278 3436 22330
rect 3448 22278 3500 22330
rect 3512 22278 3564 22330
rect 3576 22278 3628 22330
rect 4268 22278 4320 22330
rect 4332 22278 4384 22330
rect 4396 22278 4448 22330
rect 4460 22278 4512 22330
rect 4524 22278 4576 22330
rect 4252 21972 4304 22024
rect 3700 21836 3752 21888
rect 1898 21734 1950 21786
rect 1962 21734 2014 21786
rect 2026 21734 2078 21786
rect 2090 21734 2142 21786
rect 2154 21734 2206 21786
rect 2846 21734 2898 21786
rect 2910 21734 2962 21786
rect 2974 21734 3026 21786
rect 3038 21734 3090 21786
rect 3102 21734 3154 21786
rect 3794 21734 3846 21786
rect 3858 21734 3910 21786
rect 3922 21734 3974 21786
rect 3986 21734 4038 21786
rect 4050 21734 4102 21786
rect 1424 21190 1476 21242
rect 1488 21190 1540 21242
rect 1552 21190 1604 21242
rect 1616 21190 1668 21242
rect 1680 21190 1732 21242
rect 2372 21190 2424 21242
rect 2436 21190 2488 21242
rect 2500 21190 2552 21242
rect 2564 21190 2616 21242
rect 2628 21190 2680 21242
rect 3320 21190 3372 21242
rect 3384 21190 3436 21242
rect 3448 21190 3500 21242
rect 3512 21190 3564 21242
rect 3576 21190 3628 21242
rect 4268 21190 4320 21242
rect 4332 21190 4384 21242
rect 4396 21190 4448 21242
rect 4460 21190 4512 21242
rect 4524 21190 4576 21242
rect 1898 20646 1950 20698
rect 1962 20646 2014 20698
rect 2026 20646 2078 20698
rect 2090 20646 2142 20698
rect 2154 20646 2206 20698
rect 2846 20646 2898 20698
rect 2910 20646 2962 20698
rect 2974 20646 3026 20698
rect 3038 20646 3090 20698
rect 3102 20646 3154 20698
rect 3794 20646 3846 20698
rect 3858 20646 3910 20698
rect 3922 20646 3974 20698
rect 3986 20646 4038 20698
rect 4050 20646 4102 20698
rect 4712 20408 4764 20460
rect 3700 20204 3752 20256
rect 1424 20102 1476 20154
rect 1488 20102 1540 20154
rect 1552 20102 1604 20154
rect 1616 20102 1668 20154
rect 1680 20102 1732 20154
rect 2372 20102 2424 20154
rect 2436 20102 2488 20154
rect 2500 20102 2552 20154
rect 2564 20102 2616 20154
rect 2628 20102 2680 20154
rect 3320 20102 3372 20154
rect 3384 20102 3436 20154
rect 3448 20102 3500 20154
rect 3512 20102 3564 20154
rect 3576 20102 3628 20154
rect 4268 20102 4320 20154
rect 4332 20102 4384 20154
rect 4396 20102 4448 20154
rect 4460 20102 4512 20154
rect 4524 20102 4576 20154
rect 3792 19660 3844 19712
rect 4896 19660 4948 19712
rect 1898 19558 1950 19610
rect 1962 19558 2014 19610
rect 2026 19558 2078 19610
rect 2090 19558 2142 19610
rect 2154 19558 2206 19610
rect 2846 19558 2898 19610
rect 2910 19558 2962 19610
rect 2974 19558 3026 19610
rect 3038 19558 3090 19610
rect 3102 19558 3154 19610
rect 3794 19558 3846 19610
rect 3858 19558 3910 19610
rect 3922 19558 3974 19610
rect 3986 19558 4038 19610
rect 4050 19558 4102 19610
rect 1424 19014 1476 19066
rect 1488 19014 1540 19066
rect 1552 19014 1604 19066
rect 1616 19014 1668 19066
rect 1680 19014 1732 19066
rect 2372 19014 2424 19066
rect 2436 19014 2488 19066
rect 2500 19014 2552 19066
rect 2564 19014 2616 19066
rect 2628 19014 2680 19066
rect 3320 19014 3372 19066
rect 3384 19014 3436 19066
rect 3448 19014 3500 19066
rect 3512 19014 3564 19066
rect 3576 19014 3628 19066
rect 4268 19014 4320 19066
rect 4332 19014 4384 19066
rect 4396 19014 4448 19066
rect 4460 19014 4512 19066
rect 4524 19014 4576 19066
rect 4160 18751 4212 18760
rect 4160 18717 4169 18751
rect 4169 18717 4203 18751
rect 4203 18717 4212 18751
rect 4160 18708 4212 18717
rect 3332 18572 3384 18624
rect 1898 18470 1950 18522
rect 1962 18470 2014 18522
rect 2026 18470 2078 18522
rect 2090 18470 2142 18522
rect 2154 18470 2206 18522
rect 2846 18470 2898 18522
rect 2910 18470 2962 18522
rect 2974 18470 3026 18522
rect 3038 18470 3090 18522
rect 3102 18470 3154 18522
rect 3794 18470 3846 18522
rect 3858 18470 3910 18522
rect 3922 18470 3974 18522
rect 3986 18470 4038 18522
rect 4050 18470 4102 18522
rect 3148 18028 3200 18080
rect 3332 18028 3384 18080
rect 1424 17926 1476 17978
rect 1488 17926 1540 17978
rect 1552 17926 1604 17978
rect 1616 17926 1668 17978
rect 1680 17926 1732 17978
rect 2372 17926 2424 17978
rect 2436 17926 2488 17978
rect 2500 17926 2552 17978
rect 2564 17926 2616 17978
rect 2628 17926 2680 17978
rect 3320 17926 3372 17978
rect 3384 17926 3436 17978
rect 3448 17926 3500 17978
rect 3512 17926 3564 17978
rect 3576 17926 3628 17978
rect 4268 17926 4320 17978
rect 4332 17926 4384 17978
rect 4396 17926 4448 17978
rect 4460 17926 4512 17978
rect 4524 17926 4576 17978
rect 1768 17688 1820 17740
rect 2228 17620 2280 17672
rect 4160 17663 4212 17672
rect 4160 17629 4169 17663
rect 4169 17629 4203 17663
rect 4203 17629 4212 17663
rect 4160 17620 4212 17629
rect 3516 17484 3568 17536
rect 1898 17382 1950 17434
rect 1962 17382 2014 17434
rect 2026 17382 2078 17434
rect 2090 17382 2142 17434
rect 2154 17382 2206 17434
rect 2846 17382 2898 17434
rect 2910 17382 2962 17434
rect 2974 17382 3026 17434
rect 3038 17382 3090 17434
rect 3102 17382 3154 17434
rect 3794 17382 3846 17434
rect 3858 17382 3910 17434
rect 3922 17382 3974 17434
rect 3986 17382 4038 17434
rect 4050 17382 4102 17434
rect 3424 17212 3476 17264
rect 3516 17144 3568 17196
rect 4068 17144 4120 17196
rect 4804 17076 4856 17128
rect 1424 16838 1476 16890
rect 1488 16838 1540 16890
rect 1552 16838 1604 16890
rect 1616 16838 1668 16890
rect 1680 16838 1732 16890
rect 2372 16838 2424 16890
rect 2436 16838 2488 16890
rect 2500 16838 2552 16890
rect 2564 16838 2616 16890
rect 2628 16838 2680 16890
rect 3320 16838 3372 16890
rect 3384 16838 3436 16890
rect 3448 16838 3500 16890
rect 3512 16838 3564 16890
rect 3576 16838 3628 16890
rect 4268 16838 4320 16890
rect 4332 16838 4384 16890
rect 4396 16838 4448 16890
rect 4460 16838 4512 16890
rect 4524 16838 4576 16890
rect 1898 16294 1950 16346
rect 1962 16294 2014 16346
rect 2026 16294 2078 16346
rect 2090 16294 2142 16346
rect 2154 16294 2206 16346
rect 2846 16294 2898 16346
rect 2910 16294 2962 16346
rect 2974 16294 3026 16346
rect 3038 16294 3090 16346
rect 3102 16294 3154 16346
rect 3794 16294 3846 16346
rect 3858 16294 3910 16346
rect 3922 16294 3974 16346
rect 3986 16294 4038 16346
rect 4050 16294 4102 16346
rect 3792 16056 3844 16108
rect 4620 15988 4672 16040
rect 1424 15750 1476 15802
rect 1488 15750 1540 15802
rect 1552 15750 1604 15802
rect 1616 15750 1668 15802
rect 1680 15750 1732 15802
rect 2372 15750 2424 15802
rect 2436 15750 2488 15802
rect 2500 15750 2552 15802
rect 2564 15750 2616 15802
rect 2628 15750 2680 15802
rect 3320 15750 3372 15802
rect 3384 15750 3436 15802
rect 3448 15750 3500 15802
rect 3512 15750 3564 15802
rect 3576 15750 3628 15802
rect 4268 15750 4320 15802
rect 4332 15750 4384 15802
rect 4396 15750 4448 15802
rect 4460 15750 4512 15802
rect 4524 15750 4576 15802
rect 4712 15444 4764 15496
rect 3516 15376 3568 15428
rect 3792 15376 3844 15428
rect 3608 15308 3660 15360
rect 1898 15206 1950 15258
rect 1962 15206 2014 15258
rect 2026 15206 2078 15258
rect 2090 15206 2142 15258
rect 2154 15206 2206 15258
rect 2846 15206 2898 15258
rect 2910 15206 2962 15258
rect 2974 15206 3026 15258
rect 3038 15206 3090 15258
rect 3102 15206 3154 15258
rect 3794 15206 3846 15258
rect 3858 15206 3910 15258
rect 3922 15206 3974 15258
rect 3986 15206 4038 15258
rect 4050 15206 4102 15258
rect 1400 15036 1452 15088
rect 2872 14968 2924 15020
rect 3700 14968 3752 15020
rect 2228 14900 2280 14952
rect 2504 14900 2556 14952
rect 1768 14764 1820 14816
rect 2504 14764 2556 14816
rect 3516 14764 3568 14816
rect 3792 14764 3844 14816
rect 4712 14764 4764 14816
rect 1424 14662 1476 14714
rect 1488 14662 1540 14714
rect 1552 14662 1604 14714
rect 1616 14662 1668 14714
rect 1680 14662 1732 14714
rect 2372 14662 2424 14714
rect 2436 14662 2488 14714
rect 2500 14662 2552 14714
rect 2564 14662 2616 14714
rect 2628 14662 2680 14714
rect 3320 14662 3372 14714
rect 3384 14662 3436 14714
rect 3448 14662 3500 14714
rect 3512 14662 3564 14714
rect 3576 14662 3628 14714
rect 4268 14662 4320 14714
rect 4332 14662 4384 14714
rect 4396 14662 4448 14714
rect 4460 14662 4512 14714
rect 4524 14662 4576 14714
rect 2872 14560 2924 14612
rect 3332 14560 3384 14612
rect 1860 14467 1912 14476
rect 1860 14433 1872 14467
rect 1872 14433 1906 14467
rect 1906 14433 1912 14467
rect 1860 14424 1912 14433
rect 2228 14424 2280 14476
rect 2780 14356 2832 14408
rect 4252 14356 4304 14408
rect 3792 14288 3844 14340
rect 2780 14220 2832 14272
rect 3608 14220 3660 14272
rect 3700 14220 3752 14272
rect 1898 14118 1950 14170
rect 1962 14118 2014 14170
rect 2026 14118 2078 14170
rect 2090 14118 2142 14170
rect 2154 14118 2206 14170
rect 2846 14118 2898 14170
rect 2910 14118 2962 14170
rect 2974 14118 3026 14170
rect 3038 14118 3090 14170
rect 3102 14118 3154 14170
rect 3794 14118 3846 14170
rect 3858 14118 3910 14170
rect 3922 14118 3974 14170
rect 3986 14118 4038 14170
rect 4050 14118 4102 14170
rect 1400 14016 1452 14068
rect 1676 14016 1728 14068
rect 3056 14016 3108 14068
rect 3332 14016 3384 14068
rect 3424 14016 3476 14068
rect 2228 13880 2280 13932
rect 3332 13880 3384 13932
rect 3240 13812 3292 13864
rect 3608 13812 3660 13864
rect 4160 13744 4212 13796
rect 3240 13676 3292 13728
rect 3516 13676 3568 13728
rect 3608 13676 3660 13728
rect 3976 13676 4028 13728
rect 1424 13574 1476 13626
rect 1488 13574 1540 13626
rect 1552 13574 1604 13626
rect 1616 13574 1668 13626
rect 1680 13574 1732 13626
rect 2372 13574 2424 13626
rect 2436 13574 2488 13626
rect 2500 13574 2552 13626
rect 2564 13574 2616 13626
rect 2628 13574 2680 13626
rect 3320 13574 3372 13626
rect 3384 13574 3436 13626
rect 3448 13574 3500 13626
rect 3512 13574 3564 13626
rect 3576 13574 3628 13626
rect 4268 13574 4320 13626
rect 4332 13574 4384 13626
rect 4396 13574 4448 13626
rect 4460 13574 4512 13626
rect 4524 13574 4576 13626
rect 2504 13472 2556 13524
rect 4896 13472 4948 13524
rect 2228 13268 2280 13320
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 2688 13336 2740 13388
rect 3056 13336 3108 13388
rect 3332 13336 3384 13388
rect 4068 13336 4120 13388
rect 3516 13200 3568 13252
rect 3976 13200 4028 13252
rect 1400 13175 1452 13184
rect 1400 13141 1409 13175
rect 1409 13141 1443 13175
rect 1443 13141 1452 13175
rect 1400 13132 1452 13141
rect 1768 13132 1820 13184
rect 2596 13132 2648 13184
rect 4528 13132 4580 13184
rect 4712 13132 4764 13184
rect 1898 13030 1950 13082
rect 1962 13030 2014 13082
rect 2026 13030 2078 13082
rect 2090 13030 2142 13082
rect 2154 13030 2206 13082
rect 2846 13030 2898 13082
rect 2910 13030 2962 13082
rect 2974 13030 3026 13082
rect 3038 13030 3090 13082
rect 3102 13030 3154 13082
rect 3794 13030 3846 13082
rect 3858 13030 3910 13082
rect 3922 13030 3974 13082
rect 3986 13030 4038 13082
rect 4050 13030 4102 13082
rect 3516 12928 3568 12980
rect 4160 12971 4212 12980
rect 4160 12937 4169 12971
rect 4169 12937 4203 12971
rect 4203 12937 4212 12971
rect 4160 12928 4212 12937
rect 1584 12903 1636 12912
rect 1584 12869 1593 12903
rect 1593 12869 1627 12903
rect 1627 12869 1636 12903
rect 1584 12860 1636 12869
rect 1124 12792 1176 12844
rect 3332 12792 3384 12844
rect 2228 12724 2280 12776
rect 2872 12724 2924 12776
rect 3516 12588 3568 12640
rect 3792 12588 3844 12640
rect 1424 12486 1476 12538
rect 1488 12486 1540 12538
rect 1552 12486 1604 12538
rect 1616 12486 1668 12538
rect 1680 12486 1732 12538
rect 2372 12486 2424 12538
rect 2436 12486 2488 12538
rect 2500 12486 2552 12538
rect 2564 12486 2616 12538
rect 2628 12486 2680 12538
rect 3320 12486 3372 12538
rect 3384 12486 3436 12538
rect 3448 12486 3500 12538
rect 3512 12486 3564 12538
rect 3576 12486 3628 12538
rect 4268 12486 4320 12538
rect 4332 12486 4384 12538
rect 4396 12486 4448 12538
rect 4460 12486 4512 12538
rect 4524 12486 4576 12538
rect 2504 12384 2556 12436
rect 3700 12384 3752 12436
rect 2504 12291 2556 12300
rect 2504 12257 2513 12291
rect 2513 12257 2547 12291
rect 2547 12257 2556 12291
rect 2504 12248 2556 12257
rect 3608 12248 3660 12300
rect 2596 12180 2648 12232
rect 4068 12180 4120 12232
rect 1400 12087 1452 12096
rect 1400 12053 1409 12087
rect 1409 12053 1443 12087
rect 1443 12053 1452 12087
rect 1400 12044 1452 12053
rect 4712 12112 4764 12164
rect 3332 12044 3384 12096
rect 1898 11942 1950 11994
rect 1962 11942 2014 11994
rect 2026 11942 2078 11994
rect 2090 11942 2142 11994
rect 2154 11942 2206 11994
rect 2846 11942 2898 11994
rect 2910 11942 2962 11994
rect 2974 11942 3026 11994
rect 3038 11942 3090 11994
rect 3102 11942 3154 11994
rect 3794 11942 3846 11994
rect 3858 11942 3910 11994
rect 3922 11942 3974 11994
rect 3986 11942 4038 11994
rect 4050 11942 4102 11994
rect 3148 11840 3200 11892
rect 3332 11840 3384 11892
rect 3700 11883 3752 11892
rect 3700 11849 3702 11883
rect 3702 11849 3736 11883
rect 3736 11849 3752 11883
rect 3700 11840 3752 11849
rect 2228 11704 2280 11756
rect 2596 11704 2648 11756
rect 3240 11636 3292 11688
rect 3608 11636 3660 11688
rect 1308 11568 1360 11620
rect 2320 11611 2372 11620
rect 2320 11577 2329 11611
rect 2329 11577 2363 11611
rect 2363 11577 2372 11611
rect 2320 11568 2372 11577
rect 1400 11500 1452 11552
rect 3240 11500 3292 11552
rect 3608 11500 3660 11552
rect 1424 11398 1476 11450
rect 1488 11398 1540 11450
rect 1552 11398 1604 11450
rect 1616 11398 1668 11450
rect 1680 11398 1732 11450
rect 2372 11398 2424 11450
rect 2436 11398 2488 11450
rect 2500 11398 2552 11450
rect 2564 11398 2616 11450
rect 2628 11398 2680 11450
rect 3320 11398 3372 11450
rect 3384 11398 3436 11450
rect 3448 11398 3500 11450
rect 3512 11398 3564 11450
rect 3576 11398 3628 11450
rect 4268 11398 4320 11450
rect 4332 11398 4384 11450
rect 4396 11398 4448 11450
rect 4460 11398 4512 11450
rect 4524 11398 4576 11450
rect 3424 11228 3476 11280
rect 2780 11092 2832 11144
rect 3608 11024 3660 11076
rect 3700 11024 3752 11076
rect 1898 10854 1950 10906
rect 1962 10854 2014 10906
rect 2026 10854 2078 10906
rect 2090 10854 2142 10906
rect 2154 10854 2206 10906
rect 2846 10854 2898 10906
rect 2910 10854 2962 10906
rect 2974 10854 3026 10906
rect 3038 10854 3090 10906
rect 3102 10854 3154 10906
rect 3794 10854 3846 10906
rect 3858 10854 3910 10906
rect 3922 10854 3974 10906
rect 3986 10854 4038 10906
rect 4050 10854 4102 10906
rect 1124 10752 1176 10804
rect 2136 10752 2188 10804
rect 2780 10752 2832 10804
rect 3332 10752 3384 10804
rect 4804 10752 4856 10804
rect 2688 10727 2740 10736
rect 2688 10693 2697 10727
rect 2697 10693 2731 10727
rect 2731 10693 2740 10727
rect 2688 10684 2740 10693
rect 3700 10684 3752 10736
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 2228 10548 2280 10600
rect 1424 10310 1476 10362
rect 1488 10310 1540 10362
rect 1552 10310 1604 10362
rect 1616 10310 1668 10362
rect 1680 10310 1732 10362
rect 2372 10310 2424 10362
rect 2436 10310 2488 10362
rect 2500 10310 2552 10362
rect 2564 10310 2616 10362
rect 2628 10310 2680 10362
rect 3320 10310 3372 10362
rect 3384 10310 3436 10362
rect 3448 10310 3500 10362
rect 3512 10310 3564 10362
rect 3576 10310 3628 10362
rect 4268 10310 4320 10362
rect 4332 10310 4384 10362
rect 4396 10310 4448 10362
rect 4460 10310 4512 10362
rect 4524 10310 4576 10362
rect 1308 10208 1360 10260
rect 1676 10208 1728 10260
rect 1768 10140 1820 10192
rect 2136 10072 2188 10124
rect 4712 10072 4764 10124
rect 2596 10004 2648 10056
rect 2780 10004 2832 10056
rect 2136 9936 2188 9988
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 3700 9868 3752 9920
rect 1898 9766 1950 9818
rect 1962 9766 2014 9818
rect 2026 9766 2078 9818
rect 2090 9766 2142 9818
rect 2154 9766 2206 9818
rect 2846 9766 2898 9818
rect 2910 9766 2962 9818
rect 2974 9766 3026 9818
rect 3038 9766 3090 9818
rect 3102 9766 3154 9818
rect 3794 9766 3846 9818
rect 3858 9766 3910 9818
rect 3922 9766 3974 9818
rect 3986 9766 4038 9818
rect 4050 9766 4102 9818
rect 2504 9664 2556 9716
rect 1400 9596 1452 9648
rect 1860 9596 1912 9648
rect 1952 9528 2004 9580
rect 2228 9503 2280 9512
rect 2228 9469 2237 9503
rect 2237 9469 2271 9503
rect 2271 9469 2280 9503
rect 2228 9460 2280 9469
rect 3332 9528 3384 9580
rect 3608 9324 3660 9376
rect 4804 9324 4856 9376
rect 1424 9222 1476 9274
rect 1488 9222 1540 9274
rect 1552 9222 1604 9274
rect 1616 9222 1668 9274
rect 1680 9222 1732 9274
rect 2372 9222 2424 9274
rect 2436 9222 2488 9274
rect 2500 9222 2552 9274
rect 2564 9222 2616 9274
rect 2628 9222 2680 9274
rect 3320 9222 3372 9274
rect 3384 9222 3436 9274
rect 3448 9222 3500 9274
rect 3512 9222 3564 9274
rect 3576 9222 3628 9274
rect 4268 9222 4320 9274
rect 4332 9222 4384 9274
rect 4396 9222 4448 9274
rect 4460 9222 4512 9274
rect 4524 9222 4576 9274
rect 3332 9120 3384 9172
rect 3700 9120 3752 9172
rect 3240 9052 3292 9104
rect 1860 8916 1912 8968
rect 3700 8916 3752 8968
rect 1400 8780 1452 8832
rect 1952 8780 2004 8832
rect 3700 8780 3752 8832
rect 1898 8678 1950 8730
rect 1962 8678 2014 8730
rect 2026 8678 2078 8730
rect 2090 8678 2142 8730
rect 2154 8678 2206 8730
rect 2846 8678 2898 8730
rect 2910 8678 2962 8730
rect 2974 8678 3026 8730
rect 3038 8678 3090 8730
rect 3102 8678 3154 8730
rect 3794 8678 3846 8730
rect 3858 8678 3910 8730
rect 3922 8678 3974 8730
rect 3986 8678 4038 8730
rect 4050 8678 4102 8730
rect 1676 8576 1728 8628
rect 3240 8508 3292 8560
rect 2688 8440 2740 8492
rect 3332 8440 3384 8492
rect 4620 8440 4672 8492
rect 4712 8304 4764 8356
rect 1424 8134 1476 8186
rect 1488 8134 1540 8186
rect 1552 8134 1604 8186
rect 1616 8134 1668 8186
rect 1680 8134 1732 8186
rect 2372 8134 2424 8186
rect 2436 8134 2488 8186
rect 2500 8134 2552 8186
rect 2564 8134 2616 8186
rect 2628 8134 2680 8186
rect 3320 8134 3372 8186
rect 3384 8134 3436 8186
rect 3448 8134 3500 8186
rect 3512 8134 3564 8186
rect 3576 8134 3628 8186
rect 4268 8134 4320 8186
rect 4332 8134 4384 8186
rect 4396 8134 4448 8186
rect 4460 8134 4512 8186
rect 4524 8134 4576 8186
rect 1216 8032 1268 8084
rect 3240 8032 3292 8084
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 1860 7828 1912 7880
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 1898 7590 1950 7642
rect 1962 7590 2014 7642
rect 2026 7590 2078 7642
rect 2090 7590 2142 7642
rect 2154 7590 2206 7642
rect 2846 7590 2898 7642
rect 2910 7590 2962 7642
rect 2974 7590 3026 7642
rect 3038 7590 3090 7642
rect 3102 7590 3154 7642
rect 3794 7590 3846 7642
rect 3858 7590 3910 7642
rect 3922 7590 3974 7642
rect 3986 7590 4038 7642
rect 4050 7590 4102 7642
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3332 7352 3384 7404
rect 4160 7352 4212 7404
rect 4160 7191 4212 7200
rect 4160 7157 4169 7191
rect 4169 7157 4203 7191
rect 4203 7157 4212 7191
rect 4160 7148 4212 7157
rect 1424 7046 1476 7098
rect 1488 7046 1540 7098
rect 1552 7046 1604 7098
rect 1616 7046 1668 7098
rect 1680 7046 1732 7098
rect 2372 7046 2424 7098
rect 2436 7046 2488 7098
rect 2500 7046 2552 7098
rect 2564 7046 2616 7098
rect 2628 7046 2680 7098
rect 3320 7046 3372 7098
rect 3384 7046 3436 7098
rect 3448 7046 3500 7098
rect 3512 7046 3564 7098
rect 3576 7046 3628 7098
rect 4268 7046 4320 7098
rect 4332 7046 4384 7098
rect 4396 7046 4448 7098
rect 4460 7046 4512 7098
rect 4524 7046 4576 7098
rect 3148 6604 3200 6656
rect 3332 6604 3384 6656
rect 1898 6502 1950 6554
rect 1962 6502 2014 6554
rect 2026 6502 2078 6554
rect 2090 6502 2142 6554
rect 2154 6502 2206 6554
rect 2846 6502 2898 6554
rect 2910 6502 2962 6554
rect 2974 6502 3026 6554
rect 3038 6502 3090 6554
rect 3102 6502 3154 6554
rect 3794 6502 3846 6554
rect 3858 6502 3910 6554
rect 3922 6502 3974 6554
rect 3986 6502 4038 6554
rect 4050 6502 4102 6554
rect 1768 6400 1820 6452
rect 2136 6400 2188 6452
rect 2228 6332 2280 6384
rect 1768 6264 1820 6316
rect 3332 6264 3384 6316
rect 4804 6264 4856 6316
rect 4712 6060 4764 6112
rect 1424 5958 1476 6010
rect 1488 5958 1540 6010
rect 1552 5958 1604 6010
rect 1616 5958 1668 6010
rect 1680 5958 1732 6010
rect 2372 5958 2424 6010
rect 2436 5958 2488 6010
rect 2500 5958 2552 6010
rect 2564 5958 2616 6010
rect 2628 5958 2680 6010
rect 3320 5958 3372 6010
rect 3384 5958 3436 6010
rect 3448 5958 3500 6010
rect 3512 5958 3564 6010
rect 3576 5958 3628 6010
rect 4268 5958 4320 6010
rect 4332 5958 4384 6010
rect 4396 5958 4448 6010
rect 4460 5958 4512 6010
rect 4524 5958 4576 6010
rect 1898 5414 1950 5466
rect 1962 5414 2014 5466
rect 2026 5414 2078 5466
rect 2090 5414 2142 5466
rect 2154 5414 2206 5466
rect 2846 5414 2898 5466
rect 2910 5414 2962 5466
rect 2974 5414 3026 5466
rect 3038 5414 3090 5466
rect 3102 5414 3154 5466
rect 3794 5414 3846 5466
rect 3858 5414 3910 5466
rect 3922 5414 3974 5466
rect 3986 5414 4038 5466
rect 4050 5414 4102 5466
rect 1424 4870 1476 4922
rect 1488 4870 1540 4922
rect 1552 4870 1604 4922
rect 1616 4870 1668 4922
rect 1680 4870 1732 4922
rect 2372 4870 2424 4922
rect 2436 4870 2488 4922
rect 2500 4870 2552 4922
rect 2564 4870 2616 4922
rect 2628 4870 2680 4922
rect 3320 4870 3372 4922
rect 3384 4870 3436 4922
rect 3448 4870 3500 4922
rect 3512 4870 3564 4922
rect 3576 4870 3628 4922
rect 4268 4870 4320 4922
rect 4332 4870 4384 4922
rect 4396 4870 4448 4922
rect 4460 4870 4512 4922
rect 4524 4870 4576 4922
rect 1308 4768 1360 4820
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 1898 4326 1950 4378
rect 1962 4326 2014 4378
rect 2026 4326 2078 4378
rect 2090 4326 2142 4378
rect 2154 4326 2206 4378
rect 2846 4326 2898 4378
rect 2910 4326 2962 4378
rect 2974 4326 3026 4378
rect 3038 4326 3090 4378
rect 3102 4326 3154 4378
rect 3794 4326 3846 4378
rect 3858 4326 3910 4378
rect 3922 4326 3974 4378
rect 3986 4326 4038 4378
rect 4050 4326 4102 4378
rect 1424 3782 1476 3834
rect 1488 3782 1540 3834
rect 1552 3782 1604 3834
rect 1616 3782 1668 3834
rect 1680 3782 1732 3834
rect 2372 3782 2424 3834
rect 2436 3782 2488 3834
rect 2500 3782 2552 3834
rect 2564 3782 2616 3834
rect 2628 3782 2680 3834
rect 3320 3782 3372 3834
rect 3384 3782 3436 3834
rect 3448 3782 3500 3834
rect 3512 3782 3564 3834
rect 3576 3782 3628 3834
rect 4268 3782 4320 3834
rect 4332 3782 4384 3834
rect 4396 3782 4448 3834
rect 4460 3782 4512 3834
rect 4524 3782 4576 3834
rect 1898 3238 1950 3290
rect 1962 3238 2014 3290
rect 2026 3238 2078 3290
rect 2090 3238 2142 3290
rect 2154 3238 2206 3290
rect 2846 3238 2898 3290
rect 2910 3238 2962 3290
rect 2974 3238 3026 3290
rect 3038 3238 3090 3290
rect 3102 3238 3154 3290
rect 3794 3238 3846 3290
rect 3858 3238 3910 3290
rect 3922 3238 3974 3290
rect 3986 3238 4038 3290
rect 4050 3238 4102 3290
rect 1424 2694 1476 2746
rect 1488 2694 1540 2746
rect 1552 2694 1604 2746
rect 1616 2694 1668 2746
rect 1680 2694 1732 2746
rect 2372 2694 2424 2746
rect 2436 2694 2488 2746
rect 2500 2694 2552 2746
rect 2564 2694 2616 2746
rect 2628 2694 2680 2746
rect 3320 2694 3372 2746
rect 3384 2694 3436 2746
rect 3448 2694 3500 2746
rect 3512 2694 3564 2746
rect 3576 2694 3628 2746
rect 4268 2694 4320 2746
rect 4332 2694 4384 2746
rect 4396 2694 4448 2746
rect 4460 2694 4512 2746
rect 4524 2694 4576 2746
rect 1898 2150 1950 2202
rect 1962 2150 2014 2202
rect 2026 2150 2078 2202
rect 2090 2150 2142 2202
rect 2154 2150 2206 2202
rect 2846 2150 2898 2202
rect 2910 2150 2962 2202
rect 2974 2150 3026 2202
rect 3038 2150 3090 2202
rect 3102 2150 3154 2202
rect 3794 2150 3846 2202
rect 3858 2150 3910 2202
rect 3922 2150 3974 2202
rect 3986 2150 4038 2202
rect 4050 2150 4102 2202
rect 1424 1606 1476 1658
rect 1488 1606 1540 1658
rect 1552 1606 1604 1658
rect 1616 1606 1668 1658
rect 1680 1606 1732 1658
rect 2372 1606 2424 1658
rect 2436 1606 2488 1658
rect 2500 1606 2552 1658
rect 2564 1606 2616 1658
rect 2628 1606 2680 1658
rect 3320 1606 3372 1658
rect 3384 1606 3436 1658
rect 3448 1606 3500 1658
rect 3512 1606 3564 1658
rect 3576 1606 3628 1658
rect 4268 1606 4320 1658
rect 4332 1606 4384 1658
rect 4396 1606 4448 1658
rect 4460 1606 4512 1658
rect 4524 1606 4576 1658
rect 1898 1062 1950 1114
rect 1962 1062 2014 1114
rect 2026 1062 2078 1114
rect 2090 1062 2142 1114
rect 2154 1062 2206 1114
rect 2846 1062 2898 1114
rect 2910 1062 2962 1114
rect 2974 1062 3026 1114
rect 3038 1062 3090 1114
rect 3102 1062 3154 1114
rect 3794 1062 3846 1114
rect 3858 1062 3910 1114
rect 3922 1062 3974 1114
rect 3986 1062 4038 1114
rect 4050 1062 4102 1114
<< metal2 >>
rect 4158 23216 4214 23225
rect 4158 23151 4214 23160
rect 1898 22876 2206 22885
rect 1898 22874 1904 22876
rect 1960 22874 1984 22876
rect 2040 22874 2064 22876
rect 2120 22874 2144 22876
rect 2200 22874 2206 22876
rect 1960 22822 1962 22874
rect 2142 22822 2144 22874
rect 1898 22820 1904 22822
rect 1960 22820 1984 22822
rect 2040 22820 2064 22822
rect 2120 22820 2144 22822
rect 2200 22820 2206 22822
rect 1898 22811 2206 22820
rect 2846 22876 3154 22885
rect 2846 22874 2852 22876
rect 2908 22874 2932 22876
rect 2988 22874 3012 22876
rect 3068 22874 3092 22876
rect 3148 22874 3154 22876
rect 2908 22822 2910 22874
rect 3090 22822 3092 22874
rect 2846 22820 2852 22822
rect 2908 22820 2932 22822
rect 2988 22820 3012 22822
rect 3068 22820 3092 22822
rect 3148 22820 3154 22822
rect 2846 22811 3154 22820
rect 3794 22876 4102 22885
rect 3794 22874 3800 22876
rect 3856 22874 3880 22876
rect 3936 22874 3960 22876
rect 4016 22874 4040 22876
rect 4096 22874 4102 22876
rect 3856 22822 3858 22874
rect 4038 22822 4040 22874
rect 3794 22820 3800 22822
rect 3856 22820 3880 22822
rect 3936 22820 3960 22822
rect 4016 22820 4040 22822
rect 4096 22820 4102 22822
rect 3794 22811 4102 22820
rect 4172 22642 4200 23151
rect 4160 22636 4212 22642
rect 4160 22578 4212 22584
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 1424 22332 1732 22341
rect 1424 22330 1430 22332
rect 1486 22330 1510 22332
rect 1566 22330 1590 22332
rect 1646 22330 1670 22332
rect 1726 22330 1732 22332
rect 1486 22278 1488 22330
rect 1668 22278 1670 22330
rect 1424 22276 1430 22278
rect 1486 22276 1510 22278
rect 1566 22276 1590 22278
rect 1646 22276 1670 22278
rect 1726 22276 1732 22278
rect 1424 22267 1732 22276
rect 2372 22332 2680 22341
rect 2372 22330 2378 22332
rect 2434 22330 2458 22332
rect 2514 22330 2538 22332
rect 2594 22330 2618 22332
rect 2674 22330 2680 22332
rect 2434 22278 2436 22330
rect 2616 22278 2618 22330
rect 2372 22276 2378 22278
rect 2434 22276 2458 22278
rect 2514 22276 2538 22278
rect 2594 22276 2618 22278
rect 2674 22276 2680 22278
rect 2372 22267 2680 22276
rect 1766 22128 1822 22137
rect 1766 22063 1822 22072
rect 1424 21244 1732 21253
rect 1424 21242 1430 21244
rect 1486 21242 1510 21244
rect 1566 21242 1590 21244
rect 1646 21242 1670 21244
rect 1726 21242 1732 21244
rect 1486 21190 1488 21242
rect 1668 21190 1670 21242
rect 1424 21188 1430 21190
rect 1486 21188 1510 21190
rect 1566 21188 1590 21190
rect 1646 21188 1670 21190
rect 1726 21188 1732 21190
rect 1424 21179 1732 21188
rect 1424 20156 1732 20165
rect 1424 20154 1430 20156
rect 1486 20154 1510 20156
rect 1566 20154 1590 20156
rect 1646 20154 1670 20156
rect 1726 20154 1732 20156
rect 1486 20102 1488 20154
rect 1668 20102 1670 20154
rect 1424 20100 1430 20102
rect 1486 20100 1510 20102
rect 1566 20100 1590 20102
rect 1646 20100 1670 20102
rect 1726 20100 1732 20102
rect 1424 20091 1732 20100
rect 1424 19068 1732 19077
rect 1424 19066 1430 19068
rect 1486 19066 1510 19068
rect 1566 19066 1590 19068
rect 1646 19066 1670 19068
rect 1726 19066 1732 19068
rect 1486 19014 1488 19066
rect 1668 19014 1670 19066
rect 1424 19012 1430 19014
rect 1486 19012 1510 19014
rect 1566 19012 1590 19014
rect 1646 19012 1670 19014
rect 1726 19012 1732 19014
rect 1424 19003 1732 19012
rect 1424 17980 1732 17989
rect 1424 17978 1430 17980
rect 1486 17978 1510 17980
rect 1566 17978 1590 17980
rect 1646 17978 1670 17980
rect 1726 17978 1732 17980
rect 1486 17926 1488 17978
rect 1668 17926 1670 17978
rect 1424 17924 1430 17926
rect 1486 17924 1510 17926
rect 1566 17924 1590 17926
rect 1646 17924 1670 17926
rect 1726 17924 1732 17926
rect 1424 17915 1732 17924
rect 1780 17746 1808 22063
rect 2792 21842 2820 22374
rect 3320 22332 3628 22341
rect 3320 22330 3326 22332
rect 3382 22330 3406 22332
rect 3462 22330 3486 22332
rect 3542 22330 3566 22332
rect 3622 22330 3628 22332
rect 3382 22278 3384 22330
rect 3564 22278 3566 22330
rect 3320 22276 3326 22278
rect 3382 22276 3406 22278
rect 3462 22276 3486 22278
rect 3542 22276 3566 22278
rect 3622 22276 3628 22278
rect 3320 22267 3628 22276
rect 4268 22332 4576 22341
rect 4268 22330 4274 22332
rect 4330 22330 4354 22332
rect 4410 22330 4434 22332
rect 4490 22330 4514 22332
rect 4570 22330 4576 22332
rect 4330 22278 4332 22330
rect 4512 22278 4514 22330
rect 4268 22276 4274 22278
rect 4330 22276 4354 22278
rect 4410 22276 4434 22278
rect 4490 22276 4514 22278
rect 4570 22276 4576 22278
rect 4268 22267 4576 22276
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 2700 21814 2820 21842
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 1898 21788 2206 21797
rect 1898 21786 1904 21788
rect 1960 21786 1984 21788
rect 2040 21786 2064 21788
rect 2120 21786 2144 21788
rect 2200 21786 2206 21788
rect 1960 21734 1962 21786
rect 2142 21734 2144 21786
rect 1898 21732 1904 21734
rect 1960 21732 1984 21734
rect 2040 21732 2064 21734
rect 2120 21732 2144 21734
rect 2200 21732 2206 21734
rect 1898 21723 2206 21732
rect 2700 21706 2728 21814
rect 2846 21788 3154 21797
rect 2846 21786 2852 21788
rect 2908 21786 2932 21788
rect 2988 21786 3012 21788
rect 3068 21786 3092 21788
rect 3148 21786 3154 21788
rect 2908 21734 2910 21786
rect 3090 21734 3092 21786
rect 2846 21732 2852 21734
rect 2908 21732 2932 21734
rect 2988 21732 3012 21734
rect 3068 21732 3092 21734
rect 3148 21732 3154 21734
rect 2846 21723 3154 21732
rect 2700 21678 2820 21706
rect 2372 21244 2680 21253
rect 2372 21242 2378 21244
rect 2434 21242 2458 21244
rect 2514 21242 2538 21244
rect 2594 21242 2618 21244
rect 2674 21242 2680 21244
rect 2434 21190 2436 21242
rect 2616 21190 2618 21242
rect 2372 21188 2378 21190
rect 2434 21188 2458 21190
rect 2514 21188 2538 21190
rect 2594 21188 2618 21190
rect 2674 21188 2680 21190
rect 2372 21179 2680 21188
rect 2792 20754 2820 21678
rect 3320 21244 3628 21253
rect 3320 21242 3326 21244
rect 3382 21242 3406 21244
rect 3462 21242 3486 21244
rect 3542 21242 3566 21244
rect 3622 21242 3628 21244
rect 3382 21190 3384 21242
rect 3564 21190 3566 21242
rect 3320 21188 3326 21190
rect 3382 21188 3406 21190
rect 3462 21188 3486 21190
rect 3542 21188 3566 21190
rect 3622 21188 3628 21190
rect 3320 21179 3628 21188
rect 2700 20726 2820 20754
rect 1898 20700 2206 20709
rect 1898 20698 1904 20700
rect 1960 20698 1984 20700
rect 2040 20698 2064 20700
rect 2120 20698 2144 20700
rect 2200 20698 2206 20700
rect 1960 20646 1962 20698
rect 2142 20646 2144 20698
rect 1898 20644 1904 20646
rect 1960 20644 1984 20646
rect 2040 20644 2064 20646
rect 2120 20644 2144 20646
rect 2200 20644 2206 20646
rect 1898 20635 2206 20644
rect 2700 20618 2728 20726
rect 2846 20700 3154 20709
rect 2846 20698 2852 20700
rect 2908 20698 2932 20700
rect 2988 20698 3012 20700
rect 3068 20698 3092 20700
rect 3148 20698 3154 20700
rect 2908 20646 2910 20698
rect 3090 20646 3092 20698
rect 2846 20644 2852 20646
rect 2908 20644 2932 20646
rect 2988 20644 3012 20646
rect 3068 20644 3092 20646
rect 3148 20644 3154 20646
rect 2846 20635 3154 20644
rect 2700 20590 2820 20618
rect 2372 20156 2680 20165
rect 2372 20154 2378 20156
rect 2434 20154 2458 20156
rect 2514 20154 2538 20156
rect 2594 20154 2618 20156
rect 2674 20154 2680 20156
rect 2434 20102 2436 20154
rect 2616 20102 2618 20154
rect 2372 20100 2378 20102
rect 2434 20100 2458 20102
rect 2514 20100 2538 20102
rect 2594 20100 2618 20102
rect 2674 20100 2680 20102
rect 2372 20091 2680 20100
rect 2792 19666 2820 20590
rect 3712 20482 3740 21830
rect 3794 21788 4102 21797
rect 3794 21786 3800 21788
rect 3856 21786 3880 21788
rect 3936 21786 3960 21788
rect 4016 21786 4040 21788
rect 4096 21786 4102 21788
rect 3856 21734 3858 21786
rect 4038 21734 4040 21786
rect 3794 21732 3800 21734
rect 3856 21732 3880 21734
rect 3936 21732 3960 21734
rect 4016 21732 4040 21734
rect 4096 21732 4102 21734
rect 3794 21723 4102 21732
rect 4264 21729 4292 21966
rect 4250 21720 4306 21729
rect 4250 21655 4306 21664
rect 4268 21244 4576 21253
rect 4268 21242 4274 21244
rect 4330 21242 4354 21244
rect 4410 21242 4434 21244
rect 4490 21242 4514 21244
rect 4570 21242 4576 21244
rect 4330 21190 4332 21242
rect 4512 21190 4514 21242
rect 4268 21188 4274 21190
rect 4330 21188 4354 21190
rect 4410 21188 4434 21190
rect 4490 21188 4514 21190
rect 4570 21188 4576 21190
rect 4268 21179 4576 21188
rect 3794 20700 4102 20709
rect 3794 20698 3800 20700
rect 3856 20698 3880 20700
rect 3936 20698 3960 20700
rect 4016 20698 4040 20700
rect 4096 20698 4102 20700
rect 3856 20646 3858 20698
rect 4038 20646 4040 20698
rect 3794 20644 3800 20646
rect 3856 20644 3880 20646
rect 3936 20644 3960 20646
rect 4016 20644 4040 20646
rect 4096 20644 4102 20646
rect 3794 20635 4102 20644
rect 3712 20454 3832 20482
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3320 20156 3628 20165
rect 3320 20154 3326 20156
rect 3382 20154 3406 20156
rect 3462 20154 3486 20156
rect 3542 20154 3566 20156
rect 3622 20154 3628 20156
rect 3382 20102 3384 20154
rect 3564 20102 3566 20154
rect 3320 20100 3326 20102
rect 3382 20100 3406 20102
rect 3462 20100 3486 20102
rect 3542 20100 3566 20102
rect 3622 20100 3628 20102
rect 3320 20091 3628 20100
rect 2700 19638 2820 19666
rect 1898 19612 2206 19621
rect 1898 19610 1904 19612
rect 1960 19610 1984 19612
rect 2040 19610 2064 19612
rect 2120 19610 2144 19612
rect 2200 19610 2206 19612
rect 1960 19558 1962 19610
rect 2142 19558 2144 19610
rect 1898 19556 1904 19558
rect 1960 19556 1984 19558
rect 2040 19556 2064 19558
rect 2120 19556 2144 19558
rect 2200 19556 2206 19558
rect 1898 19547 2206 19556
rect 2700 19530 2728 19638
rect 2846 19612 3154 19621
rect 2846 19610 2852 19612
rect 2908 19610 2932 19612
rect 2988 19610 3012 19612
rect 3068 19610 3092 19612
rect 3148 19610 3154 19612
rect 2908 19558 2910 19610
rect 3090 19558 3092 19610
rect 2846 19556 2852 19558
rect 2908 19556 2932 19558
rect 2988 19556 3012 19558
rect 3068 19556 3092 19558
rect 3148 19556 3154 19558
rect 2846 19547 3154 19556
rect 2700 19502 2820 19530
rect 2372 19068 2680 19077
rect 2372 19066 2378 19068
rect 2434 19066 2458 19068
rect 2514 19066 2538 19068
rect 2594 19066 2618 19068
rect 2674 19066 2680 19068
rect 2434 19014 2436 19066
rect 2616 19014 2618 19066
rect 2372 19012 2378 19014
rect 2434 19012 2458 19014
rect 2514 19012 2538 19014
rect 2594 19012 2618 19014
rect 2674 19012 2680 19014
rect 2372 19003 2680 19012
rect 2792 18578 2820 19502
rect 3238 19408 3294 19417
rect 3238 19343 3294 19352
rect 2700 18550 2820 18578
rect 1898 18524 2206 18533
rect 1898 18522 1904 18524
rect 1960 18522 1984 18524
rect 2040 18522 2064 18524
rect 2120 18522 2144 18524
rect 2200 18522 2206 18524
rect 1960 18470 1962 18522
rect 2142 18470 2144 18522
rect 1898 18468 1904 18470
rect 1960 18468 1984 18470
rect 2040 18468 2064 18470
rect 2120 18468 2144 18470
rect 2200 18468 2206 18470
rect 1898 18459 2206 18468
rect 2700 18442 2728 18550
rect 2846 18524 3154 18533
rect 2846 18522 2852 18524
rect 2908 18522 2932 18524
rect 2988 18522 3012 18524
rect 3068 18522 3092 18524
rect 3148 18522 3154 18524
rect 2908 18470 2910 18522
rect 3090 18470 3092 18522
rect 2846 18468 2852 18470
rect 2908 18468 2932 18470
rect 2988 18468 3012 18470
rect 3068 18468 3092 18470
rect 3148 18468 3154 18470
rect 2846 18459 3154 18468
rect 2700 18414 2820 18442
rect 2372 17980 2680 17989
rect 2372 17978 2378 17980
rect 2434 17978 2458 17980
rect 2514 17978 2538 17980
rect 2594 17978 2618 17980
rect 2674 17978 2680 17980
rect 2434 17926 2436 17978
rect 2616 17926 2618 17978
rect 2372 17924 2378 17926
rect 2434 17924 2458 17926
rect 2514 17924 2538 17926
rect 2594 17924 2618 17926
rect 2674 17924 2680 17926
rect 2372 17915 2680 17924
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 1898 17436 2206 17445
rect 1898 17434 1904 17436
rect 1960 17434 1984 17436
rect 2040 17434 2064 17436
rect 2120 17434 2144 17436
rect 2200 17434 2206 17436
rect 1960 17382 1962 17434
rect 2142 17382 2144 17434
rect 1898 17380 1904 17382
rect 1960 17380 1984 17382
rect 2040 17380 2064 17382
rect 2120 17380 2144 17382
rect 2200 17380 2206 17382
rect 1898 17371 2206 17380
rect 1424 16892 1732 16901
rect 1424 16890 1430 16892
rect 1486 16890 1510 16892
rect 1566 16890 1590 16892
rect 1646 16890 1670 16892
rect 1726 16890 1732 16892
rect 1486 16838 1488 16890
rect 1668 16838 1670 16890
rect 1424 16836 1430 16838
rect 1486 16836 1510 16838
rect 1566 16836 1590 16838
rect 1646 16836 1670 16838
rect 1726 16836 1732 16838
rect 1424 16827 1732 16836
rect 1306 16416 1362 16425
rect 1306 16351 1362 16360
rect 1320 15178 1348 16351
rect 1898 16348 2206 16357
rect 1898 16346 1904 16348
rect 1960 16346 1984 16348
rect 2040 16346 2064 16348
rect 2120 16346 2144 16348
rect 2200 16346 2206 16348
rect 1960 16294 1962 16346
rect 2142 16294 2144 16346
rect 1898 16292 1904 16294
rect 1960 16292 1984 16294
rect 2040 16292 2064 16294
rect 2120 16292 2144 16294
rect 2200 16292 2206 16294
rect 1898 16283 2206 16292
rect 1424 15804 1732 15813
rect 1424 15802 1430 15804
rect 1486 15802 1510 15804
rect 1566 15802 1590 15804
rect 1646 15802 1670 15804
rect 1726 15802 1732 15804
rect 1486 15750 1488 15802
rect 1668 15750 1670 15802
rect 1424 15748 1430 15750
rect 1486 15748 1510 15750
rect 1566 15748 1590 15750
rect 1646 15748 1670 15750
rect 1726 15748 1732 15750
rect 1424 15739 1732 15748
rect 1898 15260 2206 15269
rect 1898 15258 1904 15260
rect 1960 15258 1984 15260
rect 2040 15258 2064 15260
rect 2120 15258 2144 15260
rect 2200 15258 2206 15260
rect 1960 15206 1962 15258
rect 2142 15206 2144 15258
rect 1898 15204 1904 15206
rect 1960 15204 1984 15206
rect 2040 15204 2064 15206
rect 2120 15204 2144 15206
rect 2200 15204 2206 15206
rect 1898 15195 2206 15204
rect 1320 15150 1440 15178
rect 1412 15094 1440 15150
rect 1400 15088 1452 15094
rect 1400 15030 1452 15036
rect 2240 14958 2268 17614
rect 2792 17490 2820 18414
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 3160 17626 3188 18022
rect 3252 17762 3280 19343
rect 3320 19068 3628 19077
rect 3320 19066 3326 19068
rect 3382 19066 3406 19068
rect 3462 19066 3486 19068
rect 3542 19066 3566 19068
rect 3622 19066 3628 19068
rect 3382 19014 3384 19066
rect 3564 19014 3566 19066
rect 3320 19012 3326 19014
rect 3382 19012 3406 19014
rect 3462 19012 3486 19014
rect 3542 19012 3566 19014
rect 3622 19012 3628 19014
rect 3320 19003 3628 19012
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3344 18086 3372 18566
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3320 17980 3628 17989
rect 3320 17978 3326 17980
rect 3382 17978 3406 17980
rect 3462 17978 3486 17980
rect 3542 17978 3566 17980
rect 3622 17978 3628 17980
rect 3382 17926 3384 17978
rect 3564 17926 3566 17978
rect 3320 17924 3326 17926
rect 3382 17924 3406 17926
rect 3462 17924 3486 17926
rect 3542 17924 3566 17926
rect 3622 17924 3628 17926
rect 3320 17915 3628 17924
rect 3252 17734 3464 17762
rect 3160 17598 3372 17626
rect 2700 17462 2820 17490
rect 2700 17354 2728 17462
rect 2846 17436 3154 17445
rect 2846 17434 2852 17436
rect 2908 17434 2932 17436
rect 2988 17434 3012 17436
rect 3068 17434 3092 17436
rect 3148 17434 3154 17436
rect 2908 17382 2910 17434
rect 3090 17382 3092 17434
rect 2846 17380 2852 17382
rect 2908 17380 2932 17382
rect 2988 17380 3012 17382
rect 3068 17380 3092 17382
rect 3148 17380 3154 17382
rect 2846 17371 3154 17380
rect 2700 17326 2820 17354
rect 2372 16892 2680 16901
rect 2372 16890 2378 16892
rect 2434 16890 2458 16892
rect 2514 16890 2538 16892
rect 2594 16890 2618 16892
rect 2674 16890 2680 16892
rect 2434 16838 2436 16890
rect 2616 16838 2618 16890
rect 2372 16836 2378 16838
rect 2434 16836 2458 16838
rect 2514 16836 2538 16838
rect 2594 16836 2618 16838
rect 2674 16836 2680 16838
rect 2372 16827 2680 16836
rect 2792 16402 2820 17326
rect 3344 17082 3372 17598
rect 3436 17270 3464 17734
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3424 17264 3476 17270
rect 3424 17206 3476 17212
rect 3528 17202 3556 17478
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 2700 16374 2820 16402
rect 3252 17054 3372 17082
rect 2700 16266 2728 16374
rect 2846 16348 3154 16357
rect 2846 16346 2852 16348
rect 2908 16346 2932 16348
rect 2988 16346 3012 16348
rect 3068 16346 3092 16348
rect 3148 16346 3154 16348
rect 2908 16294 2910 16346
rect 3090 16294 3092 16346
rect 2846 16292 2852 16294
rect 2908 16292 2932 16294
rect 2988 16292 3012 16294
rect 3068 16292 3092 16294
rect 3148 16292 3154 16294
rect 2846 16283 3154 16292
rect 2700 16238 2820 16266
rect 2372 15804 2680 15813
rect 2372 15802 2378 15804
rect 2434 15802 2458 15804
rect 2514 15802 2538 15804
rect 2594 15802 2618 15804
rect 2674 15802 2680 15804
rect 2434 15750 2436 15802
rect 2616 15750 2618 15802
rect 2372 15748 2378 15750
rect 2434 15748 2458 15750
rect 2514 15748 2538 15750
rect 2594 15748 2618 15750
rect 2674 15748 2680 15750
rect 2372 15739 2680 15748
rect 2792 15314 2820 16238
rect 2700 15286 2820 15314
rect 2700 15178 2728 15286
rect 2846 15260 3154 15269
rect 2846 15258 2852 15260
rect 2908 15258 2932 15260
rect 2988 15258 3012 15260
rect 3068 15258 3092 15260
rect 3148 15258 3154 15260
rect 2908 15206 2910 15258
rect 3090 15206 3092 15258
rect 2846 15204 2852 15206
rect 2908 15204 2932 15206
rect 2988 15204 3012 15206
rect 3068 15204 3092 15206
rect 3148 15204 3154 15206
rect 2846 15195 3154 15204
rect 2700 15150 2820 15178
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2504 14952 2556 14958
rect 2504 14894 2556 14900
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1424 14716 1732 14725
rect 1424 14714 1430 14716
rect 1486 14714 1510 14716
rect 1566 14714 1590 14716
rect 1646 14714 1670 14716
rect 1726 14714 1732 14716
rect 1486 14662 1488 14714
rect 1668 14662 1670 14714
rect 1424 14660 1430 14662
rect 1486 14660 1510 14662
rect 1566 14660 1590 14662
rect 1646 14660 1670 14662
rect 1726 14660 1732 14662
rect 1424 14651 1732 14660
rect 1780 14498 1808 14758
rect 1688 14470 1808 14498
rect 2240 14482 2268 14894
rect 2516 14822 2544 14894
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2372 14716 2680 14725
rect 2372 14714 2378 14716
rect 2434 14714 2458 14716
rect 2514 14714 2538 14716
rect 2594 14714 2618 14716
rect 2674 14714 2680 14716
rect 2434 14662 2436 14714
rect 2616 14662 2618 14714
rect 2372 14660 2378 14662
rect 2434 14660 2458 14662
rect 2514 14660 2538 14662
rect 2594 14660 2618 14662
rect 2674 14660 2680 14662
rect 2372 14651 2680 14660
rect 1860 14476 1912 14482
rect 1688 14074 1716 14470
rect 1860 14418 1912 14424
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 1872 14362 1900 14418
rect 1780 14334 1900 14362
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1412 13818 1440 14010
rect 1320 13790 1440 13818
rect 1320 13682 1348 13790
rect 1228 13654 1348 13682
rect 1124 12844 1176 12850
rect 1124 12786 1176 12792
rect 1136 10810 1164 12786
rect 1124 10804 1176 10810
rect 1124 10746 1176 10752
rect 1228 10146 1256 13654
rect 1424 13628 1732 13637
rect 1424 13626 1430 13628
rect 1486 13626 1510 13628
rect 1566 13626 1590 13628
rect 1646 13626 1670 13628
rect 1726 13626 1732 13628
rect 1486 13574 1488 13626
rect 1668 13574 1670 13626
rect 1424 13572 1430 13574
rect 1486 13572 1510 13574
rect 1566 13572 1590 13574
rect 1646 13572 1670 13574
rect 1726 13572 1732 13574
rect 1424 13563 1732 13572
rect 1582 13424 1638 13433
rect 1582 13359 1638 13368
rect 1400 13184 1452 13190
rect 1400 13126 1452 13132
rect 1412 12730 1440 13126
rect 1596 12918 1624 13359
rect 1780 13190 1808 14334
rect 1898 14172 2206 14181
rect 1898 14170 1904 14172
rect 1960 14170 1984 14172
rect 2040 14170 2064 14172
rect 2120 14170 2144 14172
rect 2200 14170 2206 14172
rect 1960 14118 1962 14170
rect 2142 14118 2144 14170
rect 1898 14116 1904 14118
rect 1960 14116 1984 14118
rect 2040 14116 2064 14118
rect 2120 14116 2144 14118
rect 2200 14116 2206 14118
rect 1898 14107 2206 14116
rect 2240 13938 2268 14418
rect 2792 14414 2820 15150
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2884 14618 2912 14962
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2780 14272 2832 14278
rect 2700 14220 2780 14226
rect 2700 14214 2832 14220
rect 2700 14198 2820 14214
rect 2700 14090 2728 14198
rect 2846 14172 3154 14181
rect 2846 14170 2852 14172
rect 2908 14170 2932 14172
rect 2988 14170 3012 14172
rect 3068 14170 3092 14172
rect 3148 14170 3154 14172
rect 2908 14118 2910 14170
rect 3090 14118 3092 14170
rect 2846 14116 2852 14118
rect 2908 14116 2932 14118
rect 2988 14116 3012 14118
rect 3068 14116 3092 14118
rect 3148 14116 3154 14118
rect 2846 14107 3154 14116
rect 2700 14062 2820 14090
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2240 13326 2268 13874
rect 2372 13628 2680 13637
rect 2372 13626 2378 13628
rect 2434 13626 2458 13628
rect 2514 13626 2538 13628
rect 2594 13626 2618 13628
rect 2674 13626 2680 13628
rect 2434 13574 2436 13626
rect 2616 13574 2618 13626
rect 2372 13572 2378 13574
rect 2434 13572 2458 13574
rect 2514 13572 2538 13574
rect 2594 13572 2618 13574
rect 2674 13572 2680 13574
rect 2372 13563 2680 13572
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2516 13326 2544 13466
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2504 13320 2556 13326
rect 2700 13274 2728 13330
rect 2504 13262 2556 13268
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1898 13084 2206 13093
rect 1898 13082 1904 13084
rect 1960 13082 1984 13084
rect 2040 13082 2064 13084
rect 2120 13082 2144 13084
rect 2200 13082 2206 13084
rect 1960 13030 1962 13082
rect 2142 13030 2144 13082
rect 1898 13028 1904 13030
rect 1960 13028 1984 13030
rect 2040 13028 2064 13030
rect 2120 13028 2144 13030
rect 2200 13028 2206 13030
rect 1898 13019 2206 13028
rect 1584 12912 1636 12918
rect 1584 12854 1636 12860
rect 2240 12782 2268 13262
rect 2608 13246 2728 13274
rect 2608 13190 2636 13246
rect 2596 13184 2648 13190
rect 2792 13138 2820 14062
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3068 13394 3096 14010
rect 3252 13870 3280 17054
rect 3320 16892 3628 16901
rect 3320 16890 3326 16892
rect 3382 16890 3406 16892
rect 3462 16890 3486 16892
rect 3542 16890 3566 16892
rect 3622 16890 3628 16892
rect 3382 16838 3384 16890
rect 3564 16838 3566 16890
rect 3320 16836 3326 16838
rect 3382 16836 3406 16838
rect 3462 16836 3486 16838
rect 3542 16836 3566 16838
rect 3622 16836 3628 16838
rect 3320 16827 3628 16836
rect 3320 15804 3628 15813
rect 3320 15802 3326 15804
rect 3382 15802 3406 15804
rect 3462 15802 3486 15804
rect 3542 15802 3566 15804
rect 3622 15802 3628 15804
rect 3382 15750 3384 15802
rect 3564 15750 3566 15802
rect 3320 15748 3326 15750
rect 3382 15748 3406 15750
rect 3462 15748 3486 15750
rect 3542 15748 3566 15750
rect 3622 15748 3628 15750
rect 3320 15739 3628 15748
rect 3516 15428 3568 15434
rect 3516 15370 3568 15376
rect 3528 14822 3556 15370
rect 3608 15360 3660 15366
rect 3608 15302 3660 15308
rect 3516 14816 3568 14822
rect 3620 14804 3648 15302
rect 3712 15026 3740 20198
rect 3804 19718 3832 20454
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4724 20233 4752 20402
rect 4710 20224 4766 20233
rect 4268 20156 4576 20165
rect 4710 20159 4766 20168
rect 4268 20154 4274 20156
rect 4330 20154 4354 20156
rect 4410 20154 4434 20156
rect 4490 20154 4514 20156
rect 4570 20154 4576 20156
rect 4330 20102 4332 20154
rect 4512 20102 4514 20154
rect 4268 20100 4274 20102
rect 4330 20100 4354 20102
rect 4410 20100 4434 20102
rect 4490 20100 4514 20102
rect 4570 20100 4576 20102
rect 4268 20091 4576 20100
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 3794 19612 4102 19621
rect 3794 19610 3800 19612
rect 3856 19610 3880 19612
rect 3936 19610 3960 19612
rect 4016 19610 4040 19612
rect 4096 19610 4102 19612
rect 3856 19558 3858 19610
rect 4038 19558 4040 19610
rect 3794 19556 3800 19558
rect 3856 19556 3880 19558
rect 3936 19556 3960 19558
rect 4016 19556 4040 19558
rect 4096 19556 4102 19558
rect 3794 19547 4102 19556
rect 4268 19068 4576 19077
rect 4268 19066 4274 19068
rect 4330 19066 4354 19068
rect 4410 19066 4434 19068
rect 4490 19066 4514 19068
rect 4570 19066 4576 19068
rect 4330 19014 4332 19066
rect 4512 19014 4514 19066
rect 4268 19012 4274 19014
rect 4330 19012 4354 19014
rect 4410 19012 4434 19014
rect 4490 19012 4514 19014
rect 4570 19012 4576 19014
rect 4268 19003 4576 19012
rect 4160 18760 4212 18766
rect 4158 18728 4160 18737
rect 4212 18728 4214 18737
rect 4158 18663 4214 18672
rect 3794 18524 4102 18533
rect 3794 18522 3800 18524
rect 3856 18522 3880 18524
rect 3936 18522 3960 18524
rect 4016 18522 4040 18524
rect 4096 18522 4102 18524
rect 3856 18470 3858 18522
rect 4038 18470 4040 18522
rect 3794 18468 3800 18470
rect 3856 18468 3880 18470
rect 3936 18468 3960 18470
rect 4016 18468 4040 18470
rect 4096 18468 4102 18470
rect 3794 18459 4102 18468
rect 4268 17980 4576 17989
rect 4268 17978 4274 17980
rect 4330 17978 4354 17980
rect 4410 17978 4434 17980
rect 4490 17978 4514 17980
rect 4570 17978 4576 17980
rect 4330 17926 4332 17978
rect 4512 17926 4514 17978
rect 4268 17924 4274 17926
rect 4330 17924 4354 17926
rect 4410 17924 4434 17926
rect 4490 17924 4514 17926
rect 4570 17924 4576 17926
rect 4268 17915 4576 17924
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 3794 17436 4102 17445
rect 3794 17434 3800 17436
rect 3856 17434 3880 17436
rect 3936 17434 3960 17436
rect 4016 17434 4040 17436
rect 4096 17434 4102 17436
rect 3856 17382 3858 17434
rect 4038 17382 4040 17434
rect 3794 17380 3800 17382
rect 3856 17380 3880 17382
rect 3936 17380 3960 17382
rect 4016 17380 4040 17382
rect 4096 17380 4102 17382
rect 3794 17371 4102 17380
rect 4172 17241 4200 17614
rect 4158 17232 4214 17241
rect 4068 17196 4120 17202
rect 4158 17167 4214 17176
rect 4068 17138 4120 17144
rect 4080 16538 4108 17138
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4268 16892 4576 16901
rect 4268 16890 4274 16892
rect 4330 16890 4354 16892
rect 4410 16890 4434 16892
rect 4490 16890 4514 16892
rect 4570 16890 4576 16892
rect 4330 16838 4332 16890
rect 4512 16838 4514 16890
rect 4268 16836 4274 16838
rect 4330 16836 4354 16838
rect 4410 16836 4434 16838
rect 4490 16836 4514 16838
rect 4570 16836 4576 16838
rect 4268 16827 4576 16836
rect 4080 16510 4200 16538
rect 3794 16348 4102 16357
rect 3794 16346 3800 16348
rect 3856 16346 3880 16348
rect 3936 16346 3960 16348
rect 4016 16346 4040 16348
rect 4096 16346 4102 16348
rect 3856 16294 3858 16346
rect 4038 16294 4040 16346
rect 3794 16292 3800 16294
rect 3856 16292 3880 16294
rect 3936 16292 3960 16294
rect 4016 16292 4040 16294
rect 4096 16292 4102 16294
rect 3794 16283 4102 16292
rect 4172 16130 4200 16510
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 4080 16102 4200 16130
rect 3804 15434 3832 16050
rect 4080 15450 4108 16102
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4268 15804 4576 15813
rect 4268 15802 4274 15804
rect 4330 15802 4354 15804
rect 4410 15802 4434 15804
rect 4490 15802 4514 15804
rect 4570 15802 4576 15804
rect 4330 15750 4332 15802
rect 4512 15750 4514 15802
rect 4268 15748 4274 15750
rect 4330 15748 4354 15750
rect 4410 15748 4434 15750
rect 4490 15748 4514 15750
rect 4570 15748 4576 15750
rect 4268 15739 4576 15748
rect 3792 15428 3844 15434
rect 4080 15422 4200 15450
rect 3792 15370 3844 15376
rect 3794 15260 4102 15269
rect 3794 15258 3800 15260
rect 3856 15258 3880 15260
rect 3936 15258 3960 15260
rect 4016 15258 4040 15260
rect 4096 15258 4102 15260
rect 3856 15206 3858 15258
rect 4038 15206 4040 15258
rect 3794 15204 3800 15206
rect 3856 15204 3880 15206
rect 3936 15204 3960 15206
rect 4016 15204 4040 15206
rect 4096 15204 4102 15206
rect 3794 15195 4102 15204
rect 4172 15042 4200 15422
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 4080 15014 4200 15042
rect 3792 14816 3844 14822
rect 3620 14776 3740 14804
rect 3516 14758 3568 14764
rect 3320 14716 3628 14725
rect 3320 14714 3326 14716
rect 3382 14714 3406 14716
rect 3462 14714 3486 14716
rect 3542 14714 3566 14716
rect 3622 14714 3628 14716
rect 3382 14662 3384 14714
rect 3564 14662 3566 14714
rect 3320 14660 3326 14662
rect 3382 14660 3406 14662
rect 3462 14660 3486 14662
rect 3542 14660 3566 14662
rect 3622 14660 3628 14662
rect 3320 14651 3628 14660
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3344 14074 3372 14554
rect 3712 14362 3740 14776
rect 3792 14758 3844 14764
rect 3528 14334 3740 14362
rect 3804 14346 3832 14758
rect 4080 14362 4108 15014
rect 4268 14716 4576 14725
rect 4268 14714 4274 14716
rect 4330 14714 4354 14716
rect 4410 14714 4434 14716
rect 4490 14714 4514 14716
rect 4570 14714 4576 14716
rect 4330 14662 4332 14714
rect 4512 14662 4514 14714
rect 4268 14660 4274 14662
rect 4330 14660 4354 14662
rect 4410 14660 4434 14662
rect 4490 14660 4514 14662
rect 4570 14660 4576 14662
rect 4268 14651 4576 14660
rect 4252 14408 4304 14414
rect 3792 14340 3844 14346
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3436 13954 3464 14010
rect 3344 13938 3464 13954
rect 3332 13932 3464 13938
rect 3384 13926 3464 13932
rect 3332 13874 3384 13880
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3528 13734 3556 14334
rect 4080 14334 4200 14362
rect 4252 14350 4304 14356
rect 3792 14282 3844 14288
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3700 14272 3752 14278
rect 3700 14214 3752 14220
rect 3620 13870 3648 14214
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3620 13734 3648 13806
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 2596 13126 2648 13132
rect 2700 13110 2820 13138
rect 2700 13002 2728 13110
rect 2846 13084 3154 13093
rect 2846 13082 2852 13084
rect 2908 13082 2932 13084
rect 2988 13082 3012 13084
rect 3068 13082 3092 13084
rect 3148 13082 3154 13084
rect 2908 13030 2910 13082
rect 3090 13030 3092 13082
rect 2846 13028 2852 13030
rect 2908 13028 2932 13030
rect 2988 13028 3012 13030
rect 3068 13028 3092 13030
rect 3148 13028 3154 13030
rect 2846 13019 3154 13028
rect 2700 12974 2820 13002
rect 1320 12702 1440 12730
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 1320 12434 1348 12702
rect 1424 12540 1732 12549
rect 1424 12538 1430 12540
rect 1486 12538 1510 12540
rect 1566 12538 1590 12540
rect 1646 12538 1670 12540
rect 1726 12538 1732 12540
rect 1486 12486 1488 12538
rect 1668 12486 1670 12538
rect 1424 12484 1430 12486
rect 1486 12484 1510 12486
rect 1566 12484 1590 12486
rect 1646 12484 1670 12486
rect 1726 12484 1732 12486
rect 1424 12475 1732 12484
rect 1320 12406 1716 12434
rect 1688 12322 1716 12406
rect 1688 12294 1808 12322
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1308 11620 1360 11626
rect 1308 11562 1360 11568
rect 1320 10266 1348 11562
rect 1412 11558 1440 12038
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1424 11452 1732 11461
rect 1424 11450 1430 11452
rect 1486 11450 1510 11452
rect 1566 11450 1590 11452
rect 1646 11450 1670 11452
rect 1726 11450 1732 11452
rect 1486 11398 1488 11450
rect 1668 11398 1670 11450
rect 1424 11396 1430 11398
rect 1486 11396 1510 11398
rect 1566 11396 1590 11398
rect 1646 11396 1670 11398
rect 1726 11396 1732 11398
rect 1424 11387 1732 11396
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 10577 1440 10610
rect 1398 10568 1454 10577
rect 1398 10503 1454 10512
rect 1424 10364 1732 10373
rect 1424 10362 1430 10364
rect 1486 10362 1510 10364
rect 1566 10362 1590 10364
rect 1646 10362 1670 10364
rect 1726 10362 1732 10364
rect 1486 10310 1488 10362
rect 1668 10310 1670 10362
rect 1424 10308 1430 10310
rect 1486 10308 1510 10310
rect 1566 10308 1590 10310
rect 1646 10308 1670 10310
rect 1726 10308 1732 10310
rect 1424 10299 1732 10308
rect 1308 10260 1360 10266
rect 1308 10202 1360 10208
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1228 10118 1440 10146
rect 1412 9654 1440 10118
rect 1688 9674 1716 10202
rect 1780 10198 1808 12294
rect 1898 11996 2206 12005
rect 1898 11994 1904 11996
rect 1960 11994 1984 11996
rect 2040 11994 2064 11996
rect 2120 11994 2144 11996
rect 2200 11994 2206 11996
rect 1960 11942 1962 11994
rect 2142 11942 2144 11994
rect 1898 11940 1904 11942
rect 1960 11940 1984 11942
rect 2040 11940 2064 11942
rect 2120 11940 2144 11942
rect 2200 11940 2206 11942
rect 1898 11931 2206 11940
rect 2240 11762 2268 12718
rect 2372 12540 2680 12549
rect 2372 12538 2378 12540
rect 2434 12538 2458 12540
rect 2514 12538 2538 12540
rect 2594 12538 2618 12540
rect 2674 12538 2680 12540
rect 2434 12486 2436 12538
rect 2616 12486 2618 12538
rect 2372 12484 2378 12486
rect 2434 12484 2458 12486
rect 2514 12484 2538 12486
rect 2594 12484 2618 12486
rect 2674 12484 2680 12486
rect 2372 12475 2680 12484
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2318 12336 2374 12345
rect 2516 12306 2544 12378
rect 2318 12271 2374 12280
rect 2504 12300 2556 12306
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 1898 10908 2206 10917
rect 1898 10906 1904 10908
rect 1960 10906 1984 10908
rect 2040 10906 2064 10908
rect 2120 10906 2144 10908
rect 2200 10906 2206 10908
rect 1960 10854 1962 10906
rect 2142 10854 2144 10906
rect 1898 10852 1904 10854
rect 1960 10852 1984 10854
rect 2040 10852 2064 10854
rect 2120 10852 2144 10854
rect 2200 10852 2206 10854
rect 1898 10843 2206 10852
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 1768 10192 1820 10198
rect 1768 10134 1820 10140
rect 2148 10130 2176 10746
rect 2240 10606 2268 11698
rect 2332 11626 2360 12271
rect 2504 12242 2556 12248
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2608 11762 2636 12174
rect 2792 12050 2820 12974
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2884 12345 2912 12718
rect 2870 12336 2926 12345
rect 2870 12271 2926 12280
rect 2700 12022 2820 12050
rect 2700 11914 2728 12022
rect 2846 11996 3154 12005
rect 2846 11994 2852 11996
rect 2908 11994 2932 11996
rect 2988 11994 3012 11996
rect 3068 11994 3092 11996
rect 3148 11994 3154 11996
rect 2908 11942 2910 11994
rect 3090 11942 3092 11994
rect 2846 11940 2852 11942
rect 2908 11940 2932 11942
rect 2988 11940 3012 11942
rect 3068 11940 3092 11942
rect 3148 11940 3154 11942
rect 2846 11931 3154 11940
rect 2700 11886 2820 11914
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2372 11452 2680 11461
rect 2372 11450 2378 11452
rect 2434 11450 2458 11452
rect 2514 11450 2538 11452
rect 2594 11450 2618 11452
rect 2674 11450 2680 11452
rect 2434 11398 2436 11450
rect 2616 11398 2618 11450
rect 2372 11396 2378 11398
rect 2434 11396 2458 11398
rect 2514 11396 2538 11398
rect 2594 11396 2618 11398
rect 2674 11396 2680 11398
rect 2372 11387 2680 11396
rect 2792 11150 2820 11886
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 3160 11098 3188 11834
rect 3252 11694 3280 13670
rect 3320 13628 3628 13637
rect 3320 13626 3326 13628
rect 3382 13626 3406 13628
rect 3462 13626 3486 13628
rect 3542 13626 3566 13628
rect 3622 13626 3628 13628
rect 3382 13574 3384 13626
rect 3564 13574 3566 13626
rect 3320 13572 3326 13574
rect 3382 13572 3406 13574
rect 3462 13572 3486 13574
rect 3542 13572 3566 13574
rect 3622 13572 3628 13574
rect 3320 13563 3628 13572
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3344 12850 3372 13330
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3528 12986 3556 13194
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3528 12646 3556 12922
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3320 12540 3628 12549
rect 3320 12538 3326 12540
rect 3382 12538 3406 12540
rect 3462 12538 3486 12540
rect 3542 12538 3566 12540
rect 3622 12538 3628 12540
rect 3382 12486 3384 12538
rect 3564 12486 3566 12538
rect 3320 12484 3326 12486
rect 3382 12484 3406 12486
rect 3462 12484 3486 12486
rect 3542 12484 3566 12486
rect 3622 12484 3628 12486
rect 3320 12475 3628 12484
rect 3712 12442 3740 14214
rect 3794 14172 4102 14181
rect 3794 14170 3800 14172
rect 3856 14170 3880 14172
rect 3936 14170 3960 14172
rect 4016 14170 4040 14172
rect 4096 14170 4102 14172
rect 3856 14118 3858 14170
rect 4038 14118 4040 14170
rect 3794 14116 3800 14118
rect 3856 14116 3880 14118
rect 3936 14116 3960 14118
rect 4016 14116 4040 14118
rect 4096 14116 4102 14118
rect 3794 14107 4102 14116
rect 4172 13954 4200 14334
rect 4264 14249 4292 14350
rect 4250 14240 4306 14249
rect 4250 14175 4306 14184
rect 4080 13926 4200 13954
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 13258 4016 13670
rect 4080 13394 4108 13926
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3794 13084 4102 13093
rect 3794 13082 3800 13084
rect 3856 13082 3880 13084
rect 3936 13082 3960 13084
rect 4016 13082 4040 13084
rect 4096 13082 4102 13084
rect 3856 13030 3858 13082
rect 4038 13030 4040 13082
rect 3794 13028 3800 13030
rect 3856 13028 3880 13030
rect 3936 13028 3960 13030
rect 4016 13028 4040 13030
rect 4096 13028 4102 13030
rect 3794 13019 4102 13028
rect 4172 12986 4200 13738
rect 4268 13628 4576 13637
rect 4268 13626 4274 13628
rect 4330 13626 4354 13628
rect 4410 13626 4434 13628
rect 4490 13626 4514 13628
rect 4570 13626 4576 13628
rect 4330 13574 4332 13626
rect 4512 13574 4514 13626
rect 4268 13572 4274 13574
rect 4330 13572 4354 13574
rect 4410 13572 4434 13574
rect 4490 13572 4514 13574
rect 4570 13572 4576 13574
rect 4268 13563 4576 13572
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4066 12744 4122 12753
rect 4066 12679 4122 12688
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3344 11898 3372 12038
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3620 11778 3648 12242
rect 3804 12186 3832 12582
rect 4080 12238 4108 12679
rect 3712 12158 3832 12186
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3712 11898 3740 12158
rect 3794 11996 4102 12005
rect 3794 11994 3800 11996
rect 3856 11994 3880 11996
rect 3936 11994 3960 11996
rect 4016 11994 4040 11996
rect 4096 11994 4102 11996
rect 3856 11942 3858 11994
rect 4038 11942 4040 11994
rect 3794 11940 3800 11942
rect 3856 11940 3880 11942
rect 3936 11940 3960 11942
rect 4016 11940 4040 11942
rect 4096 11940 4102 11942
rect 3794 11931 4102 11940
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3620 11750 3832 11778
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3620 11558 3648 11630
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3252 11234 3280 11494
rect 3320 11452 3628 11461
rect 3320 11450 3326 11452
rect 3382 11450 3406 11452
rect 3462 11450 3486 11452
rect 3542 11450 3566 11452
rect 3622 11450 3628 11452
rect 3382 11398 3384 11450
rect 3564 11398 3566 11450
rect 3320 11396 3326 11398
rect 3382 11396 3406 11398
rect 3462 11396 3486 11398
rect 3542 11396 3566 11398
rect 3622 11396 3628 11398
rect 3320 11387 3628 11396
rect 3424 11280 3476 11286
rect 3422 11248 3424 11257
rect 3476 11248 3478 11257
rect 3252 11206 3372 11234
rect 2792 10962 2820 11086
rect 3160 11070 3280 11098
rect 2700 10934 2820 10962
rect 2700 10742 2728 10934
rect 2846 10908 3154 10917
rect 2846 10906 2852 10908
rect 2908 10906 2932 10908
rect 2988 10906 3012 10908
rect 3068 10906 3092 10908
rect 3148 10906 3154 10908
rect 2908 10854 2910 10906
rect 3090 10854 3092 10906
rect 2846 10852 2852 10854
rect 2908 10852 2932 10854
rect 2988 10852 3012 10854
rect 3068 10852 3092 10854
rect 3148 10852 3154 10854
rect 2846 10843 3154 10852
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2688 10736 2740 10742
rect 2688 10678 2740 10684
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2148 9994 2176 10066
rect 2136 9988 2188 9994
rect 2136 9930 2188 9936
rect 1898 9820 2206 9829
rect 1898 9818 1904 9820
rect 1960 9818 1984 9820
rect 2040 9818 2064 9820
rect 2120 9818 2144 9820
rect 2200 9818 2206 9820
rect 1960 9766 1962 9818
rect 2142 9766 2144 9818
rect 1898 9764 1904 9766
rect 1960 9764 1984 9766
rect 2040 9764 2064 9766
rect 2120 9764 2144 9766
rect 2200 9764 2206 9766
rect 1898 9755 2206 9764
rect 1400 9648 1452 9654
rect 1214 9616 1270 9625
rect 1688 9646 1808 9674
rect 1400 9590 1452 9596
rect 1214 9551 1270 9560
rect 1228 8090 1256 9551
rect 1424 9276 1732 9285
rect 1424 9274 1430 9276
rect 1486 9274 1510 9276
rect 1566 9274 1590 9276
rect 1646 9274 1670 9276
rect 1726 9274 1732 9276
rect 1486 9222 1488 9274
rect 1668 9222 1670 9274
rect 1424 9220 1430 9222
rect 1486 9220 1510 9222
rect 1566 9220 1590 9222
rect 1646 9220 1670 9222
rect 1726 9220 1732 9222
rect 1424 9211 1732 9220
rect 1400 8832 1452 8838
rect 1400 8774 1452 8780
rect 1412 8378 1440 8774
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1320 8350 1440 8378
rect 1688 8378 1716 8570
rect 1780 8514 1808 9646
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1872 8974 1900 9590
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1964 8838 1992 9522
rect 2240 9518 2268 10542
rect 2372 10364 2680 10373
rect 2372 10362 2378 10364
rect 2434 10362 2458 10364
rect 2514 10362 2538 10364
rect 2594 10362 2618 10364
rect 2674 10362 2680 10364
rect 2434 10310 2436 10362
rect 2616 10310 2618 10362
rect 2372 10308 2378 10310
rect 2434 10308 2458 10310
rect 2514 10308 2538 10310
rect 2594 10308 2618 10310
rect 2674 10308 2680 10310
rect 2372 10299 2680 10308
rect 2792 10180 2820 10746
rect 2700 10152 2820 10180
rect 2596 10056 2648 10062
rect 2516 10004 2596 10010
rect 2516 9998 2648 10004
rect 2516 9982 2636 9998
rect 2516 9722 2544 9982
rect 2700 9874 2728 10152
rect 3252 10146 3280 11070
rect 3344 10810 3372 11206
rect 3804 11234 3832 11750
rect 3422 11183 3478 11192
rect 3528 11206 3832 11234
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3528 10577 3556 11206
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3700 11076 3752 11082
rect 3700 11018 3752 11024
rect 3514 10568 3570 10577
rect 3620 10554 3648 11018
rect 3712 10742 3740 11018
rect 3794 10908 4102 10917
rect 3794 10906 3800 10908
rect 3856 10906 3880 10908
rect 3936 10906 3960 10908
rect 4016 10906 4040 10908
rect 4096 10906 4102 10908
rect 3856 10854 3858 10906
rect 4038 10854 4040 10906
rect 3794 10852 3800 10854
rect 3856 10852 3880 10854
rect 3936 10852 3960 10854
rect 4016 10852 4040 10854
rect 4096 10852 4102 10854
rect 3794 10843 4102 10852
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 3620 10526 3740 10554
rect 3514 10503 3570 10512
rect 3320 10364 3628 10373
rect 3320 10362 3326 10364
rect 3382 10362 3406 10364
rect 3462 10362 3486 10364
rect 3542 10362 3566 10364
rect 3622 10362 3628 10364
rect 3382 10310 3384 10362
rect 3564 10310 3566 10362
rect 3320 10308 3326 10310
rect 3382 10308 3406 10310
rect 3462 10308 3486 10310
rect 3542 10308 3566 10310
rect 3622 10308 3628 10310
rect 3320 10299 3628 10308
rect 3606 10160 3662 10169
rect 3252 10118 3372 10146
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 3238 10024 3294 10033
rect 2792 9874 2820 9998
rect 3238 9959 3294 9968
rect 3252 9926 3280 9959
rect 2608 9846 2728 9874
rect 2785 9846 2820 9874
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2608 9674 2636 9846
rect 2785 9704 2813 9846
rect 2846 9820 3154 9829
rect 2846 9818 2852 9820
rect 2908 9818 2932 9820
rect 2988 9818 3012 9820
rect 3068 9818 3092 9820
rect 3148 9818 3154 9820
rect 2908 9766 2910 9818
rect 3090 9766 3092 9818
rect 2846 9764 2852 9766
rect 2908 9764 2932 9766
rect 2988 9764 3012 9766
rect 3068 9764 3092 9766
rect 3148 9764 3154 9766
rect 2846 9755 3154 9764
rect 2785 9676 2820 9704
rect 2608 9646 2728 9674
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2700 9466 2728 9646
rect 2792 9625 2820 9676
rect 2778 9616 2834 9625
rect 3344 9586 3372 10118
rect 3606 10095 3662 10104
rect 2778 9551 2834 9560
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1898 8732 2206 8741
rect 1898 8730 1904 8732
rect 1960 8730 1984 8732
rect 2040 8730 2064 8732
rect 2120 8730 2144 8732
rect 2200 8730 2206 8732
rect 1960 8678 1962 8730
rect 2142 8678 2144 8730
rect 1898 8676 1904 8678
rect 1960 8676 1984 8678
rect 2040 8676 2064 8678
rect 2120 8676 2144 8678
rect 2200 8676 2206 8678
rect 1898 8667 2206 8676
rect 1780 8486 1900 8514
rect 1688 8350 1808 8378
rect 1216 8084 1268 8090
rect 1216 8026 1268 8032
rect 1320 6882 1348 8350
rect 1424 8188 1732 8197
rect 1424 8186 1430 8188
rect 1486 8186 1510 8188
rect 1566 8186 1590 8188
rect 1646 8186 1670 8188
rect 1726 8186 1732 8188
rect 1486 8134 1488 8186
rect 1668 8134 1670 8186
rect 1424 8132 1430 8134
rect 1486 8132 1510 8134
rect 1566 8132 1590 8134
rect 1646 8132 1670 8134
rect 1726 8132 1732 8134
rect 1424 8123 1732 8132
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7449 1440 7822
rect 1398 7440 1454 7449
rect 1398 7375 1454 7384
rect 1424 7100 1732 7109
rect 1424 7098 1430 7100
rect 1486 7098 1510 7100
rect 1566 7098 1590 7100
rect 1646 7098 1670 7100
rect 1726 7098 1732 7100
rect 1486 7046 1488 7098
rect 1668 7046 1670 7098
rect 1424 7044 1430 7046
rect 1486 7044 1510 7046
rect 1566 7044 1590 7046
rect 1646 7044 1670 7046
rect 1726 7044 1732 7046
rect 1424 7035 1732 7044
rect 1320 6854 1440 6882
rect 1412 6202 1440 6854
rect 1780 6458 1808 8350
rect 1872 7886 1900 8486
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1898 7644 2206 7653
rect 1898 7642 1904 7644
rect 1960 7642 1984 7644
rect 2040 7642 2064 7644
rect 2120 7642 2144 7644
rect 2200 7642 2206 7644
rect 1960 7590 1962 7642
rect 2142 7590 2144 7642
rect 1898 7588 1904 7590
rect 1960 7588 1984 7590
rect 2040 7588 2064 7590
rect 2120 7588 2144 7590
rect 2200 7588 2206 7590
rect 1898 7579 2206 7588
rect 1898 6556 2206 6565
rect 1898 6554 1904 6556
rect 1960 6554 1984 6556
rect 2040 6554 2064 6556
rect 2120 6554 2144 6556
rect 2200 6554 2206 6556
rect 1960 6502 1962 6554
rect 2142 6502 2144 6554
rect 1898 6500 1904 6502
rect 1960 6500 1984 6502
rect 2040 6500 2064 6502
rect 2120 6500 2144 6502
rect 2200 6500 2206 6502
rect 1898 6491 2206 6500
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1320 6174 1440 6202
rect 1320 5794 1348 6174
rect 1424 6012 1732 6021
rect 1424 6010 1430 6012
rect 1486 6010 1510 6012
rect 1566 6010 1590 6012
rect 1646 6010 1670 6012
rect 1726 6010 1732 6012
rect 1486 5958 1488 6010
rect 1668 5958 1670 6010
rect 1424 5956 1430 5958
rect 1486 5956 1510 5958
rect 1566 5956 1590 5958
rect 1646 5956 1670 5958
rect 1726 5956 1732 5958
rect 1424 5947 1732 5956
rect 1320 5766 1440 5794
rect 1412 5114 1440 5766
rect 1320 5086 1440 5114
rect 1320 4826 1348 5086
rect 1424 4924 1732 4933
rect 1424 4922 1430 4924
rect 1486 4922 1510 4924
rect 1566 4922 1590 4924
rect 1646 4922 1670 4924
rect 1726 4922 1732 4924
rect 1486 4870 1488 4922
rect 1668 4870 1670 4922
rect 1424 4868 1430 4870
rect 1486 4868 1510 4870
rect 1566 4868 1590 4870
rect 1646 4868 1670 4870
rect 1726 4868 1732 4870
rect 1424 4859 1732 4868
rect 1308 4820 1360 4826
rect 1308 4762 1360 4768
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1412 4457 1440 4558
rect 1398 4448 1454 4457
rect 1398 4383 1454 4392
rect 1424 3836 1732 3845
rect 1424 3834 1430 3836
rect 1486 3834 1510 3836
rect 1566 3834 1590 3836
rect 1646 3834 1670 3836
rect 1726 3834 1732 3836
rect 1486 3782 1488 3834
rect 1668 3782 1670 3834
rect 1424 3780 1430 3782
rect 1486 3780 1510 3782
rect 1566 3780 1590 3782
rect 1646 3780 1670 3782
rect 1726 3780 1732 3782
rect 1424 3771 1732 3780
rect 1424 2748 1732 2757
rect 1424 2746 1430 2748
rect 1486 2746 1510 2748
rect 1566 2746 1590 2748
rect 1646 2746 1670 2748
rect 1726 2746 1732 2748
rect 1486 2694 1488 2746
rect 1668 2694 1670 2746
rect 1424 2692 1430 2694
rect 1486 2692 1510 2694
rect 1566 2692 1590 2694
rect 1646 2692 1670 2694
rect 1726 2692 1732 2694
rect 1424 2683 1732 2692
rect 1424 1660 1732 1669
rect 1424 1658 1430 1660
rect 1486 1658 1510 1660
rect 1566 1658 1590 1660
rect 1646 1658 1670 1660
rect 1726 1658 1732 1660
rect 1486 1606 1488 1658
rect 1668 1606 1670 1658
rect 1424 1604 1430 1606
rect 1486 1604 1510 1606
rect 1566 1604 1590 1606
rect 1646 1604 1670 1606
rect 1726 1604 1732 1606
rect 1424 1595 1732 1604
rect 1780 1465 1808 6258
rect 2148 5658 2176 6394
rect 2240 6390 2268 9454
rect 2700 9438 2820 9466
rect 2372 9276 2680 9285
rect 2372 9274 2378 9276
rect 2434 9274 2458 9276
rect 2514 9274 2538 9276
rect 2594 9274 2618 9276
rect 2674 9274 2680 9276
rect 2434 9222 2436 9274
rect 2616 9222 2618 9274
rect 2372 9220 2378 9222
rect 2434 9220 2458 9222
rect 2514 9220 2538 9222
rect 2594 9220 2618 9222
rect 2674 9220 2680 9222
rect 2372 9211 2680 9220
rect 2792 9058 2820 9438
rect 3620 9382 3648 10095
rect 3712 9926 3740 10526
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3320 9276 3628 9285
rect 3320 9274 3326 9276
rect 3382 9274 3406 9276
rect 3462 9274 3486 9276
rect 3542 9274 3566 9276
rect 3622 9274 3628 9276
rect 3382 9222 3384 9274
rect 3564 9222 3566 9274
rect 3320 9220 3326 9222
rect 3382 9220 3406 9222
rect 3462 9220 3486 9222
rect 3542 9220 3566 9222
rect 3622 9220 3628 9222
rect 3320 9211 3628 9220
rect 3712 9178 3740 9862
rect 3794 9820 4102 9829
rect 3794 9818 3800 9820
rect 3856 9818 3880 9820
rect 3936 9818 3960 9820
rect 4016 9818 4040 9820
rect 4096 9818 4102 9820
rect 3856 9766 3858 9818
rect 4038 9766 4040 9818
rect 3794 9764 3800 9766
rect 3856 9764 3880 9766
rect 3936 9764 3960 9766
rect 4016 9764 4040 9766
rect 4096 9764 4102 9766
rect 3794 9755 4102 9764
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 2700 9030 2820 9058
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 2700 8498 2728 9030
rect 2846 8732 3154 8741
rect 2846 8730 2852 8732
rect 2908 8730 2932 8732
rect 2988 8730 3012 8732
rect 3068 8730 3092 8732
rect 3148 8730 3154 8732
rect 2908 8678 2910 8730
rect 3090 8678 3092 8730
rect 2846 8676 2852 8678
rect 2908 8676 2932 8678
rect 2988 8676 3012 8678
rect 3068 8676 3092 8678
rect 3148 8676 3154 8678
rect 2846 8667 3154 8676
rect 3252 8566 3280 9046
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2372 8188 2680 8197
rect 2372 8186 2378 8188
rect 2434 8186 2458 8188
rect 2514 8186 2538 8188
rect 2594 8186 2618 8188
rect 2674 8186 2680 8188
rect 2434 8134 2436 8186
rect 2616 8134 2618 8186
rect 2372 8132 2378 8134
rect 2434 8132 2458 8134
rect 2514 8132 2538 8134
rect 2594 8132 2618 8134
rect 2674 8132 2680 8134
rect 2372 8123 2680 8132
rect 3252 8090 3280 8502
rect 3344 8498 3372 9114
rect 3712 8974 3740 9114
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3320 8188 3628 8197
rect 3320 8186 3326 8188
rect 3382 8186 3406 8188
rect 3462 8186 3486 8188
rect 3542 8186 3566 8188
rect 3622 8186 3628 8188
rect 3382 8134 3384 8186
rect 3564 8134 3566 8186
rect 3320 8132 3326 8134
rect 3382 8132 3406 8134
rect 3462 8132 3486 8134
rect 3542 8132 3566 8134
rect 3622 8132 3628 8134
rect 3320 8123 3628 8132
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3252 7834 3280 8026
rect 3252 7806 3372 7834
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 2846 7644 3154 7653
rect 2846 7642 2852 7644
rect 2908 7642 2932 7644
rect 2988 7642 3012 7644
rect 3068 7642 3092 7644
rect 3148 7642 3154 7644
rect 2908 7590 2910 7642
rect 3090 7590 3092 7642
rect 2846 7588 2852 7590
rect 2908 7588 2932 7590
rect 2988 7588 3012 7590
rect 3068 7588 3092 7590
rect 3148 7588 3154 7590
rect 2846 7579 3154 7588
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2372 7100 2680 7109
rect 2372 7098 2378 7100
rect 2434 7098 2458 7100
rect 2514 7098 2538 7100
rect 2594 7098 2618 7100
rect 2674 7098 2680 7100
rect 2434 7046 2436 7098
rect 2616 7046 2618 7098
rect 2372 7044 2378 7046
rect 2434 7044 2458 7046
rect 2514 7044 2538 7046
rect 2594 7044 2618 7046
rect 2674 7044 2680 7046
rect 2372 7035 2680 7044
rect 3160 6662 3188 7346
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2846 6556 3154 6565
rect 2846 6554 2852 6556
rect 2908 6554 2932 6556
rect 2988 6554 3012 6556
rect 3068 6554 3092 6556
rect 3148 6554 3154 6556
rect 2908 6502 2910 6554
rect 3090 6502 3092 6554
rect 2846 6500 2852 6502
rect 2908 6500 2932 6502
rect 2988 6500 3012 6502
rect 3068 6500 3092 6502
rect 3148 6500 3154 6502
rect 2846 6491 3154 6500
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 2372 6012 2680 6021
rect 2372 6010 2378 6012
rect 2434 6010 2458 6012
rect 2514 6010 2538 6012
rect 2594 6010 2618 6012
rect 2674 6010 2680 6012
rect 2434 5958 2436 6010
rect 2616 5958 2618 6010
rect 2372 5956 2378 5958
rect 2434 5956 2458 5958
rect 2514 5956 2538 5958
rect 2594 5956 2618 5958
rect 2674 5956 2680 5958
rect 2372 5947 2680 5956
rect 2148 5630 2268 5658
rect 1898 5468 2206 5477
rect 1898 5466 1904 5468
rect 1960 5466 1984 5468
rect 2040 5466 2064 5468
rect 2120 5466 2144 5468
rect 2200 5466 2206 5468
rect 1960 5414 1962 5466
rect 2142 5414 2144 5466
rect 1898 5412 1904 5414
rect 1960 5412 1984 5414
rect 2040 5412 2064 5414
rect 2120 5412 2144 5414
rect 2200 5412 2206 5414
rect 1898 5403 2206 5412
rect 1898 4380 2206 4389
rect 1898 4378 1904 4380
rect 1960 4378 1984 4380
rect 2040 4378 2064 4380
rect 2120 4378 2144 4380
rect 2200 4378 2206 4380
rect 1960 4326 1962 4378
rect 2142 4326 2144 4378
rect 1898 4324 1904 4326
rect 1960 4324 1984 4326
rect 2040 4324 2064 4326
rect 2120 4324 2144 4326
rect 2200 4324 2206 4326
rect 1898 4315 2206 4324
rect 1898 3292 2206 3301
rect 1898 3290 1904 3292
rect 1960 3290 1984 3292
rect 2040 3290 2064 3292
rect 2120 3290 2144 3292
rect 2200 3290 2206 3292
rect 1960 3238 1962 3290
rect 2142 3238 2144 3290
rect 1898 3236 1904 3238
rect 1960 3236 1984 3238
rect 2040 3236 2064 3238
rect 2120 3236 2144 3238
rect 2200 3236 2206 3238
rect 1898 3227 2206 3236
rect 2240 2417 2268 5630
rect 2846 5468 3154 5477
rect 2846 5466 2852 5468
rect 2908 5466 2932 5468
rect 2988 5466 3012 5468
rect 3068 5466 3092 5468
rect 3148 5466 3154 5468
rect 2908 5414 2910 5466
rect 3090 5414 3092 5466
rect 2846 5412 2852 5414
rect 2908 5412 2932 5414
rect 2988 5412 3012 5414
rect 3068 5412 3092 5414
rect 3148 5412 3154 5414
rect 2846 5403 3154 5412
rect 2372 4924 2680 4933
rect 2372 4922 2378 4924
rect 2434 4922 2458 4924
rect 2514 4922 2538 4924
rect 2594 4922 2618 4924
rect 2674 4922 2680 4924
rect 2434 4870 2436 4922
rect 2616 4870 2618 4922
rect 2372 4868 2378 4870
rect 2434 4868 2458 4870
rect 2514 4868 2538 4870
rect 2594 4868 2618 4870
rect 2674 4868 2680 4870
rect 2372 4859 2680 4868
rect 2846 4380 3154 4389
rect 2846 4378 2852 4380
rect 2908 4378 2932 4380
rect 2988 4378 3012 4380
rect 3068 4378 3092 4380
rect 3148 4378 3154 4380
rect 2908 4326 2910 4378
rect 3090 4326 3092 4378
rect 2846 4324 2852 4326
rect 2908 4324 2932 4326
rect 2988 4324 3012 4326
rect 3068 4324 3092 4326
rect 3148 4324 3154 4326
rect 2846 4315 3154 4324
rect 3252 4049 3280 7686
rect 3344 7410 3372 7806
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3320 7100 3628 7109
rect 3320 7098 3326 7100
rect 3382 7098 3406 7100
rect 3462 7098 3486 7100
rect 3542 7098 3566 7100
rect 3622 7098 3628 7100
rect 3382 7046 3384 7098
rect 3564 7046 3566 7098
rect 3320 7044 3326 7046
rect 3382 7044 3406 7046
rect 3462 7044 3486 7046
rect 3542 7044 3566 7046
rect 3622 7044 3628 7046
rect 3320 7035 3628 7044
rect 3712 6769 3740 8774
rect 3794 8732 4102 8741
rect 3794 8730 3800 8732
rect 3856 8730 3880 8732
rect 3936 8730 3960 8732
rect 4016 8730 4040 8732
rect 4096 8730 4102 8732
rect 3856 8678 3858 8730
rect 4038 8678 4040 8730
rect 3794 8676 3800 8678
rect 3856 8676 3880 8678
rect 3936 8676 3960 8678
rect 4016 8676 4040 8678
rect 4096 8676 4102 8678
rect 3794 8667 4102 8676
rect 3794 7644 4102 7653
rect 3794 7642 3800 7644
rect 3856 7642 3880 7644
rect 3936 7642 3960 7644
rect 4016 7642 4040 7644
rect 4096 7642 4102 7644
rect 3856 7590 3858 7642
rect 4038 7590 4040 7642
rect 3794 7588 3800 7590
rect 3856 7588 3880 7590
rect 3936 7588 3960 7590
rect 4016 7588 4040 7590
rect 4096 7588 4102 7590
rect 3794 7579 4102 7588
rect 4172 7410 4200 12922
rect 4540 12730 4568 13126
rect 4632 12832 4660 15982
rect 4710 15736 4766 15745
rect 4710 15671 4766 15680
rect 4724 15502 4752 15671
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4724 13190 4752 14758
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4632 12804 4752 12832
rect 4540 12702 4660 12730
rect 4268 12540 4576 12549
rect 4268 12538 4274 12540
rect 4330 12538 4354 12540
rect 4410 12538 4434 12540
rect 4490 12538 4514 12540
rect 4570 12538 4576 12540
rect 4330 12486 4332 12538
rect 4512 12486 4514 12538
rect 4268 12484 4274 12486
rect 4330 12484 4354 12486
rect 4410 12484 4434 12486
rect 4490 12484 4514 12486
rect 4570 12484 4576 12486
rect 4268 12475 4576 12484
rect 4268 11452 4576 11461
rect 4268 11450 4274 11452
rect 4330 11450 4354 11452
rect 4410 11450 4434 11452
rect 4490 11450 4514 11452
rect 4570 11450 4576 11452
rect 4330 11398 4332 11450
rect 4512 11398 4514 11450
rect 4268 11396 4274 11398
rect 4330 11396 4354 11398
rect 4410 11396 4434 11398
rect 4490 11396 4514 11398
rect 4570 11396 4576 11398
rect 4268 11387 4576 11396
rect 4268 10364 4576 10373
rect 4268 10362 4274 10364
rect 4330 10362 4354 10364
rect 4410 10362 4434 10364
rect 4490 10362 4514 10364
rect 4570 10362 4576 10364
rect 4330 10310 4332 10362
rect 4512 10310 4514 10362
rect 4268 10308 4274 10310
rect 4330 10308 4354 10310
rect 4410 10308 4434 10310
rect 4490 10308 4514 10310
rect 4570 10308 4576 10310
rect 4268 10299 4576 10308
rect 4268 9276 4576 9285
rect 4268 9274 4274 9276
rect 4330 9274 4354 9276
rect 4410 9274 4434 9276
rect 4490 9274 4514 9276
rect 4570 9274 4576 9276
rect 4330 9222 4332 9274
rect 4512 9222 4514 9274
rect 4268 9220 4274 9222
rect 4330 9220 4354 9222
rect 4410 9220 4434 9222
rect 4490 9220 4514 9222
rect 4570 9220 4576 9222
rect 4268 9211 4576 9220
rect 4632 8498 4660 12702
rect 4724 12170 4752 12804
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4724 10130 4752 12106
rect 4816 10810 4844 17070
rect 4908 13530 4936 19654
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4724 8265 4752 8298
rect 4710 8256 4766 8265
rect 4268 8188 4576 8197
rect 4710 8191 4766 8200
rect 4268 8186 4274 8188
rect 4330 8186 4354 8188
rect 4410 8186 4434 8188
rect 4490 8186 4514 8188
rect 4570 8186 4576 8188
rect 4330 8134 4332 8186
rect 4512 8134 4514 8186
rect 4268 8132 4274 8134
rect 4330 8132 4354 8134
rect 4410 8132 4434 8134
rect 4490 8132 4514 8134
rect 4570 8132 4576 8134
rect 4268 8123 4576 8132
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 3698 6760 3754 6769
rect 3698 6695 3754 6704
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3344 6322 3372 6598
rect 3794 6556 4102 6565
rect 3794 6554 3800 6556
rect 3856 6554 3880 6556
rect 3936 6554 3960 6556
rect 4016 6554 4040 6556
rect 4096 6554 4102 6556
rect 3856 6502 3858 6554
rect 4038 6502 4040 6554
rect 3794 6500 3800 6502
rect 3856 6500 3880 6502
rect 3936 6500 3960 6502
rect 4016 6500 4040 6502
rect 4096 6500 4102 6502
rect 3794 6491 4102 6500
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3320 6012 3628 6021
rect 3320 6010 3326 6012
rect 3382 6010 3406 6012
rect 3462 6010 3486 6012
rect 3542 6010 3566 6012
rect 3622 6010 3628 6012
rect 3382 5958 3384 6010
rect 3564 5958 3566 6010
rect 3320 5956 3326 5958
rect 3382 5956 3406 5958
rect 3462 5956 3486 5958
rect 3542 5956 3566 5958
rect 3622 5956 3628 5958
rect 3320 5947 3628 5956
rect 3794 5468 4102 5477
rect 3794 5466 3800 5468
rect 3856 5466 3880 5468
rect 3936 5466 3960 5468
rect 4016 5466 4040 5468
rect 4096 5466 4102 5468
rect 3856 5414 3858 5466
rect 4038 5414 4040 5466
rect 3794 5412 3800 5414
rect 3856 5412 3880 5414
rect 3936 5412 3960 5414
rect 4016 5412 4040 5414
rect 4096 5412 4102 5414
rect 3794 5403 4102 5412
rect 4172 5273 4200 7142
rect 4268 7100 4576 7109
rect 4268 7098 4274 7100
rect 4330 7098 4354 7100
rect 4410 7098 4434 7100
rect 4490 7098 4514 7100
rect 4570 7098 4576 7100
rect 4330 7046 4332 7098
rect 4512 7046 4514 7098
rect 4268 7044 4274 7046
rect 4330 7044 4354 7046
rect 4410 7044 4434 7046
rect 4490 7044 4514 7046
rect 4570 7044 4576 7046
rect 4268 7035 4576 7044
rect 4816 6322 4844 9318
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4268 6012 4576 6021
rect 4268 6010 4274 6012
rect 4330 6010 4354 6012
rect 4410 6010 4434 6012
rect 4490 6010 4514 6012
rect 4570 6010 4576 6012
rect 4330 5958 4332 6010
rect 4512 5958 4514 6010
rect 4268 5956 4274 5958
rect 4330 5956 4354 5958
rect 4410 5956 4434 5958
rect 4490 5956 4514 5958
rect 4570 5956 4576 5958
rect 4268 5947 4576 5956
rect 4158 5264 4214 5273
rect 4158 5199 4214 5208
rect 3320 4924 3628 4933
rect 3320 4922 3326 4924
rect 3382 4922 3406 4924
rect 3462 4922 3486 4924
rect 3542 4922 3566 4924
rect 3622 4922 3628 4924
rect 3382 4870 3384 4922
rect 3564 4870 3566 4922
rect 3320 4868 3326 4870
rect 3382 4868 3406 4870
rect 3462 4868 3486 4870
rect 3542 4868 3566 4870
rect 3622 4868 3628 4870
rect 3320 4859 3628 4868
rect 4268 4924 4576 4933
rect 4268 4922 4274 4924
rect 4330 4922 4354 4924
rect 4410 4922 4434 4924
rect 4490 4922 4514 4924
rect 4570 4922 4576 4924
rect 4330 4870 4332 4922
rect 4512 4870 4514 4922
rect 4268 4868 4274 4870
rect 4330 4868 4354 4870
rect 4410 4868 4434 4870
rect 4490 4868 4514 4870
rect 4570 4868 4576 4870
rect 4268 4859 4576 4868
rect 3794 4380 4102 4389
rect 3794 4378 3800 4380
rect 3856 4378 3880 4380
rect 3936 4378 3960 4380
rect 4016 4378 4040 4380
rect 4096 4378 4102 4380
rect 3856 4326 3858 4378
rect 4038 4326 4040 4378
rect 3794 4324 3800 4326
rect 3856 4324 3880 4326
rect 3936 4324 3960 4326
rect 4016 4324 4040 4326
rect 4096 4324 4102 4326
rect 3794 4315 4102 4324
rect 3238 4040 3294 4049
rect 3238 3975 3294 3984
rect 2372 3836 2680 3845
rect 2372 3834 2378 3836
rect 2434 3834 2458 3836
rect 2514 3834 2538 3836
rect 2594 3834 2618 3836
rect 2674 3834 2680 3836
rect 2434 3782 2436 3834
rect 2616 3782 2618 3834
rect 2372 3780 2378 3782
rect 2434 3780 2458 3782
rect 2514 3780 2538 3782
rect 2594 3780 2618 3782
rect 2674 3780 2680 3782
rect 2372 3771 2680 3780
rect 3320 3836 3628 3845
rect 3320 3834 3326 3836
rect 3382 3834 3406 3836
rect 3462 3834 3486 3836
rect 3542 3834 3566 3836
rect 3622 3834 3628 3836
rect 3382 3782 3384 3834
rect 3564 3782 3566 3834
rect 3320 3780 3326 3782
rect 3382 3780 3406 3782
rect 3462 3780 3486 3782
rect 3542 3780 3566 3782
rect 3622 3780 3628 3782
rect 3320 3771 3628 3780
rect 4268 3836 4576 3845
rect 4268 3834 4274 3836
rect 4330 3834 4354 3836
rect 4410 3834 4434 3836
rect 4490 3834 4514 3836
rect 4570 3834 4576 3836
rect 4330 3782 4332 3834
rect 4512 3782 4514 3834
rect 4268 3780 4274 3782
rect 4330 3780 4354 3782
rect 4410 3780 4434 3782
rect 4490 3780 4514 3782
rect 4570 3780 4576 3782
rect 4268 3771 4576 3780
rect 2846 3292 3154 3301
rect 2846 3290 2852 3292
rect 2908 3290 2932 3292
rect 2988 3290 3012 3292
rect 3068 3290 3092 3292
rect 3148 3290 3154 3292
rect 2908 3238 2910 3290
rect 3090 3238 3092 3290
rect 2846 3236 2852 3238
rect 2908 3236 2932 3238
rect 2988 3236 3012 3238
rect 3068 3236 3092 3238
rect 3148 3236 3154 3238
rect 2846 3227 3154 3236
rect 3794 3292 4102 3301
rect 3794 3290 3800 3292
rect 3856 3290 3880 3292
rect 3936 3290 3960 3292
rect 4016 3290 4040 3292
rect 4096 3290 4102 3292
rect 3856 3238 3858 3290
rect 4038 3238 4040 3290
rect 3794 3236 3800 3238
rect 3856 3236 3880 3238
rect 3936 3236 3960 3238
rect 4016 3236 4040 3238
rect 4096 3236 4102 3238
rect 3794 3227 4102 3236
rect 2372 2748 2680 2757
rect 2372 2746 2378 2748
rect 2434 2746 2458 2748
rect 2514 2746 2538 2748
rect 2594 2746 2618 2748
rect 2674 2746 2680 2748
rect 2434 2694 2436 2746
rect 2616 2694 2618 2746
rect 2372 2692 2378 2694
rect 2434 2692 2458 2694
rect 2514 2692 2538 2694
rect 2594 2692 2618 2694
rect 2674 2692 2680 2694
rect 2372 2683 2680 2692
rect 3320 2748 3628 2757
rect 3320 2746 3326 2748
rect 3382 2746 3406 2748
rect 3462 2746 3486 2748
rect 3542 2746 3566 2748
rect 3622 2746 3628 2748
rect 3382 2694 3384 2746
rect 3564 2694 3566 2746
rect 3320 2692 3326 2694
rect 3382 2692 3406 2694
rect 3462 2692 3486 2694
rect 3542 2692 3566 2694
rect 3622 2692 3628 2694
rect 3320 2683 3628 2692
rect 4268 2748 4576 2757
rect 4268 2746 4274 2748
rect 4330 2746 4354 2748
rect 4410 2746 4434 2748
rect 4490 2746 4514 2748
rect 4570 2746 4576 2748
rect 4330 2694 4332 2746
rect 4512 2694 4514 2746
rect 4268 2692 4274 2694
rect 4330 2692 4354 2694
rect 4410 2692 4434 2694
rect 4490 2692 4514 2694
rect 4570 2692 4576 2694
rect 4268 2683 4576 2692
rect 2226 2408 2282 2417
rect 2226 2343 2282 2352
rect 1898 2204 2206 2213
rect 1898 2202 1904 2204
rect 1960 2202 1984 2204
rect 2040 2202 2064 2204
rect 2120 2202 2144 2204
rect 2200 2202 2206 2204
rect 1960 2150 1962 2202
rect 2142 2150 2144 2202
rect 1898 2148 1904 2150
rect 1960 2148 1984 2150
rect 2040 2148 2064 2150
rect 2120 2148 2144 2150
rect 2200 2148 2206 2150
rect 1898 2139 2206 2148
rect 2846 2204 3154 2213
rect 2846 2202 2852 2204
rect 2908 2202 2932 2204
rect 2988 2202 3012 2204
rect 3068 2202 3092 2204
rect 3148 2202 3154 2204
rect 2908 2150 2910 2202
rect 3090 2150 3092 2202
rect 2846 2148 2852 2150
rect 2908 2148 2932 2150
rect 2988 2148 3012 2150
rect 3068 2148 3092 2150
rect 3148 2148 3154 2150
rect 2846 2139 3154 2148
rect 3794 2204 4102 2213
rect 3794 2202 3800 2204
rect 3856 2202 3880 2204
rect 3936 2202 3960 2204
rect 4016 2202 4040 2204
rect 4096 2202 4102 2204
rect 3856 2150 3858 2202
rect 4038 2150 4040 2202
rect 3794 2148 3800 2150
rect 3856 2148 3880 2150
rect 3936 2148 3960 2150
rect 4016 2148 4040 2150
rect 4096 2148 4102 2150
rect 3794 2139 4102 2148
rect 2372 1660 2680 1669
rect 2372 1658 2378 1660
rect 2434 1658 2458 1660
rect 2514 1658 2538 1660
rect 2594 1658 2618 1660
rect 2674 1658 2680 1660
rect 2434 1606 2436 1658
rect 2616 1606 2618 1658
rect 2372 1604 2378 1606
rect 2434 1604 2458 1606
rect 2514 1604 2538 1606
rect 2594 1604 2618 1606
rect 2674 1604 2680 1606
rect 2372 1595 2680 1604
rect 3320 1660 3628 1669
rect 3320 1658 3326 1660
rect 3382 1658 3406 1660
rect 3462 1658 3486 1660
rect 3542 1658 3566 1660
rect 3622 1658 3628 1660
rect 3382 1606 3384 1658
rect 3564 1606 3566 1658
rect 3320 1604 3326 1606
rect 3382 1604 3406 1606
rect 3462 1604 3486 1606
rect 3542 1604 3566 1606
rect 3622 1604 3628 1606
rect 3320 1595 3628 1604
rect 4268 1660 4576 1669
rect 4268 1658 4274 1660
rect 4330 1658 4354 1660
rect 4410 1658 4434 1660
rect 4490 1658 4514 1660
rect 4570 1658 4576 1660
rect 4330 1606 4332 1658
rect 4512 1606 4514 1658
rect 4268 1604 4274 1606
rect 4330 1604 4354 1606
rect 4410 1604 4434 1606
rect 4490 1604 4514 1606
rect 4570 1604 4576 1606
rect 4268 1595 4576 1604
rect 1766 1456 1822 1465
rect 1766 1391 1822 1400
rect 1898 1116 2206 1125
rect 1898 1114 1904 1116
rect 1960 1114 1984 1116
rect 2040 1114 2064 1116
rect 2120 1114 2144 1116
rect 2200 1114 2206 1116
rect 1960 1062 1962 1114
rect 2142 1062 2144 1114
rect 1898 1060 1904 1062
rect 1960 1060 1984 1062
rect 2040 1060 2064 1062
rect 2120 1060 2144 1062
rect 2200 1060 2206 1062
rect 1898 1051 2206 1060
rect 2846 1116 3154 1125
rect 2846 1114 2852 1116
rect 2908 1114 2932 1116
rect 2988 1114 3012 1116
rect 3068 1114 3092 1116
rect 3148 1114 3154 1116
rect 2908 1062 2910 1114
rect 3090 1062 3092 1114
rect 2846 1060 2852 1062
rect 2908 1060 2932 1062
rect 2988 1060 3012 1062
rect 3068 1060 3092 1062
rect 3148 1060 3154 1062
rect 2846 1051 3154 1060
rect 3794 1116 4102 1125
rect 3794 1114 3800 1116
rect 3856 1114 3880 1116
rect 3936 1114 3960 1116
rect 4016 1114 4040 1116
rect 4096 1114 4102 1116
rect 3856 1062 3858 1114
rect 4038 1062 4040 1114
rect 3794 1060 3800 1062
rect 3856 1060 3880 1062
rect 3936 1060 3960 1062
rect 4016 1060 4040 1062
rect 4096 1060 4102 1062
rect 3794 1051 4102 1060
rect 4724 785 4752 6054
rect 4710 776 4766 785
rect 4710 711 4766 720
<< via2 >>
rect 4158 23160 4214 23216
rect 1904 22874 1960 22876
rect 1984 22874 2040 22876
rect 2064 22874 2120 22876
rect 2144 22874 2200 22876
rect 1904 22822 1950 22874
rect 1950 22822 1960 22874
rect 1984 22822 2014 22874
rect 2014 22822 2026 22874
rect 2026 22822 2040 22874
rect 2064 22822 2078 22874
rect 2078 22822 2090 22874
rect 2090 22822 2120 22874
rect 2144 22822 2154 22874
rect 2154 22822 2200 22874
rect 1904 22820 1960 22822
rect 1984 22820 2040 22822
rect 2064 22820 2120 22822
rect 2144 22820 2200 22822
rect 2852 22874 2908 22876
rect 2932 22874 2988 22876
rect 3012 22874 3068 22876
rect 3092 22874 3148 22876
rect 2852 22822 2898 22874
rect 2898 22822 2908 22874
rect 2932 22822 2962 22874
rect 2962 22822 2974 22874
rect 2974 22822 2988 22874
rect 3012 22822 3026 22874
rect 3026 22822 3038 22874
rect 3038 22822 3068 22874
rect 3092 22822 3102 22874
rect 3102 22822 3148 22874
rect 2852 22820 2908 22822
rect 2932 22820 2988 22822
rect 3012 22820 3068 22822
rect 3092 22820 3148 22822
rect 3800 22874 3856 22876
rect 3880 22874 3936 22876
rect 3960 22874 4016 22876
rect 4040 22874 4096 22876
rect 3800 22822 3846 22874
rect 3846 22822 3856 22874
rect 3880 22822 3910 22874
rect 3910 22822 3922 22874
rect 3922 22822 3936 22874
rect 3960 22822 3974 22874
rect 3974 22822 3986 22874
rect 3986 22822 4016 22874
rect 4040 22822 4050 22874
rect 4050 22822 4096 22874
rect 3800 22820 3856 22822
rect 3880 22820 3936 22822
rect 3960 22820 4016 22822
rect 4040 22820 4096 22822
rect 1430 22330 1486 22332
rect 1510 22330 1566 22332
rect 1590 22330 1646 22332
rect 1670 22330 1726 22332
rect 1430 22278 1476 22330
rect 1476 22278 1486 22330
rect 1510 22278 1540 22330
rect 1540 22278 1552 22330
rect 1552 22278 1566 22330
rect 1590 22278 1604 22330
rect 1604 22278 1616 22330
rect 1616 22278 1646 22330
rect 1670 22278 1680 22330
rect 1680 22278 1726 22330
rect 1430 22276 1486 22278
rect 1510 22276 1566 22278
rect 1590 22276 1646 22278
rect 1670 22276 1726 22278
rect 2378 22330 2434 22332
rect 2458 22330 2514 22332
rect 2538 22330 2594 22332
rect 2618 22330 2674 22332
rect 2378 22278 2424 22330
rect 2424 22278 2434 22330
rect 2458 22278 2488 22330
rect 2488 22278 2500 22330
rect 2500 22278 2514 22330
rect 2538 22278 2552 22330
rect 2552 22278 2564 22330
rect 2564 22278 2594 22330
rect 2618 22278 2628 22330
rect 2628 22278 2674 22330
rect 2378 22276 2434 22278
rect 2458 22276 2514 22278
rect 2538 22276 2594 22278
rect 2618 22276 2674 22278
rect 1766 22072 1822 22128
rect 1430 21242 1486 21244
rect 1510 21242 1566 21244
rect 1590 21242 1646 21244
rect 1670 21242 1726 21244
rect 1430 21190 1476 21242
rect 1476 21190 1486 21242
rect 1510 21190 1540 21242
rect 1540 21190 1552 21242
rect 1552 21190 1566 21242
rect 1590 21190 1604 21242
rect 1604 21190 1616 21242
rect 1616 21190 1646 21242
rect 1670 21190 1680 21242
rect 1680 21190 1726 21242
rect 1430 21188 1486 21190
rect 1510 21188 1566 21190
rect 1590 21188 1646 21190
rect 1670 21188 1726 21190
rect 1430 20154 1486 20156
rect 1510 20154 1566 20156
rect 1590 20154 1646 20156
rect 1670 20154 1726 20156
rect 1430 20102 1476 20154
rect 1476 20102 1486 20154
rect 1510 20102 1540 20154
rect 1540 20102 1552 20154
rect 1552 20102 1566 20154
rect 1590 20102 1604 20154
rect 1604 20102 1616 20154
rect 1616 20102 1646 20154
rect 1670 20102 1680 20154
rect 1680 20102 1726 20154
rect 1430 20100 1486 20102
rect 1510 20100 1566 20102
rect 1590 20100 1646 20102
rect 1670 20100 1726 20102
rect 1430 19066 1486 19068
rect 1510 19066 1566 19068
rect 1590 19066 1646 19068
rect 1670 19066 1726 19068
rect 1430 19014 1476 19066
rect 1476 19014 1486 19066
rect 1510 19014 1540 19066
rect 1540 19014 1552 19066
rect 1552 19014 1566 19066
rect 1590 19014 1604 19066
rect 1604 19014 1616 19066
rect 1616 19014 1646 19066
rect 1670 19014 1680 19066
rect 1680 19014 1726 19066
rect 1430 19012 1486 19014
rect 1510 19012 1566 19014
rect 1590 19012 1646 19014
rect 1670 19012 1726 19014
rect 1430 17978 1486 17980
rect 1510 17978 1566 17980
rect 1590 17978 1646 17980
rect 1670 17978 1726 17980
rect 1430 17926 1476 17978
rect 1476 17926 1486 17978
rect 1510 17926 1540 17978
rect 1540 17926 1552 17978
rect 1552 17926 1566 17978
rect 1590 17926 1604 17978
rect 1604 17926 1616 17978
rect 1616 17926 1646 17978
rect 1670 17926 1680 17978
rect 1680 17926 1726 17978
rect 1430 17924 1486 17926
rect 1510 17924 1566 17926
rect 1590 17924 1646 17926
rect 1670 17924 1726 17926
rect 3326 22330 3382 22332
rect 3406 22330 3462 22332
rect 3486 22330 3542 22332
rect 3566 22330 3622 22332
rect 3326 22278 3372 22330
rect 3372 22278 3382 22330
rect 3406 22278 3436 22330
rect 3436 22278 3448 22330
rect 3448 22278 3462 22330
rect 3486 22278 3500 22330
rect 3500 22278 3512 22330
rect 3512 22278 3542 22330
rect 3566 22278 3576 22330
rect 3576 22278 3622 22330
rect 3326 22276 3382 22278
rect 3406 22276 3462 22278
rect 3486 22276 3542 22278
rect 3566 22276 3622 22278
rect 4274 22330 4330 22332
rect 4354 22330 4410 22332
rect 4434 22330 4490 22332
rect 4514 22330 4570 22332
rect 4274 22278 4320 22330
rect 4320 22278 4330 22330
rect 4354 22278 4384 22330
rect 4384 22278 4396 22330
rect 4396 22278 4410 22330
rect 4434 22278 4448 22330
rect 4448 22278 4460 22330
rect 4460 22278 4490 22330
rect 4514 22278 4524 22330
rect 4524 22278 4570 22330
rect 4274 22276 4330 22278
rect 4354 22276 4410 22278
rect 4434 22276 4490 22278
rect 4514 22276 4570 22278
rect 1904 21786 1960 21788
rect 1984 21786 2040 21788
rect 2064 21786 2120 21788
rect 2144 21786 2200 21788
rect 1904 21734 1950 21786
rect 1950 21734 1960 21786
rect 1984 21734 2014 21786
rect 2014 21734 2026 21786
rect 2026 21734 2040 21786
rect 2064 21734 2078 21786
rect 2078 21734 2090 21786
rect 2090 21734 2120 21786
rect 2144 21734 2154 21786
rect 2154 21734 2200 21786
rect 1904 21732 1960 21734
rect 1984 21732 2040 21734
rect 2064 21732 2120 21734
rect 2144 21732 2200 21734
rect 2852 21786 2908 21788
rect 2932 21786 2988 21788
rect 3012 21786 3068 21788
rect 3092 21786 3148 21788
rect 2852 21734 2898 21786
rect 2898 21734 2908 21786
rect 2932 21734 2962 21786
rect 2962 21734 2974 21786
rect 2974 21734 2988 21786
rect 3012 21734 3026 21786
rect 3026 21734 3038 21786
rect 3038 21734 3068 21786
rect 3092 21734 3102 21786
rect 3102 21734 3148 21786
rect 2852 21732 2908 21734
rect 2932 21732 2988 21734
rect 3012 21732 3068 21734
rect 3092 21732 3148 21734
rect 2378 21242 2434 21244
rect 2458 21242 2514 21244
rect 2538 21242 2594 21244
rect 2618 21242 2674 21244
rect 2378 21190 2424 21242
rect 2424 21190 2434 21242
rect 2458 21190 2488 21242
rect 2488 21190 2500 21242
rect 2500 21190 2514 21242
rect 2538 21190 2552 21242
rect 2552 21190 2564 21242
rect 2564 21190 2594 21242
rect 2618 21190 2628 21242
rect 2628 21190 2674 21242
rect 2378 21188 2434 21190
rect 2458 21188 2514 21190
rect 2538 21188 2594 21190
rect 2618 21188 2674 21190
rect 3326 21242 3382 21244
rect 3406 21242 3462 21244
rect 3486 21242 3542 21244
rect 3566 21242 3622 21244
rect 3326 21190 3372 21242
rect 3372 21190 3382 21242
rect 3406 21190 3436 21242
rect 3436 21190 3448 21242
rect 3448 21190 3462 21242
rect 3486 21190 3500 21242
rect 3500 21190 3512 21242
rect 3512 21190 3542 21242
rect 3566 21190 3576 21242
rect 3576 21190 3622 21242
rect 3326 21188 3382 21190
rect 3406 21188 3462 21190
rect 3486 21188 3542 21190
rect 3566 21188 3622 21190
rect 1904 20698 1960 20700
rect 1984 20698 2040 20700
rect 2064 20698 2120 20700
rect 2144 20698 2200 20700
rect 1904 20646 1950 20698
rect 1950 20646 1960 20698
rect 1984 20646 2014 20698
rect 2014 20646 2026 20698
rect 2026 20646 2040 20698
rect 2064 20646 2078 20698
rect 2078 20646 2090 20698
rect 2090 20646 2120 20698
rect 2144 20646 2154 20698
rect 2154 20646 2200 20698
rect 1904 20644 1960 20646
rect 1984 20644 2040 20646
rect 2064 20644 2120 20646
rect 2144 20644 2200 20646
rect 2852 20698 2908 20700
rect 2932 20698 2988 20700
rect 3012 20698 3068 20700
rect 3092 20698 3148 20700
rect 2852 20646 2898 20698
rect 2898 20646 2908 20698
rect 2932 20646 2962 20698
rect 2962 20646 2974 20698
rect 2974 20646 2988 20698
rect 3012 20646 3026 20698
rect 3026 20646 3038 20698
rect 3038 20646 3068 20698
rect 3092 20646 3102 20698
rect 3102 20646 3148 20698
rect 2852 20644 2908 20646
rect 2932 20644 2988 20646
rect 3012 20644 3068 20646
rect 3092 20644 3148 20646
rect 2378 20154 2434 20156
rect 2458 20154 2514 20156
rect 2538 20154 2594 20156
rect 2618 20154 2674 20156
rect 2378 20102 2424 20154
rect 2424 20102 2434 20154
rect 2458 20102 2488 20154
rect 2488 20102 2500 20154
rect 2500 20102 2514 20154
rect 2538 20102 2552 20154
rect 2552 20102 2564 20154
rect 2564 20102 2594 20154
rect 2618 20102 2628 20154
rect 2628 20102 2674 20154
rect 2378 20100 2434 20102
rect 2458 20100 2514 20102
rect 2538 20100 2594 20102
rect 2618 20100 2674 20102
rect 3800 21786 3856 21788
rect 3880 21786 3936 21788
rect 3960 21786 4016 21788
rect 4040 21786 4096 21788
rect 3800 21734 3846 21786
rect 3846 21734 3856 21786
rect 3880 21734 3910 21786
rect 3910 21734 3922 21786
rect 3922 21734 3936 21786
rect 3960 21734 3974 21786
rect 3974 21734 3986 21786
rect 3986 21734 4016 21786
rect 4040 21734 4050 21786
rect 4050 21734 4096 21786
rect 3800 21732 3856 21734
rect 3880 21732 3936 21734
rect 3960 21732 4016 21734
rect 4040 21732 4096 21734
rect 4250 21664 4306 21720
rect 4274 21242 4330 21244
rect 4354 21242 4410 21244
rect 4434 21242 4490 21244
rect 4514 21242 4570 21244
rect 4274 21190 4320 21242
rect 4320 21190 4330 21242
rect 4354 21190 4384 21242
rect 4384 21190 4396 21242
rect 4396 21190 4410 21242
rect 4434 21190 4448 21242
rect 4448 21190 4460 21242
rect 4460 21190 4490 21242
rect 4514 21190 4524 21242
rect 4524 21190 4570 21242
rect 4274 21188 4330 21190
rect 4354 21188 4410 21190
rect 4434 21188 4490 21190
rect 4514 21188 4570 21190
rect 3800 20698 3856 20700
rect 3880 20698 3936 20700
rect 3960 20698 4016 20700
rect 4040 20698 4096 20700
rect 3800 20646 3846 20698
rect 3846 20646 3856 20698
rect 3880 20646 3910 20698
rect 3910 20646 3922 20698
rect 3922 20646 3936 20698
rect 3960 20646 3974 20698
rect 3974 20646 3986 20698
rect 3986 20646 4016 20698
rect 4040 20646 4050 20698
rect 4050 20646 4096 20698
rect 3800 20644 3856 20646
rect 3880 20644 3936 20646
rect 3960 20644 4016 20646
rect 4040 20644 4096 20646
rect 3326 20154 3382 20156
rect 3406 20154 3462 20156
rect 3486 20154 3542 20156
rect 3566 20154 3622 20156
rect 3326 20102 3372 20154
rect 3372 20102 3382 20154
rect 3406 20102 3436 20154
rect 3436 20102 3448 20154
rect 3448 20102 3462 20154
rect 3486 20102 3500 20154
rect 3500 20102 3512 20154
rect 3512 20102 3542 20154
rect 3566 20102 3576 20154
rect 3576 20102 3622 20154
rect 3326 20100 3382 20102
rect 3406 20100 3462 20102
rect 3486 20100 3542 20102
rect 3566 20100 3622 20102
rect 1904 19610 1960 19612
rect 1984 19610 2040 19612
rect 2064 19610 2120 19612
rect 2144 19610 2200 19612
rect 1904 19558 1950 19610
rect 1950 19558 1960 19610
rect 1984 19558 2014 19610
rect 2014 19558 2026 19610
rect 2026 19558 2040 19610
rect 2064 19558 2078 19610
rect 2078 19558 2090 19610
rect 2090 19558 2120 19610
rect 2144 19558 2154 19610
rect 2154 19558 2200 19610
rect 1904 19556 1960 19558
rect 1984 19556 2040 19558
rect 2064 19556 2120 19558
rect 2144 19556 2200 19558
rect 2852 19610 2908 19612
rect 2932 19610 2988 19612
rect 3012 19610 3068 19612
rect 3092 19610 3148 19612
rect 2852 19558 2898 19610
rect 2898 19558 2908 19610
rect 2932 19558 2962 19610
rect 2962 19558 2974 19610
rect 2974 19558 2988 19610
rect 3012 19558 3026 19610
rect 3026 19558 3038 19610
rect 3038 19558 3068 19610
rect 3092 19558 3102 19610
rect 3102 19558 3148 19610
rect 2852 19556 2908 19558
rect 2932 19556 2988 19558
rect 3012 19556 3068 19558
rect 3092 19556 3148 19558
rect 2378 19066 2434 19068
rect 2458 19066 2514 19068
rect 2538 19066 2594 19068
rect 2618 19066 2674 19068
rect 2378 19014 2424 19066
rect 2424 19014 2434 19066
rect 2458 19014 2488 19066
rect 2488 19014 2500 19066
rect 2500 19014 2514 19066
rect 2538 19014 2552 19066
rect 2552 19014 2564 19066
rect 2564 19014 2594 19066
rect 2618 19014 2628 19066
rect 2628 19014 2674 19066
rect 2378 19012 2434 19014
rect 2458 19012 2514 19014
rect 2538 19012 2594 19014
rect 2618 19012 2674 19014
rect 3238 19352 3294 19408
rect 1904 18522 1960 18524
rect 1984 18522 2040 18524
rect 2064 18522 2120 18524
rect 2144 18522 2200 18524
rect 1904 18470 1950 18522
rect 1950 18470 1960 18522
rect 1984 18470 2014 18522
rect 2014 18470 2026 18522
rect 2026 18470 2040 18522
rect 2064 18470 2078 18522
rect 2078 18470 2090 18522
rect 2090 18470 2120 18522
rect 2144 18470 2154 18522
rect 2154 18470 2200 18522
rect 1904 18468 1960 18470
rect 1984 18468 2040 18470
rect 2064 18468 2120 18470
rect 2144 18468 2200 18470
rect 2852 18522 2908 18524
rect 2932 18522 2988 18524
rect 3012 18522 3068 18524
rect 3092 18522 3148 18524
rect 2852 18470 2898 18522
rect 2898 18470 2908 18522
rect 2932 18470 2962 18522
rect 2962 18470 2974 18522
rect 2974 18470 2988 18522
rect 3012 18470 3026 18522
rect 3026 18470 3038 18522
rect 3038 18470 3068 18522
rect 3092 18470 3102 18522
rect 3102 18470 3148 18522
rect 2852 18468 2908 18470
rect 2932 18468 2988 18470
rect 3012 18468 3068 18470
rect 3092 18468 3148 18470
rect 2378 17978 2434 17980
rect 2458 17978 2514 17980
rect 2538 17978 2594 17980
rect 2618 17978 2674 17980
rect 2378 17926 2424 17978
rect 2424 17926 2434 17978
rect 2458 17926 2488 17978
rect 2488 17926 2500 17978
rect 2500 17926 2514 17978
rect 2538 17926 2552 17978
rect 2552 17926 2564 17978
rect 2564 17926 2594 17978
rect 2618 17926 2628 17978
rect 2628 17926 2674 17978
rect 2378 17924 2434 17926
rect 2458 17924 2514 17926
rect 2538 17924 2594 17926
rect 2618 17924 2674 17926
rect 1904 17434 1960 17436
rect 1984 17434 2040 17436
rect 2064 17434 2120 17436
rect 2144 17434 2200 17436
rect 1904 17382 1950 17434
rect 1950 17382 1960 17434
rect 1984 17382 2014 17434
rect 2014 17382 2026 17434
rect 2026 17382 2040 17434
rect 2064 17382 2078 17434
rect 2078 17382 2090 17434
rect 2090 17382 2120 17434
rect 2144 17382 2154 17434
rect 2154 17382 2200 17434
rect 1904 17380 1960 17382
rect 1984 17380 2040 17382
rect 2064 17380 2120 17382
rect 2144 17380 2200 17382
rect 1430 16890 1486 16892
rect 1510 16890 1566 16892
rect 1590 16890 1646 16892
rect 1670 16890 1726 16892
rect 1430 16838 1476 16890
rect 1476 16838 1486 16890
rect 1510 16838 1540 16890
rect 1540 16838 1552 16890
rect 1552 16838 1566 16890
rect 1590 16838 1604 16890
rect 1604 16838 1616 16890
rect 1616 16838 1646 16890
rect 1670 16838 1680 16890
rect 1680 16838 1726 16890
rect 1430 16836 1486 16838
rect 1510 16836 1566 16838
rect 1590 16836 1646 16838
rect 1670 16836 1726 16838
rect 1306 16360 1362 16416
rect 1904 16346 1960 16348
rect 1984 16346 2040 16348
rect 2064 16346 2120 16348
rect 2144 16346 2200 16348
rect 1904 16294 1950 16346
rect 1950 16294 1960 16346
rect 1984 16294 2014 16346
rect 2014 16294 2026 16346
rect 2026 16294 2040 16346
rect 2064 16294 2078 16346
rect 2078 16294 2090 16346
rect 2090 16294 2120 16346
rect 2144 16294 2154 16346
rect 2154 16294 2200 16346
rect 1904 16292 1960 16294
rect 1984 16292 2040 16294
rect 2064 16292 2120 16294
rect 2144 16292 2200 16294
rect 1430 15802 1486 15804
rect 1510 15802 1566 15804
rect 1590 15802 1646 15804
rect 1670 15802 1726 15804
rect 1430 15750 1476 15802
rect 1476 15750 1486 15802
rect 1510 15750 1540 15802
rect 1540 15750 1552 15802
rect 1552 15750 1566 15802
rect 1590 15750 1604 15802
rect 1604 15750 1616 15802
rect 1616 15750 1646 15802
rect 1670 15750 1680 15802
rect 1680 15750 1726 15802
rect 1430 15748 1486 15750
rect 1510 15748 1566 15750
rect 1590 15748 1646 15750
rect 1670 15748 1726 15750
rect 1904 15258 1960 15260
rect 1984 15258 2040 15260
rect 2064 15258 2120 15260
rect 2144 15258 2200 15260
rect 1904 15206 1950 15258
rect 1950 15206 1960 15258
rect 1984 15206 2014 15258
rect 2014 15206 2026 15258
rect 2026 15206 2040 15258
rect 2064 15206 2078 15258
rect 2078 15206 2090 15258
rect 2090 15206 2120 15258
rect 2144 15206 2154 15258
rect 2154 15206 2200 15258
rect 1904 15204 1960 15206
rect 1984 15204 2040 15206
rect 2064 15204 2120 15206
rect 2144 15204 2200 15206
rect 3326 19066 3382 19068
rect 3406 19066 3462 19068
rect 3486 19066 3542 19068
rect 3566 19066 3622 19068
rect 3326 19014 3372 19066
rect 3372 19014 3382 19066
rect 3406 19014 3436 19066
rect 3436 19014 3448 19066
rect 3448 19014 3462 19066
rect 3486 19014 3500 19066
rect 3500 19014 3512 19066
rect 3512 19014 3542 19066
rect 3566 19014 3576 19066
rect 3576 19014 3622 19066
rect 3326 19012 3382 19014
rect 3406 19012 3462 19014
rect 3486 19012 3542 19014
rect 3566 19012 3622 19014
rect 3326 17978 3382 17980
rect 3406 17978 3462 17980
rect 3486 17978 3542 17980
rect 3566 17978 3622 17980
rect 3326 17926 3372 17978
rect 3372 17926 3382 17978
rect 3406 17926 3436 17978
rect 3436 17926 3448 17978
rect 3448 17926 3462 17978
rect 3486 17926 3500 17978
rect 3500 17926 3512 17978
rect 3512 17926 3542 17978
rect 3566 17926 3576 17978
rect 3576 17926 3622 17978
rect 3326 17924 3382 17926
rect 3406 17924 3462 17926
rect 3486 17924 3542 17926
rect 3566 17924 3622 17926
rect 2852 17434 2908 17436
rect 2932 17434 2988 17436
rect 3012 17434 3068 17436
rect 3092 17434 3148 17436
rect 2852 17382 2898 17434
rect 2898 17382 2908 17434
rect 2932 17382 2962 17434
rect 2962 17382 2974 17434
rect 2974 17382 2988 17434
rect 3012 17382 3026 17434
rect 3026 17382 3038 17434
rect 3038 17382 3068 17434
rect 3092 17382 3102 17434
rect 3102 17382 3148 17434
rect 2852 17380 2908 17382
rect 2932 17380 2988 17382
rect 3012 17380 3068 17382
rect 3092 17380 3148 17382
rect 2378 16890 2434 16892
rect 2458 16890 2514 16892
rect 2538 16890 2594 16892
rect 2618 16890 2674 16892
rect 2378 16838 2424 16890
rect 2424 16838 2434 16890
rect 2458 16838 2488 16890
rect 2488 16838 2500 16890
rect 2500 16838 2514 16890
rect 2538 16838 2552 16890
rect 2552 16838 2564 16890
rect 2564 16838 2594 16890
rect 2618 16838 2628 16890
rect 2628 16838 2674 16890
rect 2378 16836 2434 16838
rect 2458 16836 2514 16838
rect 2538 16836 2594 16838
rect 2618 16836 2674 16838
rect 2852 16346 2908 16348
rect 2932 16346 2988 16348
rect 3012 16346 3068 16348
rect 3092 16346 3148 16348
rect 2852 16294 2898 16346
rect 2898 16294 2908 16346
rect 2932 16294 2962 16346
rect 2962 16294 2974 16346
rect 2974 16294 2988 16346
rect 3012 16294 3026 16346
rect 3026 16294 3038 16346
rect 3038 16294 3068 16346
rect 3092 16294 3102 16346
rect 3102 16294 3148 16346
rect 2852 16292 2908 16294
rect 2932 16292 2988 16294
rect 3012 16292 3068 16294
rect 3092 16292 3148 16294
rect 2378 15802 2434 15804
rect 2458 15802 2514 15804
rect 2538 15802 2594 15804
rect 2618 15802 2674 15804
rect 2378 15750 2424 15802
rect 2424 15750 2434 15802
rect 2458 15750 2488 15802
rect 2488 15750 2500 15802
rect 2500 15750 2514 15802
rect 2538 15750 2552 15802
rect 2552 15750 2564 15802
rect 2564 15750 2594 15802
rect 2618 15750 2628 15802
rect 2628 15750 2674 15802
rect 2378 15748 2434 15750
rect 2458 15748 2514 15750
rect 2538 15748 2594 15750
rect 2618 15748 2674 15750
rect 2852 15258 2908 15260
rect 2932 15258 2988 15260
rect 3012 15258 3068 15260
rect 3092 15258 3148 15260
rect 2852 15206 2898 15258
rect 2898 15206 2908 15258
rect 2932 15206 2962 15258
rect 2962 15206 2974 15258
rect 2974 15206 2988 15258
rect 3012 15206 3026 15258
rect 3026 15206 3038 15258
rect 3038 15206 3068 15258
rect 3092 15206 3102 15258
rect 3102 15206 3148 15258
rect 2852 15204 2908 15206
rect 2932 15204 2988 15206
rect 3012 15204 3068 15206
rect 3092 15204 3148 15206
rect 1430 14714 1486 14716
rect 1510 14714 1566 14716
rect 1590 14714 1646 14716
rect 1670 14714 1726 14716
rect 1430 14662 1476 14714
rect 1476 14662 1486 14714
rect 1510 14662 1540 14714
rect 1540 14662 1552 14714
rect 1552 14662 1566 14714
rect 1590 14662 1604 14714
rect 1604 14662 1616 14714
rect 1616 14662 1646 14714
rect 1670 14662 1680 14714
rect 1680 14662 1726 14714
rect 1430 14660 1486 14662
rect 1510 14660 1566 14662
rect 1590 14660 1646 14662
rect 1670 14660 1726 14662
rect 2378 14714 2434 14716
rect 2458 14714 2514 14716
rect 2538 14714 2594 14716
rect 2618 14714 2674 14716
rect 2378 14662 2424 14714
rect 2424 14662 2434 14714
rect 2458 14662 2488 14714
rect 2488 14662 2500 14714
rect 2500 14662 2514 14714
rect 2538 14662 2552 14714
rect 2552 14662 2564 14714
rect 2564 14662 2594 14714
rect 2618 14662 2628 14714
rect 2628 14662 2674 14714
rect 2378 14660 2434 14662
rect 2458 14660 2514 14662
rect 2538 14660 2594 14662
rect 2618 14660 2674 14662
rect 1430 13626 1486 13628
rect 1510 13626 1566 13628
rect 1590 13626 1646 13628
rect 1670 13626 1726 13628
rect 1430 13574 1476 13626
rect 1476 13574 1486 13626
rect 1510 13574 1540 13626
rect 1540 13574 1552 13626
rect 1552 13574 1566 13626
rect 1590 13574 1604 13626
rect 1604 13574 1616 13626
rect 1616 13574 1646 13626
rect 1670 13574 1680 13626
rect 1680 13574 1726 13626
rect 1430 13572 1486 13574
rect 1510 13572 1566 13574
rect 1590 13572 1646 13574
rect 1670 13572 1726 13574
rect 1582 13368 1638 13424
rect 1904 14170 1960 14172
rect 1984 14170 2040 14172
rect 2064 14170 2120 14172
rect 2144 14170 2200 14172
rect 1904 14118 1950 14170
rect 1950 14118 1960 14170
rect 1984 14118 2014 14170
rect 2014 14118 2026 14170
rect 2026 14118 2040 14170
rect 2064 14118 2078 14170
rect 2078 14118 2090 14170
rect 2090 14118 2120 14170
rect 2144 14118 2154 14170
rect 2154 14118 2200 14170
rect 1904 14116 1960 14118
rect 1984 14116 2040 14118
rect 2064 14116 2120 14118
rect 2144 14116 2200 14118
rect 2852 14170 2908 14172
rect 2932 14170 2988 14172
rect 3012 14170 3068 14172
rect 3092 14170 3148 14172
rect 2852 14118 2898 14170
rect 2898 14118 2908 14170
rect 2932 14118 2962 14170
rect 2962 14118 2974 14170
rect 2974 14118 2988 14170
rect 3012 14118 3026 14170
rect 3026 14118 3038 14170
rect 3038 14118 3068 14170
rect 3092 14118 3102 14170
rect 3102 14118 3148 14170
rect 2852 14116 2908 14118
rect 2932 14116 2988 14118
rect 3012 14116 3068 14118
rect 3092 14116 3148 14118
rect 2378 13626 2434 13628
rect 2458 13626 2514 13628
rect 2538 13626 2594 13628
rect 2618 13626 2674 13628
rect 2378 13574 2424 13626
rect 2424 13574 2434 13626
rect 2458 13574 2488 13626
rect 2488 13574 2500 13626
rect 2500 13574 2514 13626
rect 2538 13574 2552 13626
rect 2552 13574 2564 13626
rect 2564 13574 2594 13626
rect 2618 13574 2628 13626
rect 2628 13574 2674 13626
rect 2378 13572 2434 13574
rect 2458 13572 2514 13574
rect 2538 13572 2594 13574
rect 2618 13572 2674 13574
rect 1904 13082 1960 13084
rect 1984 13082 2040 13084
rect 2064 13082 2120 13084
rect 2144 13082 2200 13084
rect 1904 13030 1950 13082
rect 1950 13030 1960 13082
rect 1984 13030 2014 13082
rect 2014 13030 2026 13082
rect 2026 13030 2040 13082
rect 2064 13030 2078 13082
rect 2078 13030 2090 13082
rect 2090 13030 2120 13082
rect 2144 13030 2154 13082
rect 2154 13030 2200 13082
rect 1904 13028 1960 13030
rect 1984 13028 2040 13030
rect 2064 13028 2120 13030
rect 2144 13028 2200 13030
rect 3326 16890 3382 16892
rect 3406 16890 3462 16892
rect 3486 16890 3542 16892
rect 3566 16890 3622 16892
rect 3326 16838 3372 16890
rect 3372 16838 3382 16890
rect 3406 16838 3436 16890
rect 3436 16838 3448 16890
rect 3448 16838 3462 16890
rect 3486 16838 3500 16890
rect 3500 16838 3512 16890
rect 3512 16838 3542 16890
rect 3566 16838 3576 16890
rect 3576 16838 3622 16890
rect 3326 16836 3382 16838
rect 3406 16836 3462 16838
rect 3486 16836 3542 16838
rect 3566 16836 3622 16838
rect 3326 15802 3382 15804
rect 3406 15802 3462 15804
rect 3486 15802 3542 15804
rect 3566 15802 3622 15804
rect 3326 15750 3372 15802
rect 3372 15750 3382 15802
rect 3406 15750 3436 15802
rect 3436 15750 3448 15802
rect 3448 15750 3462 15802
rect 3486 15750 3500 15802
rect 3500 15750 3512 15802
rect 3512 15750 3542 15802
rect 3566 15750 3576 15802
rect 3576 15750 3622 15802
rect 3326 15748 3382 15750
rect 3406 15748 3462 15750
rect 3486 15748 3542 15750
rect 3566 15748 3622 15750
rect 4710 20168 4766 20224
rect 4274 20154 4330 20156
rect 4354 20154 4410 20156
rect 4434 20154 4490 20156
rect 4514 20154 4570 20156
rect 4274 20102 4320 20154
rect 4320 20102 4330 20154
rect 4354 20102 4384 20154
rect 4384 20102 4396 20154
rect 4396 20102 4410 20154
rect 4434 20102 4448 20154
rect 4448 20102 4460 20154
rect 4460 20102 4490 20154
rect 4514 20102 4524 20154
rect 4524 20102 4570 20154
rect 4274 20100 4330 20102
rect 4354 20100 4410 20102
rect 4434 20100 4490 20102
rect 4514 20100 4570 20102
rect 3800 19610 3856 19612
rect 3880 19610 3936 19612
rect 3960 19610 4016 19612
rect 4040 19610 4096 19612
rect 3800 19558 3846 19610
rect 3846 19558 3856 19610
rect 3880 19558 3910 19610
rect 3910 19558 3922 19610
rect 3922 19558 3936 19610
rect 3960 19558 3974 19610
rect 3974 19558 3986 19610
rect 3986 19558 4016 19610
rect 4040 19558 4050 19610
rect 4050 19558 4096 19610
rect 3800 19556 3856 19558
rect 3880 19556 3936 19558
rect 3960 19556 4016 19558
rect 4040 19556 4096 19558
rect 4274 19066 4330 19068
rect 4354 19066 4410 19068
rect 4434 19066 4490 19068
rect 4514 19066 4570 19068
rect 4274 19014 4320 19066
rect 4320 19014 4330 19066
rect 4354 19014 4384 19066
rect 4384 19014 4396 19066
rect 4396 19014 4410 19066
rect 4434 19014 4448 19066
rect 4448 19014 4460 19066
rect 4460 19014 4490 19066
rect 4514 19014 4524 19066
rect 4524 19014 4570 19066
rect 4274 19012 4330 19014
rect 4354 19012 4410 19014
rect 4434 19012 4490 19014
rect 4514 19012 4570 19014
rect 4158 18708 4160 18728
rect 4160 18708 4212 18728
rect 4212 18708 4214 18728
rect 4158 18672 4214 18708
rect 3800 18522 3856 18524
rect 3880 18522 3936 18524
rect 3960 18522 4016 18524
rect 4040 18522 4096 18524
rect 3800 18470 3846 18522
rect 3846 18470 3856 18522
rect 3880 18470 3910 18522
rect 3910 18470 3922 18522
rect 3922 18470 3936 18522
rect 3960 18470 3974 18522
rect 3974 18470 3986 18522
rect 3986 18470 4016 18522
rect 4040 18470 4050 18522
rect 4050 18470 4096 18522
rect 3800 18468 3856 18470
rect 3880 18468 3936 18470
rect 3960 18468 4016 18470
rect 4040 18468 4096 18470
rect 4274 17978 4330 17980
rect 4354 17978 4410 17980
rect 4434 17978 4490 17980
rect 4514 17978 4570 17980
rect 4274 17926 4320 17978
rect 4320 17926 4330 17978
rect 4354 17926 4384 17978
rect 4384 17926 4396 17978
rect 4396 17926 4410 17978
rect 4434 17926 4448 17978
rect 4448 17926 4460 17978
rect 4460 17926 4490 17978
rect 4514 17926 4524 17978
rect 4524 17926 4570 17978
rect 4274 17924 4330 17926
rect 4354 17924 4410 17926
rect 4434 17924 4490 17926
rect 4514 17924 4570 17926
rect 3800 17434 3856 17436
rect 3880 17434 3936 17436
rect 3960 17434 4016 17436
rect 4040 17434 4096 17436
rect 3800 17382 3846 17434
rect 3846 17382 3856 17434
rect 3880 17382 3910 17434
rect 3910 17382 3922 17434
rect 3922 17382 3936 17434
rect 3960 17382 3974 17434
rect 3974 17382 3986 17434
rect 3986 17382 4016 17434
rect 4040 17382 4050 17434
rect 4050 17382 4096 17434
rect 3800 17380 3856 17382
rect 3880 17380 3936 17382
rect 3960 17380 4016 17382
rect 4040 17380 4096 17382
rect 4158 17176 4214 17232
rect 4274 16890 4330 16892
rect 4354 16890 4410 16892
rect 4434 16890 4490 16892
rect 4514 16890 4570 16892
rect 4274 16838 4320 16890
rect 4320 16838 4330 16890
rect 4354 16838 4384 16890
rect 4384 16838 4396 16890
rect 4396 16838 4410 16890
rect 4434 16838 4448 16890
rect 4448 16838 4460 16890
rect 4460 16838 4490 16890
rect 4514 16838 4524 16890
rect 4524 16838 4570 16890
rect 4274 16836 4330 16838
rect 4354 16836 4410 16838
rect 4434 16836 4490 16838
rect 4514 16836 4570 16838
rect 3800 16346 3856 16348
rect 3880 16346 3936 16348
rect 3960 16346 4016 16348
rect 4040 16346 4096 16348
rect 3800 16294 3846 16346
rect 3846 16294 3856 16346
rect 3880 16294 3910 16346
rect 3910 16294 3922 16346
rect 3922 16294 3936 16346
rect 3960 16294 3974 16346
rect 3974 16294 3986 16346
rect 3986 16294 4016 16346
rect 4040 16294 4050 16346
rect 4050 16294 4096 16346
rect 3800 16292 3856 16294
rect 3880 16292 3936 16294
rect 3960 16292 4016 16294
rect 4040 16292 4096 16294
rect 4274 15802 4330 15804
rect 4354 15802 4410 15804
rect 4434 15802 4490 15804
rect 4514 15802 4570 15804
rect 4274 15750 4320 15802
rect 4320 15750 4330 15802
rect 4354 15750 4384 15802
rect 4384 15750 4396 15802
rect 4396 15750 4410 15802
rect 4434 15750 4448 15802
rect 4448 15750 4460 15802
rect 4460 15750 4490 15802
rect 4514 15750 4524 15802
rect 4524 15750 4570 15802
rect 4274 15748 4330 15750
rect 4354 15748 4410 15750
rect 4434 15748 4490 15750
rect 4514 15748 4570 15750
rect 3800 15258 3856 15260
rect 3880 15258 3936 15260
rect 3960 15258 4016 15260
rect 4040 15258 4096 15260
rect 3800 15206 3846 15258
rect 3846 15206 3856 15258
rect 3880 15206 3910 15258
rect 3910 15206 3922 15258
rect 3922 15206 3936 15258
rect 3960 15206 3974 15258
rect 3974 15206 3986 15258
rect 3986 15206 4016 15258
rect 4040 15206 4050 15258
rect 4050 15206 4096 15258
rect 3800 15204 3856 15206
rect 3880 15204 3936 15206
rect 3960 15204 4016 15206
rect 4040 15204 4096 15206
rect 3326 14714 3382 14716
rect 3406 14714 3462 14716
rect 3486 14714 3542 14716
rect 3566 14714 3622 14716
rect 3326 14662 3372 14714
rect 3372 14662 3382 14714
rect 3406 14662 3436 14714
rect 3436 14662 3448 14714
rect 3448 14662 3462 14714
rect 3486 14662 3500 14714
rect 3500 14662 3512 14714
rect 3512 14662 3542 14714
rect 3566 14662 3576 14714
rect 3576 14662 3622 14714
rect 3326 14660 3382 14662
rect 3406 14660 3462 14662
rect 3486 14660 3542 14662
rect 3566 14660 3622 14662
rect 4274 14714 4330 14716
rect 4354 14714 4410 14716
rect 4434 14714 4490 14716
rect 4514 14714 4570 14716
rect 4274 14662 4320 14714
rect 4320 14662 4330 14714
rect 4354 14662 4384 14714
rect 4384 14662 4396 14714
rect 4396 14662 4410 14714
rect 4434 14662 4448 14714
rect 4448 14662 4460 14714
rect 4460 14662 4490 14714
rect 4514 14662 4524 14714
rect 4524 14662 4570 14714
rect 4274 14660 4330 14662
rect 4354 14660 4410 14662
rect 4434 14660 4490 14662
rect 4514 14660 4570 14662
rect 2852 13082 2908 13084
rect 2932 13082 2988 13084
rect 3012 13082 3068 13084
rect 3092 13082 3148 13084
rect 2852 13030 2898 13082
rect 2898 13030 2908 13082
rect 2932 13030 2962 13082
rect 2962 13030 2974 13082
rect 2974 13030 2988 13082
rect 3012 13030 3026 13082
rect 3026 13030 3038 13082
rect 3038 13030 3068 13082
rect 3092 13030 3102 13082
rect 3102 13030 3148 13082
rect 2852 13028 2908 13030
rect 2932 13028 2988 13030
rect 3012 13028 3068 13030
rect 3092 13028 3148 13030
rect 1430 12538 1486 12540
rect 1510 12538 1566 12540
rect 1590 12538 1646 12540
rect 1670 12538 1726 12540
rect 1430 12486 1476 12538
rect 1476 12486 1486 12538
rect 1510 12486 1540 12538
rect 1540 12486 1552 12538
rect 1552 12486 1566 12538
rect 1590 12486 1604 12538
rect 1604 12486 1616 12538
rect 1616 12486 1646 12538
rect 1670 12486 1680 12538
rect 1680 12486 1726 12538
rect 1430 12484 1486 12486
rect 1510 12484 1566 12486
rect 1590 12484 1646 12486
rect 1670 12484 1726 12486
rect 1430 11450 1486 11452
rect 1510 11450 1566 11452
rect 1590 11450 1646 11452
rect 1670 11450 1726 11452
rect 1430 11398 1476 11450
rect 1476 11398 1486 11450
rect 1510 11398 1540 11450
rect 1540 11398 1552 11450
rect 1552 11398 1566 11450
rect 1590 11398 1604 11450
rect 1604 11398 1616 11450
rect 1616 11398 1646 11450
rect 1670 11398 1680 11450
rect 1680 11398 1726 11450
rect 1430 11396 1486 11398
rect 1510 11396 1566 11398
rect 1590 11396 1646 11398
rect 1670 11396 1726 11398
rect 1398 10512 1454 10568
rect 1430 10362 1486 10364
rect 1510 10362 1566 10364
rect 1590 10362 1646 10364
rect 1670 10362 1726 10364
rect 1430 10310 1476 10362
rect 1476 10310 1486 10362
rect 1510 10310 1540 10362
rect 1540 10310 1552 10362
rect 1552 10310 1566 10362
rect 1590 10310 1604 10362
rect 1604 10310 1616 10362
rect 1616 10310 1646 10362
rect 1670 10310 1680 10362
rect 1680 10310 1726 10362
rect 1430 10308 1486 10310
rect 1510 10308 1566 10310
rect 1590 10308 1646 10310
rect 1670 10308 1726 10310
rect 1904 11994 1960 11996
rect 1984 11994 2040 11996
rect 2064 11994 2120 11996
rect 2144 11994 2200 11996
rect 1904 11942 1950 11994
rect 1950 11942 1960 11994
rect 1984 11942 2014 11994
rect 2014 11942 2026 11994
rect 2026 11942 2040 11994
rect 2064 11942 2078 11994
rect 2078 11942 2090 11994
rect 2090 11942 2120 11994
rect 2144 11942 2154 11994
rect 2154 11942 2200 11994
rect 1904 11940 1960 11942
rect 1984 11940 2040 11942
rect 2064 11940 2120 11942
rect 2144 11940 2200 11942
rect 2378 12538 2434 12540
rect 2458 12538 2514 12540
rect 2538 12538 2594 12540
rect 2618 12538 2674 12540
rect 2378 12486 2424 12538
rect 2424 12486 2434 12538
rect 2458 12486 2488 12538
rect 2488 12486 2500 12538
rect 2500 12486 2514 12538
rect 2538 12486 2552 12538
rect 2552 12486 2564 12538
rect 2564 12486 2594 12538
rect 2618 12486 2628 12538
rect 2628 12486 2674 12538
rect 2378 12484 2434 12486
rect 2458 12484 2514 12486
rect 2538 12484 2594 12486
rect 2618 12484 2674 12486
rect 2318 12280 2374 12336
rect 1904 10906 1960 10908
rect 1984 10906 2040 10908
rect 2064 10906 2120 10908
rect 2144 10906 2200 10908
rect 1904 10854 1950 10906
rect 1950 10854 1960 10906
rect 1984 10854 2014 10906
rect 2014 10854 2026 10906
rect 2026 10854 2040 10906
rect 2064 10854 2078 10906
rect 2078 10854 2090 10906
rect 2090 10854 2120 10906
rect 2144 10854 2154 10906
rect 2154 10854 2200 10906
rect 1904 10852 1960 10854
rect 1984 10852 2040 10854
rect 2064 10852 2120 10854
rect 2144 10852 2200 10854
rect 2870 12280 2926 12336
rect 2852 11994 2908 11996
rect 2932 11994 2988 11996
rect 3012 11994 3068 11996
rect 3092 11994 3148 11996
rect 2852 11942 2898 11994
rect 2898 11942 2908 11994
rect 2932 11942 2962 11994
rect 2962 11942 2974 11994
rect 2974 11942 2988 11994
rect 3012 11942 3026 11994
rect 3026 11942 3038 11994
rect 3038 11942 3068 11994
rect 3092 11942 3102 11994
rect 3102 11942 3148 11994
rect 2852 11940 2908 11942
rect 2932 11940 2988 11942
rect 3012 11940 3068 11942
rect 3092 11940 3148 11942
rect 2378 11450 2434 11452
rect 2458 11450 2514 11452
rect 2538 11450 2594 11452
rect 2618 11450 2674 11452
rect 2378 11398 2424 11450
rect 2424 11398 2434 11450
rect 2458 11398 2488 11450
rect 2488 11398 2500 11450
rect 2500 11398 2514 11450
rect 2538 11398 2552 11450
rect 2552 11398 2564 11450
rect 2564 11398 2594 11450
rect 2618 11398 2628 11450
rect 2628 11398 2674 11450
rect 2378 11396 2434 11398
rect 2458 11396 2514 11398
rect 2538 11396 2594 11398
rect 2618 11396 2674 11398
rect 3326 13626 3382 13628
rect 3406 13626 3462 13628
rect 3486 13626 3542 13628
rect 3566 13626 3622 13628
rect 3326 13574 3372 13626
rect 3372 13574 3382 13626
rect 3406 13574 3436 13626
rect 3436 13574 3448 13626
rect 3448 13574 3462 13626
rect 3486 13574 3500 13626
rect 3500 13574 3512 13626
rect 3512 13574 3542 13626
rect 3566 13574 3576 13626
rect 3576 13574 3622 13626
rect 3326 13572 3382 13574
rect 3406 13572 3462 13574
rect 3486 13572 3542 13574
rect 3566 13572 3622 13574
rect 3326 12538 3382 12540
rect 3406 12538 3462 12540
rect 3486 12538 3542 12540
rect 3566 12538 3622 12540
rect 3326 12486 3372 12538
rect 3372 12486 3382 12538
rect 3406 12486 3436 12538
rect 3436 12486 3448 12538
rect 3448 12486 3462 12538
rect 3486 12486 3500 12538
rect 3500 12486 3512 12538
rect 3512 12486 3542 12538
rect 3566 12486 3576 12538
rect 3576 12486 3622 12538
rect 3326 12484 3382 12486
rect 3406 12484 3462 12486
rect 3486 12484 3542 12486
rect 3566 12484 3622 12486
rect 3800 14170 3856 14172
rect 3880 14170 3936 14172
rect 3960 14170 4016 14172
rect 4040 14170 4096 14172
rect 3800 14118 3846 14170
rect 3846 14118 3856 14170
rect 3880 14118 3910 14170
rect 3910 14118 3922 14170
rect 3922 14118 3936 14170
rect 3960 14118 3974 14170
rect 3974 14118 3986 14170
rect 3986 14118 4016 14170
rect 4040 14118 4050 14170
rect 4050 14118 4096 14170
rect 3800 14116 3856 14118
rect 3880 14116 3936 14118
rect 3960 14116 4016 14118
rect 4040 14116 4096 14118
rect 4250 14184 4306 14240
rect 3800 13082 3856 13084
rect 3880 13082 3936 13084
rect 3960 13082 4016 13084
rect 4040 13082 4096 13084
rect 3800 13030 3846 13082
rect 3846 13030 3856 13082
rect 3880 13030 3910 13082
rect 3910 13030 3922 13082
rect 3922 13030 3936 13082
rect 3960 13030 3974 13082
rect 3974 13030 3986 13082
rect 3986 13030 4016 13082
rect 4040 13030 4050 13082
rect 4050 13030 4096 13082
rect 3800 13028 3856 13030
rect 3880 13028 3936 13030
rect 3960 13028 4016 13030
rect 4040 13028 4096 13030
rect 4274 13626 4330 13628
rect 4354 13626 4410 13628
rect 4434 13626 4490 13628
rect 4514 13626 4570 13628
rect 4274 13574 4320 13626
rect 4320 13574 4330 13626
rect 4354 13574 4384 13626
rect 4384 13574 4396 13626
rect 4396 13574 4410 13626
rect 4434 13574 4448 13626
rect 4448 13574 4460 13626
rect 4460 13574 4490 13626
rect 4514 13574 4524 13626
rect 4524 13574 4570 13626
rect 4274 13572 4330 13574
rect 4354 13572 4410 13574
rect 4434 13572 4490 13574
rect 4514 13572 4570 13574
rect 4066 12688 4122 12744
rect 3800 11994 3856 11996
rect 3880 11994 3936 11996
rect 3960 11994 4016 11996
rect 4040 11994 4096 11996
rect 3800 11942 3846 11994
rect 3846 11942 3856 11994
rect 3880 11942 3910 11994
rect 3910 11942 3922 11994
rect 3922 11942 3936 11994
rect 3960 11942 3974 11994
rect 3974 11942 3986 11994
rect 3986 11942 4016 11994
rect 4040 11942 4050 11994
rect 4050 11942 4096 11994
rect 3800 11940 3856 11942
rect 3880 11940 3936 11942
rect 3960 11940 4016 11942
rect 4040 11940 4096 11942
rect 3326 11450 3382 11452
rect 3406 11450 3462 11452
rect 3486 11450 3542 11452
rect 3566 11450 3622 11452
rect 3326 11398 3372 11450
rect 3372 11398 3382 11450
rect 3406 11398 3436 11450
rect 3436 11398 3448 11450
rect 3448 11398 3462 11450
rect 3486 11398 3500 11450
rect 3500 11398 3512 11450
rect 3512 11398 3542 11450
rect 3566 11398 3576 11450
rect 3576 11398 3622 11450
rect 3326 11396 3382 11398
rect 3406 11396 3462 11398
rect 3486 11396 3542 11398
rect 3566 11396 3622 11398
rect 2852 10906 2908 10908
rect 2932 10906 2988 10908
rect 3012 10906 3068 10908
rect 3092 10906 3148 10908
rect 2852 10854 2898 10906
rect 2898 10854 2908 10906
rect 2932 10854 2962 10906
rect 2962 10854 2974 10906
rect 2974 10854 2988 10906
rect 3012 10854 3026 10906
rect 3026 10854 3038 10906
rect 3038 10854 3068 10906
rect 3092 10854 3102 10906
rect 3102 10854 3148 10906
rect 2852 10852 2908 10854
rect 2932 10852 2988 10854
rect 3012 10852 3068 10854
rect 3092 10852 3148 10854
rect 1904 9818 1960 9820
rect 1984 9818 2040 9820
rect 2064 9818 2120 9820
rect 2144 9818 2200 9820
rect 1904 9766 1950 9818
rect 1950 9766 1960 9818
rect 1984 9766 2014 9818
rect 2014 9766 2026 9818
rect 2026 9766 2040 9818
rect 2064 9766 2078 9818
rect 2078 9766 2090 9818
rect 2090 9766 2120 9818
rect 2144 9766 2154 9818
rect 2154 9766 2200 9818
rect 1904 9764 1960 9766
rect 1984 9764 2040 9766
rect 2064 9764 2120 9766
rect 2144 9764 2200 9766
rect 1214 9560 1270 9616
rect 1430 9274 1486 9276
rect 1510 9274 1566 9276
rect 1590 9274 1646 9276
rect 1670 9274 1726 9276
rect 1430 9222 1476 9274
rect 1476 9222 1486 9274
rect 1510 9222 1540 9274
rect 1540 9222 1552 9274
rect 1552 9222 1566 9274
rect 1590 9222 1604 9274
rect 1604 9222 1616 9274
rect 1616 9222 1646 9274
rect 1670 9222 1680 9274
rect 1680 9222 1726 9274
rect 1430 9220 1486 9222
rect 1510 9220 1566 9222
rect 1590 9220 1646 9222
rect 1670 9220 1726 9222
rect 2378 10362 2434 10364
rect 2458 10362 2514 10364
rect 2538 10362 2594 10364
rect 2618 10362 2674 10364
rect 2378 10310 2424 10362
rect 2424 10310 2434 10362
rect 2458 10310 2488 10362
rect 2488 10310 2500 10362
rect 2500 10310 2514 10362
rect 2538 10310 2552 10362
rect 2552 10310 2564 10362
rect 2564 10310 2594 10362
rect 2618 10310 2628 10362
rect 2628 10310 2674 10362
rect 2378 10308 2434 10310
rect 2458 10308 2514 10310
rect 2538 10308 2594 10310
rect 2618 10308 2674 10310
rect 3422 11228 3424 11248
rect 3424 11228 3476 11248
rect 3476 11228 3478 11248
rect 3422 11192 3478 11228
rect 3514 10512 3570 10568
rect 3800 10906 3856 10908
rect 3880 10906 3936 10908
rect 3960 10906 4016 10908
rect 4040 10906 4096 10908
rect 3800 10854 3846 10906
rect 3846 10854 3856 10906
rect 3880 10854 3910 10906
rect 3910 10854 3922 10906
rect 3922 10854 3936 10906
rect 3960 10854 3974 10906
rect 3974 10854 3986 10906
rect 3986 10854 4016 10906
rect 4040 10854 4050 10906
rect 4050 10854 4096 10906
rect 3800 10852 3856 10854
rect 3880 10852 3936 10854
rect 3960 10852 4016 10854
rect 4040 10852 4096 10854
rect 3326 10362 3382 10364
rect 3406 10362 3462 10364
rect 3486 10362 3542 10364
rect 3566 10362 3622 10364
rect 3326 10310 3372 10362
rect 3372 10310 3382 10362
rect 3406 10310 3436 10362
rect 3436 10310 3448 10362
rect 3448 10310 3462 10362
rect 3486 10310 3500 10362
rect 3500 10310 3512 10362
rect 3512 10310 3542 10362
rect 3566 10310 3576 10362
rect 3576 10310 3622 10362
rect 3326 10308 3382 10310
rect 3406 10308 3462 10310
rect 3486 10308 3542 10310
rect 3566 10308 3622 10310
rect 3238 9968 3294 10024
rect 2852 9818 2908 9820
rect 2932 9818 2988 9820
rect 3012 9818 3068 9820
rect 3092 9818 3148 9820
rect 2852 9766 2898 9818
rect 2898 9766 2908 9818
rect 2932 9766 2962 9818
rect 2962 9766 2974 9818
rect 2974 9766 2988 9818
rect 3012 9766 3026 9818
rect 3026 9766 3038 9818
rect 3038 9766 3068 9818
rect 3092 9766 3102 9818
rect 3102 9766 3148 9818
rect 2852 9764 2908 9766
rect 2932 9764 2988 9766
rect 3012 9764 3068 9766
rect 3092 9764 3148 9766
rect 2778 9560 2834 9616
rect 3606 10104 3662 10160
rect 1904 8730 1960 8732
rect 1984 8730 2040 8732
rect 2064 8730 2120 8732
rect 2144 8730 2200 8732
rect 1904 8678 1950 8730
rect 1950 8678 1960 8730
rect 1984 8678 2014 8730
rect 2014 8678 2026 8730
rect 2026 8678 2040 8730
rect 2064 8678 2078 8730
rect 2078 8678 2090 8730
rect 2090 8678 2120 8730
rect 2144 8678 2154 8730
rect 2154 8678 2200 8730
rect 1904 8676 1960 8678
rect 1984 8676 2040 8678
rect 2064 8676 2120 8678
rect 2144 8676 2200 8678
rect 1430 8186 1486 8188
rect 1510 8186 1566 8188
rect 1590 8186 1646 8188
rect 1670 8186 1726 8188
rect 1430 8134 1476 8186
rect 1476 8134 1486 8186
rect 1510 8134 1540 8186
rect 1540 8134 1552 8186
rect 1552 8134 1566 8186
rect 1590 8134 1604 8186
rect 1604 8134 1616 8186
rect 1616 8134 1646 8186
rect 1670 8134 1680 8186
rect 1680 8134 1726 8186
rect 1430 8132 1486 8134
rect 1510 8132 1566 8134
rect 1590 8132 1646 8134
rect 1670 8132 1726 8134
rect 1398 7384 1454 7440
rect 1430 7098 1486 7100
rect 1510 7098 1566 7100
rect 1590 7098 1646 7100
rect 1670 7098 1726 7100
rect 1430 7046 1476 7098
rect 1476 7046 1486 7098
rect 1510 7046 1540 7098
rect 1540 7046 1552 7098
rect 1552 7046 1566 7098
rect 1590 7046 1604 7098
rect 1604 7046 1616 7098
rect 1616 7046 1646 7098
rect 1670 7046 1680 7098
rect 1680 7046 1726 7098
rect 1430 7044 1486 7046
rect 1510 7044 1566 7046
rect 1590 7044 1646 7046
rect 1670 7044 1726 7046
rect 1904 7642 1960 7644
rect 1984 7642 2040 7644
rect 2064 7642 2120 7644
rect 2144 7642 2200 7644
rect 1904 7590 1950 7642
rect 1950 7590 1960 7642
rect 1984 7590 2014 7642
rect 2014 7590 2026 7642
rect 2026 7590 2040 7642
rect 2064 7590 2078 7642
rect 2078 7590 2090 7642
rect 2090 7590 2120 7642
rect 2144 7590 2154 7642
rect 2154 7590 2200 7642
rect 1904 7588 1960 7590
rect 1984 7588 2040 7590
rect 2064 7588 2120 7590
rect 2144 7588 2200 7590
rect 1904 6554 1960 6556
rect 1984 6554 2040 6556
rect 2064 6554 2120 6556
rect 2144 6554 2200 6556
rect 1904 6502 1950 6554
rect 1950 6502 1960 6554
rect 1984 6502 2014 6554
rect 2014 6502 2026 6554
rect 2026 6502 2040 6554
rect 2064 6502 2078 6554
rect 2078 6502 2090 6554
rect 2090 6502 2120 6554
rect 2144 6502 2154 6554
rect 2154 6502 2200 6554
rect 1904 6500 1960 6502
rect 1984 6500 2040 6502
rect 2064 6500 2120 6502
rect 2144 6500 2200 6502
rect 1430 6010 1486 6012
rect 1510 6010 1566 6012
rect 1590 6010 1646 6012
rect 1670 6010 1726 6012
rect 1430 5958 1476 6010
rect 1476 5958 1486 6010
rect 1510 5958 1540 6010
rect 1540 5958 1552 6010
rect 1552 5958 1566 6010
rect 1590 5958 1604 6010
rect 1604 5958 1616 6010
rect 1616 5958 1646 6010
rect 1670 5958 1680 6010
rect 1680 5958 1726 6010
rect 1430 5956 1486 5958
rect 1510 5956 1566 5958
rect 1590 5956 1646 5958
rect 1670 5956 1726 5958
rect 1430 4922 1486 4924
rect 1510 4922 1566 4924
rect 1590 4922 1646 4924
rect 1670 4922 1726 4924
rect 1430 4870 1476 4922
rect 1476 4870 1486 4922
rect 1510 4870 1540 4922
rect 1540 4870 1552 4922
rect 1552 4870 1566 4922
rect 1590 4870 1604 4922
rect 1604 4870 1616 4922
rect 1616 4870 1646 4922
rect 1670 4870 1680 4922
rect 1680 4870 1726 4922
rect 1430 4868 1486 4870
rect 1510 4868 1566 4870
rect 1590 4868 1646 4870
rect 1670 4868 1726 4870
rect 1398 4392 1454 4448
rect 1430 3834 1486 3836
rect 1510 3834 1566 3836
rect 1590 3834 1646 3836
rect 1670 3834 1726 3836
rect 1430 3782 1476 3834
rect 1476 3782 1486 3834
rect 1510 3782 1540 3834
rect 1540 3782 1552 3834
rect 1552 3782 1566 3834
rect 1590 3782 1604 3834
rect 1604 3782 1616 3834
rect 1616 3782 1646 3834
rect 1670 3782 1680 3834
rect 1680 3782 1726 3834
rect 1430 3780 1486 3782
rect 1510 3780 1566 3782
rect 1590 3780 1646 3782
rect 1670 3780 1726 3782
rect 1430 2746 1486 2748
rect 1510 2746 1566 2748
rect 1590 2746 1646 2748
rect 1670 2746 1726 2748
rect 1430 2694 1476 2746
rect 1476 2694 1486 2746
rect 1510 2694 1540 2746
rect 1540 2694 1552 2746
rect 1552 2694 1566 2746
rect 1590 2694 1604 2746
rect 1604 2694 1616 2746
rect 1616 2694 1646 2746
rect 1670 2694 1680 2746
rect 1680 2694 1726 2746
rect 1430 2692 1486 2694
rect 1510 2692 1566 2694
rect 1590 2692 1646 2694
rect 1670 2692 1726 2694
rect 1430 1658 1486 1660
rect 1510 1658 1566 1660
rect 1590 1658 1646 1660
rect 1670 1658 1726 1660
rect 1430 1606 1476 1658
rect 1476 1606 1486 1658
rect 1510 1606 1540 1658
rect 1540 1606 1552 1658
rect 1552 1606 1566 1658
rect 1590 1606 1604 1658
rect 1604 1606 1616 1658
rect 1616 1606 1646 1658
rect 1670 1606 1680 1658
rect 1680 1606 1726 1658
rect 1430 1604 1486 1606
rect 1510 1604 1566 1606
rect 1590 1604 1646 1606
rect 1670 1604 1726 1606
rect 2378 9274 2434 9276
rect 2458 9274 2514 9276
rect 2538 9274 2594 9276
rect 2618 9274 2674 9276
rect 2378 9222 2424 9274
rect 2424 9222 2434 9274
rect 2458 9222 2488 9274
rect 2488 9222 2500 9274
rect 2500 9222 2514 9274
rect 2538 9222 2552 9274
rect 2552 9222 2564 9274
rect 2564 9222 2594 9274
rect 2618 9222 2628 9274
rect 2628 9222 2674 9274
rect 2378 9220 2434 9222
rect 2458 9220 2514 9222
rect 2538 9220 2594 9222
rect 2618 9220 2674 9222
rect 3326 9274 3382 9276
rect 3406 9274 3462 9276
rect 3486 9274 3542 9276
rect 3566 9274 3622 9276
rect 3326 9222 3372 9274
rect 3372 9222 3382 9274
rect 3406 9222 3436 9274
rect 3436 9222 3448 9274
rect 3448 9222 3462 9274
rect 3486 9222 3500 9274
rect 3500 9222 3512 9274
rect 3512 9222 3542 9274
rect 3566 9222 3576 9274
rect 3576 9222 3622 9274
rect 3326 9220 3382 9222
rect 3406 9220 3462 9222
rect 3486 9220 3542 9222
rect 3566 9220 3622 9222
rect 3800 9818 3856 9820
rect 3880 9818 3936 9820
rect 3960 9818 4016 9820
rect 4040 9818 4096 9820
rect 3800 9766 3846 9818
rect 3846 9766 3856 9818
rect 3880 9766 3910 9818
rect 3910 9766 3922 9818
rect 3922 9766 3936 9818
rect 3960 9766 3974 9818
rect 3974 9766 3986 9818
rect 3986 9766 4016 9818
rect 4040 9766 4050 9818
rect 4050 9766 4096 9818
rect 3800 9764 3856 9766
rect 3880 9764 3936 9766
rect 3960 9764 4016 9766
rect 4040 9764 4096 9766
rect 2852 8730 2908 8732
rect 2932 8730 2988 8732
rect 3012 8730 3068 8732
rect 3092 8730 3148 8732
rect 2852 8678 2898 8730
rect 2898 8678 2908 8730
rect 2932 8678 2962 8730
rect 2962 8678 2974 8730
rect 2974 8678 2988 8730
rect 3012 8678 3026 8730
rect 3026 8678 3038 8730
rect 3038 8678 3068 8730
rect 3092 8678 3102 8730
rect 3102 8678 3148 8730
rect 2852 8676 2908 8678
rect 2932 8676 2988 8678
rect 3012 8676 3068 8678
rect 3092 8676 3148 8678
rect 2378 8186 2434 8188
rect 2458 8186 2514 8188
rect 2538 8186 2594 8188
rect 2618 8186 2674 8188
rect 2378 8134 2424 8186
rect 2424 8134 2434 8186
rect 2458 8134 2488 8186
rect 2488 8134 2500 8186
rect 2500 8134 2514 8186
rect 2538 8134 2552 8186
rect 2552 8134 2564 8186
rect 2564 8134 2594 8186
rect 2618 8134 2628 8186
rect 2628 8134 2674 8186
rect 2378 8132 2434 8134
rect 2458 8132 2514 8134
rect 2538 8132 2594 8134
rect 2618 8132 2674 8134
rect 3326 8186 3382 8188
rect 3406 8186 3462 8188
rect 3486 8186 3542 8188
rect 3566 8186 3622 8188
rect 3326 8134 3372 8186
rect 3372 8134 3382 8186
rect 3406 8134 3436 8186
rect 3436 8134 3448 8186
rect 3448 8134 3462 8186
rect 3486 8134 3500 8186
rect 3500 8134 3512 8186
rect 3512 8134 3542 8186
rect 3566 8134 3576 8186
rect 3576 8134 3622 8186
rect 3326 8132 3382 8134
rect 3406 8132 3462 8134
rect 3486 8132 3542 8134
rect 3566 8132 3622 8134
rect 2852 7642 2908 7644
rect 2932 7642 2988 7644
rect 3012 7642 3068 7644
rect 3092 7642 3148 7644
rect 2852 7590 2898 7642
rect 2898 7590 2908 7642
rect 2932 7590 2962 7642
rect 2962 7590 2974 7642
rect 2974 7590 2988 7642
rect 3012 7590 3026 7642
rect 3026 7590 3038 7642
rect 3038 7590 3068 7642
rect 3092 7590 3102 7642
rect 3102 7590 3148 7642
rect 2852 7588 2908 7590
rect 2932 7588 2988 7590
rect 3012 7588 3068 7590
rect 3092 7588 3148 7590
rect 2378 7098 2434 7100
rect 2458 7098 2514 7100
rect 2538 7098 2594 7100
rect 2618 7098 2674 7100
rect 2378 7046 2424 7098
rect 2424 7046 2434 7098
rect 2458 7046 2488 7098
rect 2488 7046 2500 7098
rect 2500 7046 2514 7098
rect 2538 7046 2552 7098
rect 2552 7046 2564 7098
rect 2564 7046 2594 7098
rect 2618 7046 2628 7098
rect 2628 7046 2674 7098
rect 2378 7044 2434 7046
rect 2458 7044 2514 7046
rect 2538 7044 2594 7046
rect 2618 7044 2674 7046
rect 2852 6554 2908 6556
rect 2932 6554 2988 6556
rect 3012 6554 3068 6556
rect 3092 6554 3148 6556
rect 2852 6502 2898 6554
rect 2898 6502 2908 6554
rect 2932 6502 2962 6554
rect 2962 6502 2974 6554
rect 2974 6502 2988 6554
rect 3012 6502 3026 6554
rect 3026 6502 3038 6554
rect 3038 6502 3068 6554
rect 3092 6502 3102 6554
rect 3102 6502 3148 6554
rect 2852 6500 2908 6502
rect 2932 6500 2988 6502
rect 3012 6500 3068 6502
rect 3092 6500 3148 6502
rect 2378 6010 2434 6012
rect 2458 6010 2514 6012
rect 2538 6010 2594 6012
rect 2618 6010 2674 6012
rect 2378 5958 2424 6010
rect 2424 5958 2434 6010
rect 2458 5958 2488 6010
rect 2488 5958 2500 6010
rect 2500 5958 2514 6010
rect 2538 5958 2552 6010
rect 2552 5958 2564 6010
rect 2564 5958 2594 6010
rect 2618 5958 2628 6010
rect 2628 5958 2674 6010
rect 2378 5956 2434 5958
rect 2458 5956 2514 5958
rect 2538 5956 2594 5958
rect 2618 5956 2674 5958
rect 1904 5466 1960 5468
rect 1984 5466 2040 5468
rect 2064 5466 2120 5468
rect 2144 5466 2200 5468
rect 1904 5414 1950 5466
rect 1950 5414 1960 5466
rect 1984 5414 2014 5466
rect 2014 5414 2026 5466
rect 2026 5414 2040 5466
rect 2064 5414 2078 5466
rect 2078 5414 2090 5466
rect 2090 5414 2120 5466
rect 2144 5414 2154 5466
rect 2154 5414 2200 5466
rect 1904 5412 1960 5414
rect 1984 5412 2040 5414
rect 2064 5412 2120 5414
rect 2144 5412 2200 5414
rect 1904 4378 1960 4380
rect 1984 4378 2040 4380
rect 2064 4378 2120 4380
rect 2144 4378 2200 4380
rect 1904 4326 1950 4378
rect 1950 4326 1960 4378
rect 1984 4326 2014 4378
rect 2014 4326 2026 4378
rect 2026 4326 2040 4378
rect 2064 4326 2078 4378
rect 2078 4326 2090 4378
rect 2090 4326 2120 4378
rect 2144 4326 2154 4378
rect 2154 4326 2200 4378
rect 1904 4324 1960 4326
rect 1984 4324 2040 4326
rect 2064 4324 2120 4326
rect 2144 4324 2200 4326
rect 1904 3290 1960 3292
rect 1984 3290 2040 3292
rect 2064 3290 2120 3292
rect 2144 3290 2200 3292
rect 1904 3238 1950 3290
rect 1950 3238 1960 3290
rect 1984 3238 2014 3290
rect 2014 3238 2026 3290
rect 2026 3238 2040 3290
rect 2064 3238 2078 3290
rect 2078 3238 2090 3290
rect 2090 3238 2120 3290
rect 2144 3238 2154 3290
rect 2154 3238 2200 3290
rect 1904 3236 1960 3238
rect 1984 3236 2040 3238
rect 2064 3236 2120 3238
rect 2144 3236 2200 3238
rect 2852 5466 2908 5468
rect 2932 5466 2988 5468
rect 3012 5466 3068 5468
rect 3092 5466 3148 5468
rect 2852 5414 2898 5466
rect 2898 5414 2908 5466
rect 2932 5414 2962 5466
rect 2962 5414 2974 5466
rect 2974 5414 2988 5466
rect 3012 5414 3026 5466
rect 3026 5414 3038 5466
rect 3038 5414 3068 5466
rect 3092 5414 3102 5466
rect 3102 5414 3148 5466
rect 2852 5412 2908 5414
rect 2932 5412 2988 5414
rect 3012 5412 3068 5414
rect 3092 5412 3148 5414
rect 2378 4922 2434 4924
rect 2458 4922 2514 4924
rect 2538 4922 2594 4924
rect 2618 4922 2674 4924
rect 2378 4870 2424 4922
rect 2424 4870 2434 4922
rect 2458 4870 2488 4922
rect 2488 4870 2500 4922
rect 2500 4870 2514 4922
rect 2538 4870 2552 4922
rect 2552 4870 2564 4922
rect 2564 4870 2594 4922
rect 2618 4870 2628 4922
rect 2628 4870 2674 4922
rect 2378 4868 2434 4870
rect 2458 4868 2514 4870
rect 2538 4868 2594 4870
rect 2618 4868 2674 4870
rect 2852 4378 2908 4380
rect 2932 4378 2988 4380
rect 3012 4378 3068 4380
rect 3092 4378 3148 4380
rect 2852 4326 2898 4378
rect 2898 4326 2908 4378
rect 2932 4326 2962 4378
rect 2962 4326 2974 4378
rect 2974 4326 2988 4378
rect 3012 4326 3026 4378
rect 3026 4326 3038 4378
rect 3038 4326 3068 4378
rect 3092 4326 3102 4378
rect 3102 4326 3148 4378
rect 2852 4324 2908 4326
rect 2932 4324 2988 4326
rect 3012 4324 3068 4326
rect 3092 4324 3148 4326
rect 3326 7098 3382 7100
rect 3406 7098 3462 7100
rect 3486 7098 3542 7100
rect 3566 7098 3622 7100
rect 3326 7046 3372 7098
rect 3372 7046 3382 7098
rect 3406 7046 3436 7098
rect 3436 7046 3448 7098
rect 3448 7046 3462 7098
rect 3486 7046 3500 7098
rect 3500 7046 3512 7098
rect 3512 7046 3542 7098
rect 3566 7046 3576 7098
rect 3576 7046 3622 7098
rect 3326 7044 3382 7046
rect 3406 7044 3462 7046
rect 3486 7044 3542 7046
rect 3566 7044 3622 7046
rect 3800 8730 3856 8732
rect 3880 8730 3936 8732
rect 3960 8730 4016 8732
rect 4040 8730 4096 8732
rect 3800 8678 3846 8730
rect 3846 8678 3856 8730
rect 3880 8678 3910 8730
rect 3910 8678 3922 8730
rect 3922 8678 3936 8730
rect 3960 8678 3974 8730
rect 3974 8678 3986 8730
rect 3986 8678 4016 8730
rect 4040 8678 4050 8730
rect 4050 8678 4096 8730
rect 3800 8676 3856 8678
rect 3880 8676 3936 8678
rect 3960 8676 4016 8678
rect 4040 8676 4096 8678
rect 3800 7642 3856 7644
rect 3880 7642 3936 7644
rect 3960 7642 4016 7644
rect 4040 7642 4096 7644
rect 3800 7590 3846 7642
rect 3846 7590 3856 7642
rect 3880 7590 3910 7642
rect 3910 7590 3922 7642
rect 3922 7590 3936 7642
rect 3960 7590 3974 7642
rect 3974 7590 3986 7642
rect 3986 7590 4016 7642
rect 4040 7590 4050 7642
rect 4050 7590 4096 7642
rect 3800 7588 3856 7590
rect 3880 7588 3936 7590
rect 3960 7588 4016 7590
rect 4040 7588 4096 7590
rect 4710 15680 4766 15736
rect 4274 12538 4330 12540
rect 4354 12538 4410 12540
rect 4434 12538 4490 12540
rect 4514 12538 4570 12540
rect 4274 12486 4320 12538
rect 4320 12486 4330 12538
rect 4354 12486 4384 12538
rect 4384 12486 4396 12538
rect 4396 12486 4410 12538
rect 4434 12486 4448 12538
rect 4448 12486 4460 12538
rect 4460 12486 4490 12538
rect 4514 12486 4524 12538
rect 4524 12486 4570 12538
rect 4274 12484 4330 12486
rect 4354 12484 4410 12486
rect 4434 12484 4490 12486
rect 4514 12484 4570 12486
rect 4274 11450 4330 11452
rect 4354 11450 4410 11452
rect 4434 11450 4490 11452
rect 4514 11450 4570 11452
rect 4274 11398 4320 11450
rect 4320 11398 4330 11450
rect 4354 11398 4384 11450
rect 4384 11398 4396 11450
rect 4396 11398 4410 11450
rect 4434 11398 4448 11450
rect 4448 11398 4460 11450
rect 4460 11398 4490 11450
rect 4514 11398 4524 11450
rect 4524 11398 4570 11450
rect 4274 11396 4330 11398
rect 4354 11396 4410 11398
rect 4434 11396 4490 11398
rect 4514 11396 4570 11398
rect 4274 10362 4330 10364
rect 4354 10362 4410 10364
rect 4434 10362 4490 10364
rect 4514 10362 4570 10364
rect 4274 10310 4320 10362
rect 4320 10310 4330 10362
rect 4354 10310 4384 10362
rect 4384 10310 4396 10362
rect 4396 10310 4410 10362
rect 4434 10310 4448 10362
rect 4448 10310 4460 10362
rect 4460 10310 4490 10362
rect 4514 10310 4524 10362
rect 4524 10310 4570 10362
rect 4274 10308 4330 10310
rect 4354 10308 4410 10310
rect 4434 10308 4490 10310
rect 4514 10308 4570 10310
rect 4274 9274 4330 9276
rect 4354 9274 4410 9276
rect 4434 9274 4490 9276
rect 4514 9274 4570 9276
rect 4274 9222 4320 9274
rect 4320 9222 4330 9274
rect 4354 9222 4384 9274
rect 4384 9222 4396 9274
rect 4396 9222 4410 9274
rect 4434 9222 4448 9274
rect 4448 9222 4460 9274
rect 4460 9222 4490 9274
rect 4514 9222 4524 9274
rect 4524 9222 4570 9274
rect 4274 9220 4330 9222
rect 4354 9220 4410 9222
rect 4434 9220 4490 9222
rect 4514 9220 4570 9222
rect 4710 8200 4766 8256
rect 4274 8186 4330 8188
rect 4354 8186 4410 8188
rect 4434 8186 4490 8188
rect 4514 8186 4570 8188
rect 4274 8134 4320 8186
rect 4320 8134 4330 8186
rect 4354 8134 4384 8186
rect 4384 8134 4396 8186
rect 4396 8134 4410 8186
rect 4434 8134 4448 8186
rect 4448 8134 4460 8186
rect 4460 8134 4490 8186
rect 4514 8134 4524 8186
rect 4524 8134 4570 8186
rect 4274 8132 4330 8134
rect 4354 8132 4410 8134
rect 4434 8132 4490 8134
rect 4514 8132 4570 8134
rect 3698 6704 3754 6760
rect 3800 6554 3856 6556
rect 3880 6554 3936 6556
rect 3960 6554 4016 6556
rect 4040 6554 4096 6556
rect 3800 6502 3846 6554
rect 3846 6502 3856 6554
rect 3880 6502 3910 6554
rect 3910 6502 3922 6554
rect 3922 6502 3936 6554
rect 3960 6502 3974 6554
rect 3974 6502 3986 6554
rect 3986 6502 4016 6554
rect 4040 6502 4050 6554
rect 4050 6502 4096 6554
rect 3800 6500 3856 6502
rect 3880 6500 3936 6502
rect 3960 6500 4016 6502
rect 4040 6500 4096 6502
rect 3326 6010 3382 6012
rect 3406 6010 3462 6012
rect 3486 6010 3542 6012
rect 3566 6010 3622 6012
rect 3326 5958 3372 6010
rect 3372 5958 3382 6010
rect 3406 5958 3436 6010
rect 3436 5958 3448 6010
rect 3448 5958 3462 6010
rect 3486 5958 3500 6010
rect 3500 5958 3512 6010
rect 3512 5958 3542 6010
rect 3566 5958 3576 6010
rect 3576 5958 3622 6010
rect 3326 5956 3382 5958
rect 3406 5956 3462 5958
rect 3486 5956 3542 5958
rect 3566 5956 3622 5958
rect 3800 5466 3856 5468
rect 3880 5466 3936 5468
rect 3960 5466 4016 5468
rect 4040 5466 4096 5468
rect 3800 5414 3846 5466
rect 3846 5414 3856 5466
rect 3880 5414 3910 5466
rect 3910 5414 3922 5466
rect 3922 5414 3936 5466
rect 3960 5414 3974 5466
rect 3974 5414 3986 5466
rect 3986 5414 4016 5466
rect 4040 5414 4050 5466
rect 4050 5414 4096 5466
rect 3800 5412 3856 5414
rect 3880 5412 3936 5414
rect 3960 5412 4016 5414
rect 4040 5412 4096 5414
rect 4274 7098 4330 7100
rect 4354 7098 4410 7100
rect 4434 7098 4490 7100
rect 4514 7098 4570 7100
rect 4274 7046 4320 7098
rect 4320 7046 4330 7098
rect 4354 7046 4384 7098
rect 4384 7046 4396 7098
rect 4396 7046 4410 7098
rect 4434 7046 4448 7098
rect 4448 7046 4460 7098
rect 4460 7046 4490 7098
rect 4514 7046 4524 7098
rect 4524 7046 4570 7098
rect 4274 7044 4330 7046
rect 4354 7044 4410 7046
rect 4434 7044 4490 7046
rect 4514 7044 4570 7046
rect 4274 6010 4330 6012
rect 4354 6010 4410 6012
rect 4434 6010 4490 6012
rect 4514 6010 4570 6012
rect 4274 5958 4320 6010
rect 4320 5958 4330 6010
rect 4354 5958 4384 6010
rect 4384 5958 4396 6010
rect 4396 5958 4410 6010
rect 4434 5958 4448 6010
rect 4448 5958 4460 6010
rect 4460 5958 4490 6010
rect 4514 5958 4524 6010
rect 4524 5958 4570 6010
rect 4274 5956 4330 5958
rect 4354 5956 4410 5958
rect 4434 5956 4490 5958
rect 4514 5956 4570 5958
rect 4158 5208 4214 5264
rect 3326 4922 3382 4924
rect 3406 4922 3462 4924
rect 3486 4922 3542 4924
rect 3566 4922 3622 4924
rect 3326 4870 3372 4922
rect 3372 4870 3382 4922
rect 3406 4870 3436 4922
rect 3436 4870 3448 4922
rect 3448 4870 3462 4922
rect 3486 4870 3500 4922
rect 3500 4870 3512 4922
rect 3512 4870 3542 4922
rect 3566 4870 3576 4922
rect 3576 4870 3622 4922
rect 3326 4868 3382 4870
rect 3406 4868 3462 4870
rect 3486 4868 3542 4870
rect 3566 4868 3622 4870
rect 4274 4922 4330 4924
rect 4354 4922 4410 4924
rect 4434 4922 4490 4924
rect 4514 4922 4570 4924
rect 4274 4870 4320 4922
rect 4320 4870 4330 4922
rect 4354 4870 4384 4922
rect 4384 4870 4396 4922
rect 4396 4870 4410 4922
rect 4434 4870 4448 4922
rect 4448 4870 4460 4922
rect 4460 4870 4490 4922
rect 4514 4870 4524 4922
rect 4524 4870 4570 4922
rect 4274 4868 4330 4870
rect 4354 4868 4410 4870
rect 4434 4868 4490 4870
rect 4514 4868 4570 4870
rect 3800 4378 3856 4380
rect 3880 4378 3936 4380
rect 3960 4378 4016 4380
rect 4040 4378 4096 4380
rect 3800 4326 3846 4378
rect 3846 4326 3856 4378
rect 3880 4326 3910 4378
rect 3910 4326 3922 4378
rect 3922 4326 3936 4378
rect 3960 4326 3974 4378
rect 3974 4326 3986 4378
rect 3986 4326 4016 4378
rect 4040 4326 4050 4378
rect 4050 4326 4096 4378
rect 3800 4324 3856 4326
rect 3880 4324 3936 4326
rect 3960 4324 4016 4326
rect 4040 4324 4096 4326
rect 3238 3984 3294 4040
rect 2378 3834 2434 3836
rect 2458 3834 2514 3836
rect 2538 3834 2594 3836
rect 2618 3834 2674 3836
rect 2378 3782 2424 3834
rect 2424 3782 2434 3834
rect 2458 3782 2488 3834
rect 2488 3782 2500 3834
rect 2500 3782 2514 3834
rect 2538 3782 2552 3834
rect 2552 3782 2564 3834
rect 2564 3782 2594 3834
rect 2618 3782 2628 3834
rect 2628 3782 2674 3834
rect 2378 3780 2434 3782
rect 2458 3780 2514 3782
rect 2538 3780 2594 3782
rect 2618 3780 2674 3782
rect 3326 3834 3382 3836
rect 3406 3834 3462 3836
rect 3486 3834 3542 3836
rect 3566 3834 3622 3836
rect 3326 3782 3372 3834
rect 3372 3782 3382 3834
rect 3406 3782 3436 3834
rect 3436 3782 3448 3834
rect 3448 3782 3462 3834
rect 3486 3782 3500 3834
rect 3500 3782 3512 3834
rect 3512 3782 3542 3834
rect 3566 3782 3576 3834
rect 3576 3782 3622 3834
rect 3326 3780 3382 3782
rect 3406 3780 3462 3782
rect 3486 3780 3542 3782
rect 3566 3780 3622 3782
rect 4274 3834 4330 3836
rect 4354 3834 4410 3836
rect 4434 3834 4490 3836
rect 4514 3834 4570 3836
rect 4274 3782 4320 3834
rect 4320 3782 4330 3834
rect 4354 3782 4384 3834
rect 4384 3782 4396 3834
rect 4396 3782 4410 3834
rect 4434 3782 4448 3834
rect 4448 3782 4460 3834
rect 4460 3782 4490 3834
rect 4514 3782 4524 3834
rect 4524 3782 4570 3834
rect 4274 3780 4330 3782
rect 4354 3780 4410 3782
rect 4434 3780 4490 3782
rect 4514 3780 4570 3782
rect 2852 3290 2908 3292
rect 2932 3290 2988 3292
rect 3012 3290 3068 3292
rect 3092 3290 3148 3292
rect 2852 3238 2898 3290
rect 2898 3238 2908 3290
rect 2932 3238 2962 3290
rect 2962 3238 2974 3290
rect 2974 3238 2988 3290
rect 3012 3238 3026 3290
rect 3026 3238 3038 3290
rect 3038 3238 3068 3290
rect 3092 3238 3102 3290
rect 3102 3238 3148 3290
rect 2852 3236 2908 3238
rect 2932 3236 2988 3238
rect 3012 3236 3068 3238
rect 3092 3236 3148 3238
rect 3800 3290 3856 3292
rect 3880 3290 3936 3292
rect 3960 3290 4016 3292
rect 4040 3290 4096 3292
rect 3800 3238 3846 3290
rect 3846 3238 3856 3290
rect 3880 3238 3910 3290
rect 3910 3238 3922 3290
rect 3922 3238 3936 3290
rect 3960 3238 3974 3290
rect 3974 3238 3986 3290
rect 3986 3238 4016 3290
rect 4040 3238 4050 3290
rect 4050 3238 4096 3290
rect 3800 3236 3856 3238
rect 3880 3236 3936 3238
rect 3960 3236 4016 3238
rect 4040 3236 4096 3238
rect 2378 2746 2434 2748
rect 2458 2746 2514 2748
rect 2538 2746 2594 2748
rect 2618 2746 2674 2748
rect 2378 2694 2424 2746
rect 2424 2694 2434 2746
rect 2458 2694 2488 2746
rect 2488 2694 2500 2746
rect 2500 2694 2514 2746
rect 2538 2694 2552 2746
rect 2552 2694 2564 2746
rect 2564 2694 2594 2746
rect 2618 2694 2628 2746
rect 2628 2694 2674 2746
rect 2378 2692 2434 2694
rect 2458 2692 2514 2694
rect 2538 2692 2594 2694
rect 2618 2692 2674 2694
rect 3326 2746 3382 2748
rect 3406 2746 3462 2748
rect 3486 2746 3542 2748
rect 3566 2746 3622 2748
rect 3326 2694 3372 2746
rect 3372 2694 3382 2746
rect 3406 2694 3436 2746
rect 3436 2694 3448 2746
rect 3448 2694 3462 2746
rect 3486 2694 3500 2746
rect 3500 2694 3512 2746
rect 3512 2694 3542 2746
rect 3566 2694 3576 2746
rect 3576 2694 3622 2746
rect 3326 2692 3382 2694
rect 3406 2692 3462 2694
rect 3486 2692 3542 2694
rect 3566 2692 3622 2694
rect 4274 2746 4330 2748
rect 4354 2746 4410 2748
rect 4434 2746 4490 2748
rect 4514 2746 4570 2748
rect 4274 2694 4320 2746
rect 4320 2694 4330 2746
rect 4354 2694 4384 2746
rect 4384 2694 4396 2746
rect 4396 2694 4410 2746
rect 4434 2694 4448 2746
rect 4448 2694 4460 2746
rect 4460 2694 4490 2746
rect 4514 2694 4524 2746
rect 4524 2694 4570 2746
rect 4274 2692 4330 2694
rect 4354 2692 4410 2694
rect 4434 2692 4490 2694
rect 4514 2692 4570 2694
rect 2226 2352 2282 2408
rect 1904 2202 1960 2204
rect 1984 2202 2040 2204
rect 2064 2202 2120 2204
rect 2144 2202 2200 2204
rect 1904 2150 1950 2202
rect 1950 2150 1960 2202
rect 1984 2150 2014 2202
rect 2014 2150 2026 2202
rect 2026 2150 2040 2202
rect 2064 2150 2078 2202
rect 2078 2150 2090 2202
rect 2090 2150 2120 2202
rect 2144 2150 2154 2202
rect 2154 2150 2200 2202
rect 1904 2148 1960 2150
rect 1984 2148 2040 2150
rect 2064 2148 2120 2150
rect 2144 2148 2200 2150
rect 2852 2202 2908 2204
rect 2932 2202 2988 2204
rect 3012 2202 3068 2204
rect 3092 2202 3148 2204
rect 2852 2150 2898 2202
rect 2898 2150 2908 2202
rect 2932 2150 2962 2202
rect 2962 2150 2974 2202
rect 2974 2150 2988 2202
rect 3012 2150 3026 2202
rect 3026 2150 3038 2202
rect 3038 2150 3068 2202
rect 3092 2150 3102 2202
rect 3102 2150 3148 2202
rect 2852 2148 2908 2150
rect 2932 2148 2988 2150
rect 3012 2148 3068 2150
rect 3092 2148 3148 2150
rect 3800 2202 3856 2204
rect 3880 2202 3936 2204
rect 3960 2202 4016 2204
rect 4040 2202 4096 2204
rect 3800 2150 3846 2202
rect 3846 2150 3856 2202
rect 3880 2150 3910 2202
rect 3910 2150 3922 2202
rect 3922 2150 3936 2202
rect 3960 2150 3974 2202
rect 3974 2150 3986 2202
rect 3986 2150 4016 2202
rect 4040 2150 4050 2202
rect 4050 2150 4096 2202
rect 3800 2148 3856 2150
rect 3880 2148 3936 2150
rect 3960 2148 4016 2150
rect 4040 2148 4096 2150
rect 2378 1658 2434 1660
rect 2458 1658 2514 1660
rect 2538 1658 2594 1660
rect 2618 1658 2674 1660
rect 2378 1606 2424 1658
rect 2424 1606 2434 1658
rect 2458 1606 2488 1658
rect 2488 1606 2500 1658
rect 2500 1606 2514 1658
rect 2538 1606 2552 1658
rect 2552 1606 2564 1658
rect 2564 1606 2594 1658
rect 2618 1606 2628 1658
rect 2628 1606 2674 1658
rect 2378 1604 2434 1606
rect 2458 1604 2514 1606
rect 2538 1604 2594 1606
rect 2618 1604 2674 1606
rect 3326 1658 3382 1660
rect 3406 1658 3462 1660
rect 3486 1658 3542 1660
rect 3566 1658 3622 1660
rect 3326 1606 3372 1658
rect 3372 1606 3382 1658
rect 3406 1606 3436 1658
rect 3436 1606 3448 1658
rect 3448 1606 3462 1658
rect 3486 1606 3500 1658
rect 3500 1606 3512 1658
rect 3512 1606 3542 1658
rect 3566 1606 3576 1658
rect 3576 1606 3622 1658
rect 3326 1604 3382 1606
rect 3406 1604 3462 1606
rect 3486 1604 3542 1606
rect 3566 1604 3622 1606
rect 4274 1658 4330 1660
rect 4354 1658 4410 1660
rect 4434 1658 4490 1660
rect 4514 1658 4570 1660
rect 4274 1606 4320 1658
rect 4320 1606 4330 1658
rect 4354 1606 4384 1658
rect 4384 1606 4396 1658
rect 4396 1606 4410 1658
rect 4434 1606 4448 1658
rect 4448 1606 4460 1658
rect 4460 1606 4490 1658
rect 4514 1606 4524 1658
rect 4524 1606 4570 1658
rect 4274 1604 4330 1606
rect 4354 1604 4410 1606
rect 4434 1604 4490 1606
rect 4514 1604 4570 1606
rect 1766 1400 1822 1456
rect 1904 1114 1960 1116
rect 1984 1114 2040 1116
rect 2064 1114 2120 1116
rect 2144 1114 2200 1116
rect 1904 1062 1950 1114
rect 1950 1062 1960 1114
rect 1984 1062 2014 1114
rect 2014 1062 2026 1114
rect 2026 1062 2040 1114
rect 2064 1062 2078 1114
rect 2078 1062 2090 1114
rect 2090 1062 2120 1114
rect 2144 1062 2154 1114
rect 2154 1062 2200 1114
rect 1904 1060 1960 1062
rect 1984 1060 2040 1062
rect 2064 1060 2120 1062
rect 2144 1060 2200 1062
rect 2852 1114 2908 1116
rect 2932 1114 2988 1116
rect 3012 1114 3068 1116
rect 3092 1114 3148 1116
rect 2852 1062 2898 1114
rect 2898 1062 2908 1114
rect 2932 1062 2962 1114
rect 2962 1062 2974 1114
rect 2974 1062 2988 1114
rect 3012 1062 3026 1114
rect 3026 1062 3038 1114
rect 3038 1062 3068 1114
rect 3092 1062 3102 1114
rect 3102 1062 3148 1114
rect 2852 1060 2908 1062
rect 2932 1060 2988 1062
rect 3012 1060 3068 1062
rect 3092 1060 3148 1062
rect 3800 1114 3856 1116
rect 3880 1114 3936 1116
rect 3960 1114 4016 1116
rect 4040 1114 4096 1116
rect 3800 1062 3846 1114
rect 3846 1062 3856 1114
rect 3880 1062 3910 1114
rect 3910 1062 3922 1114
rect 3922 1062 3936 1114
rect 3960 1062 3974 1114
rect 3974 1062 3986 1114
rect 3986 1062 4016 1114
rect 4040 1062 4050 1114
rect 4050 1062 4096 1114
rect 3800 1060 3856 1062
rect 3880 1060 3936 1062
rect 3960 1060 4016 1062
rect 4040 1060 4096 1062
rect 4710 720 4766 776
<< metal3 >>
rect 4153 23218 4219 23221
rect 5200 23218 6000 23248
rect 4153 23216 6000 23218
rect 4153 23160 4158 23216
rect 4214 23160 6000 23216
rect 4153 23158 6000 23160
rect 4153 23155 4219 23158
rect 5200 23128 6000 23158
rect 1894 22880 2210 22881
rect 1894 22816 1900 22880
rect 1964 22816 1980 22880
rect 2044 22816 2060 22880
rect 2124 22816 2140 22880
rect 2204 22816 2210 22880
rect 1894 22815 2210 22816
rect 2842 22880 3158 22881
rect 2842 22816 2848 22880
rect 2912 22816 2928 22880
rect 2992 22816 3008 22880
rect 3072 22816 3088 22880
rect 3152 22816 3158 22880
rect 2842 22815 3158 22816
rect 3790 22880 4106 22881
rect 3790 22816 3796 22880
rect 3860 22816 3876 22880
rect 3940 22816 3956 22880
rect 4020 22816 4036 22880
rect 4100 22816 4106 22880
rect 3790 22815 4106 22816
rect 0 22402 800 22432
rect 0 22342 1226 22402
rect 0 22312 800 22342
rect 1166 22130 1226 22342
rect 1420 22336 1736 22337
rect 1420 22272 1426 22336
rect 1490 22272 1506 22336
rect 1570 22272 1586 22336
rect 1650 22272 1666 22336
rect 1730 22272 1736 22336
rect 1420 22271 1736 22272
rect 2368 22336 2684 22337
rect 2368 22272 2374 22336
rect 2438 22272 2454 22336
rect 2518 22272 2534 22336
rect 2598 22272 2614 22336
rect 2678 22272 2684 22336
rect 2368 22271 2684 22272
rect 3316 22336 3632 22337
rect 3316 22272 3322 22336
rect 3386 22272 3402 22336
rect 3466 22272 3482 22336
rect 3546 22272 3562 22336
rect 3626 22272 3632 22336
rect 3316 22271 3632 22272
rect 4264 22336 4580 22337
rect 4264 22272 4270 22336
rect 4334 22272 4350 22336
rect 4414 22272 4430 22336
rect 4494 22272 4510 22336
rect 4574 22272 4580 22336
rect 4264 22271 4580 22272
rect 1761 22130 1827 22133
rect 1166 22128 1827 22130
rect 1166 22072 1766 22128
rect 1822 22072 1827 22128
rect 1166 22070 1827 22072
rect 1761 22067 1827 22070
rect 1894 21792 2210 21793
rect 1894 21728 1900 21792
rect 1964 21728 1980 21792
rect 2044 21728 2060 21792
rect 2124 21728 2140 21792
rect 2204 21728 2210 21792
rect 1894 21727 2210 21728
rect 2842 21792 3158 21793
rect 2842 21728 2848 21792
rect 2912 21728 2928 21792
rect 2992 21728 3008 21792
rect 3072 21728 3088 21792
rect 3152 21728 3158 21792
rect 2842 21727 3158 21728
rect 3790 21792 4106 21793
rect 3790 21728 3796 21792
rect 3860 21728 3876 21792
rect 3940 21728 3956 21792
rect 4020 21728 4036 21792
rect 4100 21728 4106 21792
rect 3790 21727 4106 21728
rect 4245 21722 4311 21725
rect 5200 21722 6000 21752
rect 4245 21720 6000 21722
rect 4245 21664 4250 21720
rect 4306 21664 6000 21720
rect 4245 21662 6000 21664
rect 4245 21659 4311 21662
rect 5200 21632 6000 21662
rect 1420 21248 1736 21249
rect 1420 21184 1426 21248
rect 1490 21184 1506 21248
rect 1570 21184 1586 21248
rect 1650 21184 1666 21248
rect 1730 21184 1736 21248
rect 1420 21183 1736 21184
rect 2368 21248 2684 21249
rect 2368 21184 2374 21248
rect 2438 21184 2454 21248
rect 2518 21184 2534 21248
rect 2598 21184 2614 21248
rect 2678 21184 2684 21248
rect 2368 21183 2684 21184
rect 3316 21248 3632 21249
rect 3316 21184 3322 21248
rect 3386 21184 3402 21248
rect 3466 21184 3482 21248
rect 3546 21184 3562 21248
rect 3626 21184 3632 21248
rect 3316 21183 3632 21184
rect 4264 21248 4580 21249
rect 4264 21184 4270 21248
rect 4334 21184 4350 21248
rect 4414 21184 4430 21248
rect 4494 21184 4510 21248
rect 4574 21184 4580 21248
rect 4264 21183 4580 21184
rect 1894 20704 2210 20705
rect 1894 20640 1900 20704
rect 1964 20640 1980 20704
rect 2044 20640 2060 20704
rect 2124 20640 2140 20704
rect 2204 20640 2210 20704
rect 1894 20639 2210 20640
rect 2842 20704 3158 20705
rect 2842 20640 2848 20704
rect 2912 20640 2928 20704
rect 2992 20640 3008 20704
rect 3072 20640 3088 20704
rect 3152 20640 3158 20704
rect 2842 20639 3158 20640
rect 3790 20704 4106 20705
rect 3790 20640 3796 20704
rect 3860 20640 3876 20704
rect 3940 20640 3956 20704
rect 4020 20640 4036 20704
rect 4100 20640 4106 20704
rect 3790 20639 4106 20640
rect 4705 20226 4771 20229
rect 5200 20226 6000 20256
rect 4705 20224 6000 20226
rect 4705 20168 4710 20224
rect 4766 20168 6000 20224
rect 4705 20166 6000 20168
rect 4705 20163 4771 20166
rect 1420 20160 1736 20161
rect 1420 20096 1426 20160
rect 1490 20096 1506 20160
rect 1570 20096 1586 20160
rect 1650 20096 1666 20160
rect 1730 20096 1736 20160
rect 1420 20095 1736 20096
rect 2368 20160 2684 20161
rect 2368 20096 2374 20160
rect 2438 20096 2454 20160
rect 2518 20096 2534 20160
rect 2598 20096 2614 20160
rect 2678 20096 2684 20160
rect 2368 20095 2684 20096
rect 3316 20160 3632 20161
rect 3316 20096 3322 20160
rect 3386 20096 3402 20160
rect 3466 20096 3482 20160
rect 3546 20096 3562 20160
rect 3626 20096 3632 20160
rect 3316 20095 3632 20096
rect 4264 20160 4580 20161
rect 4264 20096 4270 20160
rect 4334 20096 4350 20160
rect 4414 20096 4430 20160
rect 4494 20096 4510 20160
rect 4574 20096 4580 20160
rect 5200 20136 6000 20166
rect 4264 20095 4580 20096
rect 1894 19616 2210 19617
rect 1894 19552 1900 19616
rect 1964 19552 1980 19616
rect 2044 19552 2060 19616
rect 2124 19552 2140 19616
rect 2204 19552 2210 19616
rect 1894 19551 2210 19552
rect 2842 19616 3158 19617
rect 2842 19552 2848 19616
rect 2912 19552 2928 19616
rect 2992 19552 3008 19616
rect 3072 19552 3088 19616
rect 3152 19552 3158 19616
rect 2842 19551 3158 19552
rect 3790 19616 4106 19617
rect 3790 19552 3796 19616
rect 3860 19552 3876 19616
rect 3940 19552 3956 19616
rect 4020 19552 4036 19616
rect 4100 19552 4106 19616
rect 3790 19551 4106 19552
rect 0 19410 800 19440
rect 3233 19410 3299 19413
rect 0 19408 3299 19410
rect 0 19352 3238 19408
rect 3294 19352 3299 19408
rect 0 19350 3299 19352
rect 0 19320 800 19350
rect 3233 19347 3299 19350
rect 1420 19072 1736 19073
rect 1420 19008 1426 19072
rect 1490 19008 1506 19072
rect 1570 19008 1586 19072
rect 1650 19008 1666 19072
rect 1730 19008 1736 19072
rect 1420 19007 1736 19008
rect 2368 19072 2684 19073
rect 2368 19008 2374 19072
rect 2438 19008 2454 19072
rect 2518 19008 2534 19072
rect 2598 19008 2614 19072
rect 2678 19008 2684 19072
rect 2368 19007 2684 19008
rect 3316 19072 3632 19073
rect 3316 19008 3322 19072
rect 3386 19008 3402 19072
rect 3466 19008 3482 19072
rect 3546 19008 3562 19072
rect 3626 19008 3632 19072
rect 3316 19007 3632 19008
rect 4264 19072 4580 19073
rect 4264 19008 4270 19072
rect 4334 19008 4350 19072
rect 4414 19008 4430 19072
rect 4494 19008 4510 19072
rect 4574 19008 4580 19072
rect 4264 19007 4580 19008
rect 4153 18730 4219 18733
rect 5200 18730 6000 18760
rect 4153 18728 6000 18730
rect 4153 18672 4158 18728
rect 4214 18672 6000 18728
rect 4153 18670 6000 18672
rect 4153 18667 4219 18670
rect 5200 18640 6000 18670
rect 1894 18528 2210 18529
rect 1894 18464 1900 18528
rect 1964 18464 1980 18528
rect 2044 18464 2060 18528
rect 2124 18464 2140 18528
rect 2204 18464 2210 18528
rect 1894 18463 2210 18464
rect 2842 18528 3158 18529
rect 2842 18464 2848 18528
rect 2912 18464 2928 18528
rect 2992 18464 3008 18528
rect 3072 18464 3088 18528
rect 3152 18464 3158 18528
rect 2842 18463 3158 18464
rect 3790 18528 4106 18529
rect 3790 18464 3796 18528
rect 3860 18464 3876 18528
rect 3940 18464 3956 18528
rect 4020 18464 4036 18528
rect 4100 18464 4106 18528
rect 3790 18463 4106 18464
rect 1420 17984 1736 17985
rect 1420 17920 1426 17984
rect 1490 17920 1506 17984
rect 1570 17920 1586 17984
rect 1650 17920 1666 17984
rect 1730 17920 1736 17984
rect 1420 17919 1736 17920
rect 2368 17984 2684 17985
rect 2368 17920 2374 17984
rect 2438 17920 2454 17984
rect 2518 17920 2534 17984
rect 2598 17920 2614 17984
rect 2678 17920 2684 17984
rect 2368 17919 2684 17920
rect 3316 17984 3632 17985
rect 3316 17920 3322 17984
rect 3386 17920 3402 17984
rect 3466 17920 3482 17984
rect 3546 17920 3562 17984
rect 3626 17920 3632 17984
rect 3316 17919 3632 17920
rect 4264 17984 4580 17985
rect 4264 17920 4270 17984
rect 4334 17920 4350 17984
rect 4414 17920 4430 17984
rect 4494 17920 4510 17984
rect 4574 17920 4580 17984
rect 4264 17919 4580 17920
rect 1894 17440 2210 17441
rect 1894 17376 1900 17440
rect 1964 17376 1980 17440
rect 2044 17376 2060 17440
rect 2124 17376 2140 17440
rect 2204 17376 2210 17440
rect 1894 17375 2210 17376
rect 2842 17440 3158 17441
rect 2842 17376 2848 17440
rect 2912 17376 2928 17440
rect 2992 17376 3008 17440
rect 3072 17376 3088 17440
rect 3152 17376 3158 17440
rect 2842 17375 3158 17376
rect 3790 17440 4106 17441
rect 3790 17376 3796 17440
rect 3860 17376 3876 17440
rect 3940 17376 3956 17440
rect 4020 17376 4036 17440
rect 4100 17376 4106 17440
rect 3790 17375 4106 17376
rect 4153 17234 4219 17237
rect 5200 17234 6000 17264
rect 4153 17232 6000 17234
rect 4153 17176 4158 17232
rect 4214 17176 6000 17232
rect 4153 17174 6000 17176
rect 4153 17171 4219 17174
rect 5200 17144 6000 17174
rect 1420 16896 1736 16897
rect 1420 16832 1426 16896
rect 1490 16832 1506 16896
rect 1570 16832 1586 16896
rect 1650 16832 1666 16896
rect 1730 16832 1736 16896
rect 1420 16831 1736 16832
rect 2368 16896 2684 16897
rect 2368 16832 2374 16896
rect 2438 16832 2454 16896
rect 2518 16832 2534 16896
rect 2598 16832 2614 16896
rect 2678 16832 2684 16896
rect 2368 16831 2684 16832
rect 3316 16896 3632 16897
rect 3316 16832 3322 16896
rect 3386 16832 3402 16896
rect 3466 16832 3482 16896
rect 3546 16832 3562 16896
rect 3626 16832 3632 16896
rect 3316 16831 3632 16832
rect 4264 16896 4580 16897
rect 4264 16832 4270 16896
rect 4334 16832 4350 16896
rect 4414 16832 4430 16896
rect 4494 16832 4510 16896
rect 4574 16832 4580 16896
rect 4264 16831 4580 16832
rect 0 16418 800 16448
rect 1301 16418 1367 16421
rect 0 16416 1367 16418
rect 0 16360 1306 16416
rect 1362 16360 1367 16416
rect 0 16358 1367 16360
rect 0 16328 800 16358
rect 1301 16355 1367 16358
rect 1894 16352 2210 16353
rect 1894 16288 1900 16352
rect 1964 16288 1980 16352
rect 2044 16288 2060 16352
rect 2124 16288 2140 16352
rect 2204 16288 2210 16352
rect 1894 16287 2210 16288
rect 2842 16352 3158 16353
rect 2842 16288 2848 16352
rect 2912 16288 2928 16352
rect 2992 16288 3008 16352
rect 3072 16288 3088 16352
rect 3152 16288 3158 16352
rect 2842 16287 3158 16288
rect 3790 16352 4106 16353
rect 3790 16288 3796 16352
rect 3860 16288 3876 16352
rect 3940 16288 3956 16352
rect 4020 16288 4036 16352
rect 4100 16288 4106 16352
rect 3790 16287 4106 16288
rect 1420 15808 1736 15809
rect 1420 15744 1426 15808
rect 1490 15744 1506 15808
rect 1570 15744 1586 15808
rect 1650 15744 1666 15808
rect 1730 15744 1736 15808
rect 1420 15743 1736 15744
rect 2368 15808 2684 15809
rect 2368 15744 2374 15808
rect 2438 15744 2454 15808
rect 2518 15744 2534 15808
rect 2598 15744 2614 15808
rect 2678 15744 2684 15808
rect 2368 15743 2684 15744
rect 3316 15808 3632 15809
rect 3316 15744 3322 15808
rect 3386 15744 3402 15808
rect 3466 15744 3482 15808
rect 3546 15744 3562 15808
rect 3626 15744 3632 15808
rect 3316 15743 3632 15744
rect 4264 15808 4580 15809
rect 4264 15744 4270 15808
rect 4334 15744 4350 15808
rect 4414 15744 4430 15808
rect 4494 15744 4510 15808
rect 4574 15744 4580 15808
rect 4264 15743 4580 15744
rect 4705 15738 4771 15741
rect 5200 15738 6000 15768
rect 4705 15736 6000 15738
rect 4705 15680 4710 15736
rect 4766 15680 6000 15736
rect 4705 15678 6000 15680
rect 4705 15675 4771 15678
rect 5200 15648 6000 15678
rect 1894 15264 2210 15265
rect 1894 15200 1900 15264
rect 1964 15200 1980 15264
rect 2044 15200 2060 15264
rect 2124 15200 2140 15264
rect 2204 15200 2210 15264
rect 1894 15199 2210 15200
rect 2842 15264 3158 15265
rect 2842 15200 2848 15264
rect 2912 15200 2928 15264
rect 2992 15200 3008 15264
rect 3072 15200 3088 15264
rect 3152 15200 3158 15264
rect 2842 15199 3158 15200
rect 3790 15264 4106 15265
rect 3790 15200 3796 15264
rect 3860 15200 3876 15264
rect 3940 15200 3956 15264
rect 4020 15200 4036 15264
rect 4100 15200 4106 15264
rect 3790 15199 4106 15200
rect 1420 14720 1736 14721
rect 1420 14656 1426 14720
rect 1490 14656 1506 14720
rect 1570 14656 1586 14720
rect 1650 14656 1666 14720
rect 1730 14656 1736 14720
rect 1420 14655 1736 14656
rect 2368 14720 2684 14721
rect 2368 14656 2374 14720
rect 2438 14656 2454 14720
rect 2518 14656 2534 14720
rect 2598 14656 2614 14720
rect 2678 14656 2684 14720
rect 2368 14655 2684 14656
rect 3316 14720 3632 14721
rect 3316 14656 3322 14720
rect 3386 14656 3402 14720
rect 3466 14656 3482 14720
rect 3546 14656 3562 14720
rect 3626 14656 3632 14720
rect 3316 14655 3632 14656
rect 4264 14720 4580 14721
rect 4264 14656 4270 14720
rect 4334 14656 4350 14720
rect 4414 14656 4430 14720
rect 4494 14656 4510 14720
rect 4574 14656 4580 14720
rect 4264 14655 4580 14656
rect 4245 14242 4311 14245
rect 5200 14242 6000 14272
rect 4245 14240 6000 14242
rect 4245 14184 4250 14240
rect 4306 14184 6000 14240
rect 4245 14182 6000 14184
rect 4245 14179 4311 14182
rect 1894 14176 2210 14177
rect 1894 14112 1900 14176
rect 1964 14112 1980 14176
rect 2044 14112 2060 14176
rect 2124 14112 2140 14176
rect 2204 14112 2210 14176
rect 1894 14111 2210 14112
rect 2842 14176 3158 14177
rect 2842 14112 2848 14176
rect 2912 14112 2928 14176
rect 2992 14112 3008 14176
rect 3072 14112 3088 14176
rect 3152 14112 3158 14176
rect 2842 14111 3158 14112
rect 3790 14176 4106 14177
rect 3790 14112 3796 14176
rect 3860 14112 3876 14176
rect 3940 14112 3956 14176
rect 4020 14112 4036 14176
rect 4100 14112 4106 14176
rect 5200 14152 6000 14182
rect 3790 14111 4106 14112
rect 1420 13632 1736 13633
rect 1420 13568 1426 13632
rect 1490 13568 1506 13632
rect 1570 13568 1586 13632
rect 1650 13568 1666 13632
rect 1730 13568 1736 13632
rect 1420 13567 1736 13568
rect 2368 13632 2684 13633
rect 2368 13568 2374 13632
rect 2438 13568 2454 13632
rect 2518 13568 2534 13632
rect 2598 13568 2614 13632
rect 2678 13568 2684 13632
rect 2368 13567 2684 13568
rect 3316 13632 3632 13633
rect 3316 13568 3322 13632
rect 3386 13568 3402 13632
rect 3466 13568 3482 13632
rect 3546 13568 3562 13632
rect 3626 13568 3632 13632
rect 3316 13567 3632 13568
rect 4264 13632 4580 13633
rect 4264 13568 4270 13632
rect 4334 13568 4350 13632
rect 4414 13568 4430 13632
rect 4494 13568 4510 13632
rect 4574 13568 4580 13632
rect 4264 13567 4580 13568
rect 0 13426 800 13456
rect 1577 13426 1643 13429
rect 0 13424 1643 13426
rect 0 13368 1582 13424
rect 1638 13368 1643 13424
rect 0 13366 1643 13368
rect 0 13336 800 13366
rect 1577 13363 1643 13366
rect 1894 13088 2210 13089
rect 1894 13024 1900 13088
rect 1964 13024 1980 13088
rect 2044 13024 2060 13088
rect 2124 13024 2140 13088
rect 2204 13024 2210 13088
rect 1894 13023 2210 13024
rect 2842 13088 3158 13089
rect 2842 13024 2848 13088
rect 2912 13024 2928 13088
rect 2992 13024 3008 13088
rect 3072 13024 3088 13088
rect 3152 13024 3158 13088
rect 2842 13023 3158 13024
rect 3790 13088 4106 13089
rect 3790 13024 3796 13088
rect 3860 13024 3876 13088
rect 3940 13024 3956 13088
rect 4020 13024 4036 13088
rect 4100 13024 4106 13088
rect 3790 13023 4106 13024
rect 4061 12746 4127 12749
rect 5200 12746 6000 12776
rect 4061 12744 6000 12746
rect 4061 12688 4066 12744
rect 4122 12688 6000 12744
rect 4061 12686 6000 12688
rect 4061 12683 4127 12686
rect 5200 12656 6000 12686
rect 1420 12544 1736 12545
rect 1420 12480 1426 12544
rect 1490 12480 1506 12544
rect 1570 12480 1586 12544
rect 1650 12480 1666 12544
rect 1730 12480 1736 12544
rect 1420 12479 1736 12480
rect 2368 12544 2684 12545
rect 2368 12480 2374 12544
rect 2438 12480 2454 12544
rect 2518 12480 2534 12544
rect 2598 12480 2614 12544
rect 2678 12480 2684 12544
rect 2368 12479 2684 12480
rect 3316 12544 3632 12545
rect 3316 12480 3322 12544
rect 3386 12480 3402 12544
rect 3466 12480 3482 12544
rect 3546 12480 3562 12544
rect 3626 12480 3632 12544
rect 3316 12479 3632 12480
rect 4264 12544 4580 12545
rect 4264 12480 4270 12544
rect 4334 12480 4350 12544
rect 4414 12480 4430 12544
rect 4494 12480 4510 12544
rect 4574 12480 4580 12544
rect 4264 12479 4580 12480
rect 2313 12338 2379 12341
rect 2865 12338 2931 12341
rect 2313 12336 2931 12338
rect 2313 12280 2318 12336
rect 2374 12280 2870 12336
rect 2926 12280 2931 12336
rect 2313 12278 2931 12280
rect 2313 12275 2379 12278
rect 2865 12275 2931 12278
rect 1894 12000 2210 12001
rect 1894 11936 1900 12000
rect 1964 11936 1980 12000
rect 2044 11936 2060 12000
rect 2124 11936 2140 12000
rect 2204 11936 2210 12000
rect 1894 11935 2210 11936
rect 2842 12000 3158 12001
rect 2842 11936 2848 12000
rect 2912 11936 2928 12000
rect 2992 11936 3008 12000
rect 3072 11936 3088 12000
rect 3152 11936 3158 12000
rect 2842 11935 3158 11936
rect 3790 12000 4106 12001
rect 3790 11936 3796 12000
rect 3860 11936 3876 12000
rect 3940 11936 3956 12000
rect 4020 11936 4036 12000
rect 4100 11936 4106 12000
rect 3790 11935 4106 11936
rect 1420 11456 1736 11457
rect 1420 11392 1426 11456
rect 1490 11392 1506 11456
rect 1570 11392 1586 11456
rect 1650 11392 1666 11456
rect 1730 11392 1736 11456
rect 1420 11391 1736 11392
rect 2368 11456 2684 11457
rect 2368 11392 2374 11456
rect 2438 11392 2454 11456
rect 2518 11392 2534 11456
rect 2598 11392 2614 11456
rect 2678 11392 2684 11456
rect 2368 11391 2684 11392
rect 3316 11456 3632 11457
rect 3316 11392 3322 11456
rect 3386 11392 3402 11456
rect 3466 11392 3482 11456
rect 3546 11392 3562 11456
rect 3626 11392 3632 11456
rect 3316 11391 3632 11392
rect 4264 11456 4580 11457
rect 4264 11392 4270 11456
rect 4334 11392 4350 11456
rect 4414 11392 4430 11456
rect 4494 11392 4510 11456
rect 4574 11392 4580 11456
rect 4264 11391 4580 11392
rect 3417 11250 3483 11253
rect 5200 11250 6000 11280
rect 3417 11248 6000 11250
rect 3417 11192 3422 11248
rect 3478 11192 6000 11248
rect 3417 11190 6000 11192
rect 3417 11187 3483 11190
rect 5200 11160 6000 11190
rect 1894 10912 2210 10913
rect 1894 10848 1900 10912
rect 1964 10848 1980 10912
rect 2044 10848 2060 10912
rect 2124 10848 2140 10912
rect 2204 10848 2210 10912
rect 1894 10847 2210 10848
rect 2842 10912 3158 10913
rect 2842 10848 2848 10912
rect 2912 10848 2928 10912
rect 2992 10848 3008 10912
rect 3072 10848 3088 10912
rect 3152 10848 3158 10912
rect 2842 10847 3158 10848
rect 3790 10912 4106 10913
rect 3790 10848 3796 10912
rect 3860 10848 3876 10912
rect 3940 10848 3956 10912
rect 4020 10848 4036 10912
rect 4100 10848 4106 10912
rect 3790 10847 4106 10848
rect 1393 10570 1459 10573
rect 798 10568 1459 10570
rect 798 10512 1398 10568
rect 1454 10512 1459 10568
rect 798 10510 1459 10512
rect 798 10464 858 10510
rect 1393 10507 1459 10510
rect 3509 10570 3575 10573
rect 3509 10568 3802 10570
rect 3509 10512 3514 10568
rect 3570 10512 3802 10568
rect 3509 10510 3802 10512
rect 3509 10507 3575 10510
rect 0 10374 858 10464
rect 0 10344 800 10374
rect 1420 10368 1736 10369
rect 1420 10304 1426 10368
rect 1490 10304 1506 10368
rect 1570 10304 1586 10368
rect 1650 10304 1666 10368
rect 1730 10304 1736 10368
rect 1420 10303 1736 10304
rect 2368 10368 2684 10369
rect 2368 10304 2374 10368
rect 2438 10304 2454 10368
rect 2518 10304 2534 10368
rect 2598 10304 2614 10368
rect 2678 10304 2684 10368
rect 2368 10303 2684 10304
rect 3316 10368 3632 10369
rect 3316 10304 3322 10368
rect 3386 10304 3402 10368
rect 3466 10304 3482 10368
rect 3546 10304 3562 10368
rect 3626 10304 3632 10368
rect 3316 10303 3632 10304
rect 3601 10162 3667 10165
rect 3742 10162 3802 10510
rect 4264 10368 4580 10369
rect 4264 10304 4270 10368
rect 4334 10304 4350 10368
rect 4414 10304 4430 10368
rect 4494 10304 4510 10368
rect 4574 10304 4580 10368
rect 4264 10303 4580 10304
rect 3601 10160 3802 10162
rect 3601 10104 3606 10160
rect 3662 10104 3802 10160
rect 3601 10102 3802 10104
rect 3601 10099 3667 10102
rect 3233 10026 3299 10029
rect 3233 10024 4354 10026
rect 3233 9968 3238 10024
rect 3294 9968 4354 10024
rect 3233 9966 4354 9968
rect 3233 9963 3299 9966
rect 1894 9824 2210 9825
rect 1894 9760 1900 9824
rect 1964 9760 1980 9824
rect 2044 9760 2060 9824
rect 2124 9760 2140 9824
rect 2204 9760 2210 9824
rect 1894 9759 2210 9760
rect 2842 9824 3158 9825
rect 2842 9760 2848 9824
rect 2912 9760 2928 9824
rect 2992 9760 3008 9824
rect 3072 9760 3088 9824
rect 3152 9760 3158 9824
rect 2842 9759 3158 9760
rect 3790 9824 4106 9825
rect 3790 9760 3796 9824
rect 3860 9760 3876 9824
rect 3940 9760 3956 9824
rect 4020 9760 4036 9824
rect 4100 9760 4106 9824
rect 3790 9759 4106 9760
rect 4294 9754 4354 9966
rect 5200 9754 6000 9784
rect 4294 9694 6000 9754
rect 5200 9664 6000 9694
rect 1209 9618 1275 9621
rect 2773 9618 2839 9621
rect 1209 9616 2839 9618
rect 1209 9560 1214 9616
rect 1270 9560 2778 9616
rect 2834 9560 2839 9616
rect 1209 9558 2839 9560
rect 1209 9555 1275 9558
rect 2773 9555 2839 9558
rect 1420 9280 1736 9281
rect 1420 9216 1426 9280
rect 1490 9216 1506 9280
rect 1570 9216 1586 9280
rect 1650 9216 1666 9280
rect 1730 9216 1736 9280
rect 1420 9215 1736 9216
rect 2368 9280 2684 9281
rect 2368 9216 2374 9280
rect 2438 9216 2454 9280
rect 2518 9216 2534 9280
rect 2598 9216 2614 9280
rect 2678 9216 2684 9280
rect 2368 9215 2684 9216
rect 3316 9280 3632 9281
rect 3316 9216 3322 9280
rect 3386 9216 3402 9280
rect 3466 9216 3482 9280
rect 3546 9216 3562 9280
rect 3626 9216 3632 9280
rect 3316 9215 3632 9216
rect 4264 9280 4580 9281
rect 4264 9216 4270 9280
rect 4334 9216 4350 9280
rect 4414 9216 4430 9280
rect 4494 9216 4510 9280
rect 4574 9216 4580 9280
rect 4264 9215 4580 9216
rect 1894 8736 2210 8737
rect 1894 8672 1900 8736
rect 1964 8672 1980 8736
rect 2044 8672 2060 8736
rect 2124 8672 2140 8736
rect 2204 8672 2210 8736
rect 1894 8671 2210 8672
rect 2842 8736 3158 8737
rect 2842 8672 2848 8736
rect 2912 8672 2928 8736
rect 2992 8672 3008 8736
rect 3072 8672 3088 8736
rect 3152 8672 3158 8736
rect 2842 8671 3158 8672
rect 3790 8736 4106 8737
rect 3790 8672 3796 8736
rect 3860 8672 3876 8736
rect 3940 8672 3956 8736
rect 4020 8672 4036 8736
rect 4100 8672 4106 8736
rect 3790 8671 4106 8672
rect 4705 8258 4771 8261
rect 5200 8258 6000 8288
rect 4705 8256 6000 8258
rect 4705 8200 4710 8256
rect 4766 8200 6000 8256
rect 4705 8198 6000 8200
rect 4705 8195 4771 8198
rect 1420 8192 1736 8193
rect 1420 8128 1426 8192
rect 1490 8128 1506 8192
rect 1570 8128 1586 8192
rect 1650 8128 1666 8192
rect 1730 8128 1736 8192
rect 1420 8127 1736 8128
rect 2368 8192 2684 8193
rect 2368 8128 2374 8192
rect 2438 8128 2454 8192
rect 2518 8128 2534 8192
rect 2598 8128 2614 8192
rect 2678 8128 2684 8192
rect 2368 8127 2684 8128
rect 3316 8192 3632 8193
rect 3316 8128 3322 8192
rect 3386 8128 3402 8192
rect 3466 8128 3482 8192
rect 3546 8128 3562 8192
rect 3626 8128 3632 8192
rect 3316 8127 3632 8128
rect 4264 8192 4580 8193
rect 4264 8128 4270 8192
rect 4334 8128 4350 8192
rect 4414 8128 4430 8192
rect 4494 8128 4510 8192
rect 4574 8128 4580 8192
rect 5200 8168 6000 8198
rect 4264 8127 4580 8128
rect 1894 7648 2210 7649
rect 1894 7584 1900 7648
rect 1964 7584 1980 7648
rect 2044 7584 2060 7648
rect 2124 7584 2140 7648
rect 2204 7584 2210 7648
rect 1894 7583 2210 7584
rect 2842 7648 3158 7649
rect 2842 7584 2848 7648
rect 2912 7584 2928 7648
rect 2992 7584 3008 7648
rect 3072 7584 3088 7648
rect 3152 7584 3158 7648
rect 2842 7583 3158 7584
rect 3790 7648 4106 7649
rect 3790 7584 3796 7648
rect 3860 7584 3876 7648
rect 3940 7584 3956 7648
rect 4020 7584 4036 7648
rect 4100 7584 4106 7648
rect 3790 7583 4106 7584
rect 0 7442 800 7472
rect 1393 7442 1459 7445
rect 0 7440 1459 7442
rect 0 7384 1398 7440
rect 1454 7384 1459 7440
rect 0 7382 1459 7384
rect 0 7352 800 7382
rect 1393 7379 1459 7382
rect 1420 7104 1736 7105
rect 1420 7040 1426 7104
rect 1490 7040 1506 7104
rect 1570 7040 1586 7104
rect 1650 7040 1666 7104
rect 1730 7040 1736 7104
rect 1420 7039 1736 7040
rect 2368 7104 2684 7105
rect 2368 7040 2374 7104
rect 2438 7040 2454 7104
rect 2518 7040 2534 7104
rect 2598 7040 2614 7104
rect 2678 7040 2684 7104
rect 2368 7039 2684 7040
rect 3316 7104 3632 7105
rect 3316 7040 3322 7104
rect 3386 7040 3402 7104
rect 3466 7040 3482 7104
rect 3546 7040 3562 7104
rect 3626 7040 3632 7104
rect 3316 7039 3632 7040
rect 4264 7104 4580 7105
rect 4264 7040 4270 7104
rect 4334 7040 4350 7104
rect 4414 7040 4430 7104
rect 4494 7040 4510 7104
rect 4574 7040 4580 7104
rect 4264 7039 4580 7040
rect 3693 6762 3759 6765
rect 5200 6762 6000 6792
rect 3693 6760 6000 6762
rect 3693 6704 3698 6760
rect 3754 6704 6000 6760
rect 3693 6702 6000 6704
rect 3693 6699 3759 6702
rect 5200 6672 6000 6702
rect 1894 6560 2210 6561
rect 1894 6496 1900 6560
rect 1964 6496 1980 6560
rect 2044 6496 2060 6560
rect 2124 6496 2140 6560
rect 2204 6496 2210 6560
rect 1894 6495 2210 6496
rect 2842 6560 3158 6561
rect 2842 6496 2848 6560
rect 2912 6496 2928 6560
rect 2992 6496 3008 6560
rect 3072 6496 3088 6560
rect 3152 6496 3158 6560
rect 2842 6495 3158 6496
rect 3790 6560 4106 6561
rect 3790 6496 3796 6560
rect 3860 6496 3876 6560
rect 3940 6496 3956 6560
rect 4020 6496 4036 6560
rect 4100 6496 4106 6560
rect 3790 6495 4106 6496
rect 1420 6016 1736 6017
rect 1420 5952 1426 6016
rect 1490 5952 1506 6016
rect 1570 5952 1586 6016
rect 1650 5952 1666 6016
rect 1730 5952 1736 6016
rect 1420 5951 1736 5952
rect 2368 6016 2684 6017
rect 2368 5952 2374 6016
rect 2438 5952 2454 6016
rect 2518 5952 2534 6016
rect 2598 5952 2614 6016
rect 2678 5952 2684 6016
rect 2368 5951 2684 5952
rect 3316 6016 3632 6017
rect 3316 5952 3322 6016
rect 3386 5952 3402 6016
rect 3466 5952 3482 6016
rect 3546 5952 3562 6016
rect 3626 5952 3632 6016
rect 3316 5951 3632 5952
rect 4264 6016 4580 6017
rect 4264 5952 4270 6016
rect 4334 5952 4350 6016
rect 4414 5952 4430 6016
rect 4494 5952 4510 6016
rect 4574 5952 4580 6016
rect 4264 5951 4580 5952
rect 1894 5472 2210 5473
rect 1894 5408 1900 5472
rect 1964 5408 1980 5472
rect 2044 5408 2060 5472
rect 2124 5408 2140 5472
rect 2204 5408 2210 5472
rect 1894 5407 2210 5408
rect 2842 5472 3158 5473
rect 2842 5408 2848 5472
rect 2912 5408 2928 5472
rect 2992 5408 3008 5472
rect 3072 5408 3088 5472
rect 3152 5408 3158 5472
rect 2842 5407 3158 5408
rect 3790 5472 4106 5473
rect 3790 5408 3796 5472
rect 3860 5408 3876 5472
rect 3940 5408 3956 5472
rect 4020 5408 4036 5472
rect 4100 5408 4106 5472
rect 3790 5407 4106 5408
rect 4153 5266 4219 5269
rect 5200 5266 6000 5296
rect 4153 5264 6000 5266
rect 4153 5208 4158 5264
rect 4214 5208 6000 5264
rect 4153 5206 6000 5208
rect 4153 5203 4219 5206
rect 5200 5176 6000 5206
rect 1420 4928 1736 4929
rect 1420 4864 1426 4928
rect 1490 4864 1506 4928
rect 1570 4864 1586 4928
rect 1650 4864 1666 4928
rect 1730 4864 1736 4928
rect 1420 4863 1736 4864
rect 2368 4928 2684 4929
rect 2368 4864 2374 4928
rect 2438 4864 2454 4928
rect 2518 4864 2534 4928
rect 2598 4864 2614 4928
rect 2678 4864 2684 4928
rect 2368 4863 2684 4864
rect 3316 4928 3632 4929
rect 3316 4864 3322 4928
rect 3386 4864 3402 4928
rect 3466 4864 3482 4928
rect 3546 4864 3562 4928
rect 3626 4864 3632 4928
rect 3316 4863 3632 4864
rect 4264 4928 4580 4929
rect 4264 4864 4270 4928
rect 4334 4864 4350 4928
rect 4414 4864 4430 4928
rect 4494 4864 4510 4928
rect 4574 4864 4580 4928
rect 4264 4863 4580 4864
rect 0 4450 800 4480
rect 1393 4450 1459 4453
rect 0 4448 1459 4450
rect 0 4392 1398 4448
rect 1454 4392 1459 4448
rect 0 4390 1459 4392
rect 0 4360 800 4390
rect 1393 4387 1459 4390
rect 1894 4384 2210 4385
rect 1894 4320 1900 4384
rect 1964 4320 1980 4384
rect 2044 4320 2060 4384
rect 2124 4320 2140 4384
rect 2204 4320 2210 4384
rect 1894 4319 2210 4320
rect 2842 4384 3158 4385
rect 2842 4320 2848 4384
rect 2912 4320 2928 4384
rect 2992 4320 3008 4384
rect 3072 4320 3088 4384
rect 3152 4320 3158 4384
rect 2842 4319 3158 4320
rect 3790 4384 4106 4385
rect 3790 4320 3796 4384
rect 3860 4320 3876 4384
rect 3940 4320 3956 4384
rect 4020 4320 4036 4384
rect 4100 4320 4106 4384
rect 3790 4319 4106 4320
rect 3233 4042 3299 4045
rect 3233 4040 4722 4042
rect 3233 3984 3238 4040
rect 3294 3984 4722 4040
rect 3233 3982 4722 3984
rect 3233 3979 3299 3982
rect 1420 3840 1736 3841
rect 1420 3776 1426 3840
rect 1490 3776 1506 3840
rect 1570 3776 1586 3840
rect 1650 3776 1666 3840
rect 1730 3776 1736 3840
rect 1420 3775 1736 3776
rect 2368 3840 2684 3841
rect 2368 3776 2374 3840
rect 2438 3776 2454 3840
rect 2518 3776 2534 3840
rect 2598 3776 2614 3840
rect 2678 3776 2684 3840
rect 2368 3775 2684 3776
rect 3316 3840 3632 3841
rect 3316 3776 3322 3840
rect 3386 3776 3402 3840
rect 3466 3776 3482 3840
rect 3546 3776 3562 3840
rect 3626 3776 3632 3840
rect 3316 3775 3632 3776
rect 4264 3840 4580 3841
rect 4264 3776 4270 3840
rect 4334 3776 4350 3840
rect 4414 3776 4430 3840
rect 4494 3776 4510 3840
rect 4574 3776 4580 3840
rect 4264 3775 4580 3776
rect 4662 3770 4722 3982
rect 5200 3770 6000 3800
rect 4662 3710 6000 3770
rect 5200 3680 6000 3710
rect 1894 3296 2210 3297
rect 1894 3232 1900 3296
rect 1964 3232 1980 3296
rect 2044 3232 2060 3296
rect 2124 3232 2140 3296
rect 2204 3232 2210 3296
rect 1894 3231 2210 3232
rect 2842 3296 3158 3297
rect 2842 3232 2848 3296
rect 2912 3232 2928 3296
rect 2992 3232 3008 3296
rect 3072 3232 3088 3296
rect 3152 3232 3158 3296
rect 2842 3231 3158 3232
rect 3790 3296 4106 3297
rect 3790 3232 3796 3296
rect 3860 3232 3876 3296
rect 3940 3232 3956 3296
rect 4020 3232 4036 3296
rect 4100 3232 4106 3296
rect 3790 3231 4106 3232
rect 1420 2752 1736 2753
rect 1420 2688 1426 2752
rect 1490 2688 1506 2752
rect 1570 2688 1586 2752
rect 1650 2688 1666 2752
rect 1730 2688 1736 2752
rect 1420 2687 1736 2688
rect 2368 2752 2684 2753
rect 2368 2688 2374 2752
rect 2438 2688 2454 2752
rect 2518 2688 2534 2752
rect 2598 2688 2614 2752
rect 2678 2688 2684 2752
rect 2368 2687 2684 2688
rect 3316 2752 3632 2753
rect 3316 2688 3322 2752
rect 3386 2688 3402 2752
rect 3466 2688 3482 2752
rect 3546 2688 3562 2752
rect 3626 2688 3632 2752
rect 3316 2687 3632 2688
rect 4264 2752 4580 2753
rect 4264 2688 4270 2752
rect 4334 2688 4350 2752
rect 4414 2688 4430 2752
rect 4494 2688 4510 2752
rect 4574 2688 4580 2752
rect 4264 2687 4580 2688
rect 2221 2410 2287 2413
rect 2221 2408 4354 2410
rect 2221 2352 2226 2408
rect 2282 2352 4354 2408
rect 2221 2350 4354 2352
rect 2221 2347 2287 2350
rect 4294 2274 4354 2350
rect 5200 2274 6000 2304
rect 4294 2214 6000 2274
rect 1894 2208 2210 2209
rect 1894 2144 1900 2208
rect 1964 2144 1980 2208
rect 2044 2144 2060 2208
rect 2124 2144 2140 2208
rect 2204 2144 2210 2208
rect 1894 2143 2210 2144
rect 2842 2208 3158 2209
rect 2842 2144 2848 2208
rect 2912 2144 2928 2208
rect 2992 2144 3008 2208
rect 3072 2144 3088 2208
rect 3152 2144 3158 2208
rect 2842 2143 3158 2144
rect 3790 2208 4106 2209
rect 3790 2144 3796 2208
rect 3860 2144 3876 2208
rect 3940 2144 3956 2208
rect 4020 2144 4036 2208
rect 4100 2144 4106 2208
rect 5200 2184 6000 2214
rect 3790 2143 4106 2144
rect 1420 1664 1736 1665
rect 1420 1600 1426 1664
rect 1490 1600 1506 1664
rect 1570 1600 1586 1664
rect 1650 1600 1666 1664
rect 1730 1600 1736 1664
rect 1420 1599 1736 1600
rect 2368 1664 2684 1665
rect 2368 1600 2374 1664
rect 2438 1600 2454 1664
rect 2518 1600 2534 1664
rect 2598 1600 2614 1664
rect 2678 1600 2684 1664
rect 2368 1599 2684 1600
rect 3316 1664 3632 1665
rect 3316 1600 3322 1664
rect 3386 1600 3402 1664
rect 3466 1600 3482 1664
rect 3546 1600 3562 1664
rect 3626 1600 3632 1664
rect 3316 1599 3632 1600
rect 4264 1664 4580 1665
rect 4264 1600 4270 1664
rect 4334 1600 4350 1664
rect 4414 1600 4430 1664
rect 4494 1600 4510 1664
rect 4574 1600 4580 1664
rect 4264 1599 4580 1600
rect 0 1458 800 1488
rect 1761 1458 1827 1461
rect 0 1456 1827 1458
rect 0 1400 1766 1456
rect 1822 1400 1827 1456
rect 0 1398 1827 1400
rect 0 1368 800 1398
rect 1761 1395 1827 1398
rect 1894 1120 2210 1121
rect 1894 1056 1900 1120
rect 1964 1056 1980 1120
rect 2044 1056 2060 1120
rect 2124 1056 2140 1120
rect 2204 1056 2210 1120
rect 1894 1055 2210 1056
rect 2842 1120 3158 1121
rect 2842 1056 2848 1120
rect 2912 1056 2928 1120
rect 2992 1056 3008 1120
rect 3072 1056 3088 1120
rect 3152 1056 3158 1120
rect 2842 1055 3158 1056
rect 3790 1120 4106 1121
rect 3790 1056 3796 1120
rect 3860 1056 3876 1120
rect 3940 1056 3956 1120
rect 4020 1056 4036 1120
rect 4100 1056 4106 1120
rect 3790 1055 4106 1056
rect 4705 778 4771 781
rect 5200 778 6000 808
rect 4705 776 6000 778
rect 4705 720 4710 776
rect 4766 720 6000 776
rect 4705 718 6000 720
rect 4705 715 4771 718
rect 5200 688 6000 718
<< via3 >>
rect 1900 22876 1964 22880
rect 1900 22820 1904 22876
rect 1904 22820 1960 22876
rect 1960 22820 1964 22876
rect 1900 22816 1964 22820
rect 1980 22876 2044 22880
rect 1980 22820 1984 22876
rect 1984 22820 2040 22876
rect 2040 22820 2044 22876
rect 1980 22816 2044 22820
rect 2060 22876 2124 22880
rect 2060 22820 2064 22876
rect 2064 22820 2120 22876
rect 2120 22820 2124 22876
rect 2060 22816 2124 22820
rect 2140 22876 2204 22880
rect 2140 22820 2144 22876
rect 2144 22820 2200 22876
rect 2200 22820 2204 22876
rect 2140 22816 2204 22820
rect 2848 22876 2912 22880
rect 2848 22820 2852 22876
rect 2852 22820 2908 22876
rect 2908 22820 2912 22876
rect 2848 22816 2912 22820
rect 2928 22876 2992 22880
rect 2928 22820 2932 22876
rect 2932 22820 2988 22876
rect 2988 22820 2992 22876
rect 2928 22816 2992 22820
rect 3008 22876 3072 22880
rect 3008 22820 3012 22876
rect 3012 22820 3068 22876
rect 3068 22820 3072 22876
rect 3008 22816 3072 22820
rect 3088 22876 3152 22880
rect 3088 22820 3092 22876
rect 3092 22820 3148 22876
rect 3148 22820 3152 22876
rect 3088 22816 3152 22820
rect 3796 22876 3860 22880
rect 3796 22820 3800 22876
rect 3800 22820 3856 22876
rect 3856 22820 3860 22876
rect 3796 22816 3860 22820
rect 3876 22876 3940 22880
rect 3876 22820 3880 22876
rect 3880 22820 3936 22876
rect 3936 22820 3940 22876
rect 3876 22816 3940 22820
rect 3956 22876 4020 22880
rect 3956 22820 3960 22876
rect 3960 22820 4016 22876
rect 4016 22820 4020 22876
rect 3956 22816 4020 22820
rect 4036 22876 4100 22880
rect 4036 22820 4040 22876
rect 4040 22820 4096 22876
rect 4096 22820 4100 22876
rect 4036 22816 4100 22820
rect 1426 22332 1490 22336
rect 1426 22276 1430 22332
rect 1430 22276 1486 22332
rect 1486 22276 1490 22332
rect 1426 22272 1490 22276
rect 1506 22332 1570 22336
rect 1506 22276 1510 22332
rect 1510 22276 1566 22332
rect 1566 22276 1570 22332
rect 1506 22272 1570 22276
rect 1586 22332 1650 22336
rect 1586 22276 1590 22332
rect 1590 22276 1646 22332
rect 1646 22276 1650 22332
rect 1586 22272 1650 22276
rect 1666 22332 1730 22336
rect 1666 22276 1670 22332
rect 1670 22276 1726 22332
rect 1726 22276 1730 22332
rect 1666 22272 1730 22276
rect 2374 22332 2438 22336
rect 2374 22276 2378 22332
rect 2378 22276 2434 22332
rect 2434 22276 2438 22332
rect 2374 22272 2438 22276
rect 2454 22332 2518 22336
rect 2454 22276 2458 22332
rect 2458 22276 2514 22332
rect 2514 22276 2518 22332
rect 2454 22272 2518 22276
rect 2534 22332 2598 22336
rect 2534 22276 2538 22332
rect 2538 22276 2594 22332
rect 2594 22276 2598 22332
rect 2534 22272 2598 22276
rect 2614 22332 2678 22336
rect 2614 22276 2618 22332
rect 2618 22276 2674 22332
rect 2674 22276 2678 22332
rect 2614 22272 2678 22276
rect 3322 22332 3386 22336
rect 3322 22276 3326 22332
rect 3326 22276 3382 22332
rect 3382 22276 3386 22332
rect 3322 22272 3386 22276
rect 3402 22332 3466 22336
rect 3402 22276 3406 22332
rect 3406 22276 3462 22332
rect 3462 22276 3466 22332
rect 3402 22272 3466 22276
rect 3482 22332 3546 22336
rect 3482 22276 3486 22332
rect 3486 22276 3542 22332
rect 3542 22276 3546 22332
rect 3482 22272 3546 22276
rect 3562 22332 3626 22336
rect 3562 22276 3566 22332
rect 3566 22276 3622 22332
rect 3622 22276 3626 22332
rect 3562 22272 3626 22276
rect 4270 22332 4334 22336
rect 4270 22276 4274 22332
rect 4274 22276 4330 22332
rect 4330 22276 4334 22332
rect 4270 22272 4334 22276
rect 4350 22332 4414 22336
rect 4350 22276 4354 22332
rect 4354 22276 4410 22332
rect 4410 22276 4414 22332
rect 4350 22272 4414 22276
rect 4430 22332 4494 22336
rect 4430 22276 4434 22332
rect 4434 22276 4490 22332
rect 4490 22276 4494 22332
rect 4430 22272 4494 22276
rect 4510 22332 4574 22336
rect 4510 22276 4514 22332
rect 4514 22276 4570 22332
rect 4570 22276 4574 22332
rect 4510 22272 4574 22276
rect 1900 21788 1964 21792
rect 1900 21732 1904 21788
rect 1904 21732 1960 21788
rect 1960 21732 1964 21788
rect 1900 21728 1964 21732
rect 1980 21788 2044 21792
rect 1980 21732 1984 21788
rect 1984 21732 2040 21788
rect 2040 21732 2044 21788
rect 1980 21728 2044 21732
rect 2060 21788 2124 21792
rect 2060 21732 2064 21788
rect 2064 21732 2120 21788
rect 2120 21732 2124 21788
rect 2060 21728 2124 21732
rect 2140 21788 2204 21792
rect 2140 21732 2144 21788
rect 2144 21732 2200 21788
rect 2200 21732 2204 21788
rect 2140 21728 2204 21732
rect 2848 21788 2912 21792
rect 2848 21732 2852 21788
rect 2852 21732 2908 21788
rect 2908 21732 2912 21788
rect 2848 21728 2912 21732
rect 2928 21788 2992 21792
rect 2928 21732 2932 21788
rect 2932 21732 2988 21788
rect 2988 21732 2992 21788
rect 2928 21728 2992 21732
rect 3008 21788 3072 21792
rect 3008 21732 3012 21788
rect 3012 21732 3068 21788
rect 3068 21732 3072 21788
rect 3008 21728 3072 21732
rect 3088 21788 3152 21792
rect 3088 21732 3092 21788
rect 3092 21732 3148 21788
rect 3148 21732 3152 21788
rect 3088 21728 3152 21732
rect 3796 21788 3860 21792
rect 3796 21732 3800 21788
rect 3800 21732 3856 21788
rect 3856 21732 3860 21788
rect 3796 21728 3860 21732
rect 3876 21788 3940 21792
rect 3876 21732 3880 21788
rect 3880 21732 3936 21788
rect 3936 21732 3940 21788
rect 3876 21728 3940 21732
rect 3956 21788 4020 21792
rect 3956 21732 3960 21788
rect 3960 21732 4016 21788
rect 4016 21732 4020 21788
rect 3956 21728 4020 21732
rect 4036 21788 4100 21792
rect 4036 21732 4040 21788
rect 4040 21732 4096 21788
rect 4096 21732 4100 21788
rect 4036 21728 4100 21732
rect 1426 21244 1490 21248
rect 1426 21188 1430 21244
rect 1430 21188 1486 21244
rect 1486 21188 1490 21244
rect 1426 21184 1490 21188
rect 1506 21244 1570 21248
rect 1506 21188 1510 21244
rect 1510 21188 1566 21244
rect 1566 21188 1570 21244
rect 1506 21184 1570 21188
rect 1586 21244 1650 21248
rect 1586 21188 1590 21244
rect 1590 21188 1646 21244
rect 1646 21188 1650 21244
rect 1586 21184 1650 21188
rect 1666 21244 1730 21248
rect 1666 21188 1670 21244
rect 1670 21188 1726 21244
rect 1726 21188 1730 21244
rect 1666 21184 1730 21188
rect 2374 21244 2438 21248
rect 2374 21188 2378 21244
rect 2378 21188 2434 21244
rect 2434 21188 2438 21244
rect 2374 21184 2438 21188
rect 2454 21244 2518 21248
rect 2454 21188 2458 21244
rect 2458 21188 2514 21244
rect 2514 21188 2518 21244
rect 2454 21184 2518 21188
rect 2534 21244 2598 21248
rect 2534 21188 2538 21244
rect 2538 21188 2594 21244
rect 2594 21188 2598 21244
rect 2534 21184 2598 21188
rect 2614 21244 2678 21248
rect 2614 21188 2618 21244
rect 2618 21188 2674 21244
rect 2674 21188 2678 21244
rect 2614 21184 2678 21188
rect 3322 21244 3386 21248
rect 3322 21188 3326 21244
rect 3326 21188 3382 21244
rect 3382 21188 3386 21244
rect 3322 21184 3386 21188
rect 3402 21244 3466 21248
rect 3402 21188 3406 21244
rect 3406 21188 3462 21244
rect 3462 21188 3466 21244
rect 3402 21184 3466 21188
rect 3482 21244 3546 21248
rect 3482 21188 3486 21244
rect 3486 21188 3542 21244
rect 3542 21188 3546 21244
rect 3482 21184 3546 21188
rect 3562 21244 3626 21248
rect 3562 21188 3566 21244
rect 3566 21188 3622 21244
rect 3622 21188 3626 21244
rect 3562 21184 3626 21188
rect 4270 21244 4334 21248
rect 4270 21188 4274 21244
rect 4274 21188 4330 21244
rect 4330 21188 4334 21244
rect 4270 21184 4334 21188
rect 4350 21244 4414 21248
rect 4350 21188 4354 21244
rect 4354 21188 4410 21244
rect 4410 21188 4414 21244
rect 4350 21184 4414 21188
rect 4430 21244 4494 21248
rect 4430 21188 4434 21244
rect 4434 21188 4490 21244
rect 4490 21188 4494 21244
rect 4430 21184 4494 21188
rect 4510 21244 4574 21248
rect 4510 21188 4514 21244
rect 4514 21188 4570 21244
rect 4570 21188 4574 21244
rect 4510 21184 4574 21188
rect 1900 20700 1964 20704
rect 1900 20644 1904 20700
rect 1904 20644 1960 20700
rect 1960 20644 1964 20700
rect 1900 20640 1964 20644
rect 1980 20700 2044 20704
rect 1980 20644 1984 20700
rect 1984 20644 2040 20700
rect 2040 20644 2044 20700
rect 1980 20640 2044 20644
rect 2060 20700 2124 20704
rect 2060 20644 2064 20700
rect 2064 20644 2120 20700
rect 2120 20644 2124 20700
rect 2060 20640 2124 20644
rect 2140 20700 2204 20704
rect 2140 20644 2144 20700
rect 2144 20644 2200 20700
rect 2200 20644 2204 20700
rect 2140 20640 2204 20644
rect 2848 20700 2912 20704
rect 2848 20644 2852 20700
rect 2852 20644 2908 20700
rect 2908 20644 2912 20700
rect 2848 20640 2912 20644
rect 2928 20700 2992 20704
rect 2928 20644 2932 20700
rect 2932 20644 2988 20700
rect 2988 20644 2992 20700
rect 2928 20640 2992 20644
rect 3008 20700 3072 20704
rect 3008 20644 3012 20700
rect 3012 20644 3068 20700
rect 3068 20644 3072 20700
rect 3008 20640 3072 20644
rect 3088 20700 3152 20704
rect 3088 20644 3092 20700
rect 3092 20644 3148 20700
rect 3148 20644 3152 20700
rect 3088 20640 3152 20644
rect 3796 20700 3860 20704
rect 3796 20644 3800 20700
rect 3800 20644 3856 20700
rect 3856 20644 3860 20700
rect 3796 20640 3860 20644
rect 3876 20700 3940 20704
rect 3876 20644 3880 20700
rect 3880 20644 3936 20700
rect 3936 20644 3940 20700
rect 3876 20640 3940 20644
rect 3956 20700 4020 20704
rect 3956 20644 3960 20700
rect 3960 20644 4016 20700
rect 4016 20644 4020 20700
rect 3956 20640 4020 20644
rect 4036 20700 4100 20704
rect 4036 20644 4040 20700
rect 4040 20644 4096 20700
rect 4096 20644 4100 20700
rect 4036 20640 4100 20644
rect 1426 20156 1490 20160
rect 1426 20100 1430 20156
rect 1430 20100 1486 20156
rect 1486 20100 1490 20156
rect 1426 20096 1490 20100
rect 1506 20156 1570 20160
rect 1506 20100 1510 20156
rect 1510 20100 1566 20156
rect 1566 20100 1570 20156
rect 1506 20096 1570 20100
rect 1586 20156 1650 20160
rect 1586 20100 1590 20156
rect 1590 20100 1646 20156
rect 1646 20100 1650 20156
rect 1586 20096 1650 20100
rect 1666 20156 1730 20160
rect 1666 20100 1670 20156
rect 1670 20100 1726 20156
rect 1726 20100 1730 20156
rect 1666 20096 1730 20100
rect 2374 20156 2438 20160
rect 2374 20100 2378 20156
rect 2378 20100 2434 20156
rect 2434 20100 2438 20156
rect 2374 20096 2438 20100
rect 2454 20156 2518 20160
rect 2454 20100 2458 20156
rect 2458 20100 2514 20156
rect 2514 20100 2518 20156
rect 2454 20096 2518 20100
rect 2534 20156 2598 20160
rect 2534 20100 2538 20156
rect 2538 20100 2594 20156
rect 2594 20100 2598 20156
rect 2534 20096 2598 20100
rect 2614 20156 2678 20160
rect 2614 20100 2618 20156
rect 2618 20100 2674 20156
rect 2674 20100 2678 20156
rect 2614 20096 2678 20100
rect 3322 20156 3386 20160
rect 3322 20100 3326 20156
rect 3326 20100 3382 20156
rect 3382 20100 3386 20156
rect 3322 20096 3386 20100
rect 3402 20156 3466 20160
rect 3402 20100 3406 20156
rect 3406 20100 3462 20156
rect 3462 20100 3466 20156
rect 3402 20096 3466 20100
rect 3482 20156 3546 20160
rect 3482 20100 3486 20156
rect 3486 20100 3542 20156
rect 3542 20100 3546 20156
rect 3482 20096 3546 20100
rect 3562 20156 3626 20160
rect 3562 20100 3566 20156
rect 3566 20100 3622 20156
rect 3622 20100 3626 20156
rect 3562 20096 3626 20100
rect 4270 20156 4334 20160
rect 4270 20100 4274 20156
rect 4274 20100 4330 20156
rect 4330 20100 4334 20156
rect 4270 20096 4334 20100
rect 4350 20156 4414 20160
rect 4350 20100 4354 20156
rect 4354 20100 4410 20156
rect 4410 20100 4414 20156
rect 4350 20096 4414 20100
rect 4430 20156 4494 20160
rect 4430 20100 4434 20156
rect 4434 20100 4490 20156
rect 4490 20100 4494 20156
rect 4430 20096 4494 20100
rect 4510 20156 4574 20160
rect 4510 20100 4514 20156
rect 4514 20100 4570 20156
rect 4570 20100 4574 20156
rect 4510 20096 4574 20100
rect 1900 19612 1964 19616
rect 1900 19556 1904 19612
rect 1904 19556 1960 19612
rect 1960 19556 1964 19612
rect 1900 19552 1964 19556
rect 1980 19612 2044 19616
rect 1980 19556 1984 19612
rect 1984 19556 2040 19612
rect 2040 19556 2044 19612
rect 1980 19552 2044 19556
rect 2060 19612 2124 19616
rect 2060 19556 2064 19612
rect 2064 19556 2120 19612
rect 2120 19556 2124 19612
rect 2060 19552 2124 19556
rect 2140 19612 2204 19616
rect 2140 19556 2144 19612
rect 2144 19556 2200 19612
rect 2200 19556 2204 19612
rect 2140 19552 2204 19556
rect 2848 19612 2912 19616
rect 2848 19556 2852 19612
rect 2852 19556 2908 19612
rect 2908 19556 2912 19612
rect 2848 19552 2912 19556
rect 2928 19612 2992 19616
rect 2928 19556 2932 19612
rect 2932 19556 2988 19612
rect 2988 19556 2992 19612
rect 2928 19552 2992 19556
rect 3008 19612 3072 19616
rect 3008 19556 3012 19612
rect 3012 19556 3068 19612
rect 3068 19556 3072 19612
rect 3008 19552 3072 19556
rect 3088 19612 3152 19616
rect 3088 19556 3092 19612
rect 3092 19556 3148 19612
rect 3148 19556 3152 19612
rect 3088 19552 3152 19556
rect 3796 19612 3860 19616
rect 3796 19556 3800 19612
rect 3800 19556 3856 19612
rect 3856 19556 3860 19612
rect 3796 19552 3860 19556
rect 3876 19612 3940 19616
rect 3876 19556 3880 19612
rect 3880 19556 3936 19612
rect 3936 19556 3940 19612
rect 3876 19552 3940 19556
rect 3956 19612 4020 19616
rect 3956 19556 3960 19612
rect 3960 19556 4016 19612
rect 4016 19556 4020 19612
rect 3956 19552 4020 19556
rect 4036 19612 4100 19616
rect 4036 19556 4040 19612
rect 4040 19556 4096 19612
rect 4096 19556 4100 19612
rect 4036 19552 4100 19556
rect 1426 19068 1490 19072
rect 1426 19012 1430 19068
rect 1430 19012 1486 19068
rect 1486 19012 1490 19068
rect 1426 19008 1490 19012
rect 1506 19068 1570 19072
rect 1506 19012 1510 19068
rect 1510 19012 1566 19068
rect 1566 19012 1570 19068
rect 1506 19008 1570 19012
rect 1586 19068 1650 19072
rect 1586 19012 1590 19068
rect 1590 19012 1646 19068
rect 1646 19012 1650 19068
rect 1586 19008 1650 19012
rect 1666 19068 1730 19072
rect 1666 19012 1670 19068
rect 1670 19012 1726 19068
rect 1726 19012 1730 19068
rect 1666 19008 1730 19012
rect 2374 19068 2438 19072
rect 2374 19012 2378 19068
rect 2378 19012 2434 19068
rect 2434 19012 2438 19068
rect 2374 19008 2438 19012
rect 2454 19068 2518 19072
rect 2454 19012 2458 19068
rect 2458 19012 2514 19068
rect 2514 19012 2518 19068
rect 2454 19008 2518 19012
rect 2534 19068 2598 19072
rect 2534 19012 2538 19068
rect 2538 19012 2594 19068
rect 2594 19012 2598 19068
rect 2534 19008 2598 19012
rect 2614 19068 2678 19072
rect 2614 19012 2618 19068
rect 2618 19012 2674 19068
rect 2674 19012 2678 19068
rect 2614 19008 2678 19012
rect 3322 19068 3386 19072
rect 3322 19012 3326 19068
rect 3326 19012 3382 19068
rect 3382 19012 3386 19068
rect 3322 19008 3386 19012
rect 3402 19068 3466 19072
rect 3402 19012 3406 19068
rect 3406 19012 3462 19068
rect 3462 19012 3466 19068
rect 3402 19008 3466 19012
rect 3482 19068 3546 19072
rect 3482 19012 3486 19068
rect 3486 19012 3542 19068
rect 3542 19012 3546 19068
rect 3482 19008 3546 19012
rect 3562 19068 3626 19072
rect 3562 19012 3566 19068
rect 3566 19012 3622 19068
rect 3622 19012 3626 19068
rect 3562 19008 3626 19012
rect 4270 19068 4334 19072
rect 4270 19012 4274 19068
rect 4274 19012 4330 19068
rect 4330 19012 4334 19068
rect 4270 19008 4334 19012
rect 4350 19068 4414 19072
rect 4350 19012 4354 19068
rect 4354 19012 4410 19068
rect 4410 19012 4414 19068
rect 4350 19008 4414 19012
rect 4430 19068 4494 19072
rect 4430 19012 4434 19068
rect 4434 19012 4490 19068
rect 4490 19012 4494 19068
rect 4430 19008 4494 19012
rect 4510 19068 4574 19072
rect 4510 19012 4514 19068
rect 4514 19012 4570 19068
rect 4570 19012 4574 19068
rect 4510 19008 4574 19012
rect 1900 18524 1964 18528
rect 1900 18468 1904 18524
rect 1904 18468 1960 18524
rect 1960 18468 1964 18524
rect 1900 18464 1964 18468
rect 1980 18524 2044 18528
rect 1980 18468 1984 18524
rect 1984 18468 2040 18524
rect 2040 18468 2044 18524
rect 1980 18464 2044 18468
rect 2060 18524 2124 18528
rect 2060 18468 2064 18524
rect 2064 18468 2120 18524
rect 2120 18468 2124 18524
rect 2060 18464 2124 18468
rect 2140 18524 2204 18528
rect 2140 18468 2144 18524
rect 2144 18468 2200 18524
rect 2200 18468 2204 18524
rect 2140 18464 2204 18468
rect 2848 18524 2912 18528
rect 2848 18468 2852 18524
rect 2852 18468 2908 18524
rect 2908 18468 2912 18524
rect 2848 18464 2912 18468
rect 2928 18524 2992 18528
rect 2928 18468 2932 18524
rect 2932 18468 2988 18524
rect 2988 18468 2992 18524
rect 2928 18464 2992 18468
rect 3008 18524 3072 18528
rect 3008 18468 3012 18524
rect 3012 18468 3068 18524
rect 3068 18468 3072 18524
rect 3008 18464 3072 18468
rect 3088 18524 3152 18528
rect 3088 18468 3092 18524
rect 3092 18468 3148 18524
rect 3148 18468 3152 18524
rect 3088 18464 3152 18468
rect 3796 18524 3860 18528
rect 3796 18468 3800 18524
rect 3800 18468 3856 18524
rect 3856 18468 3860 18524
rect 3796 18464 3860 18468
rect 3876 18524 3940 18528
rect 3876 18468 3880 18524
rect 3880 18468 3936 18524
rect 3936 18468 3940 18524
rect 3876 18464 3940 18468
rect 3956 18524 4020 18528
rect 3956 18468 3960 18524
rect 3960 18468 4016 18524
rect 4016 18468 4020 18524
rect 3956 18464 4020 18468
rect 4036 18524 4100 18528
rect 4036 18468 4040 18524
rect 4040 18468 4096 18524
rect 4096 18468 4100 18524
rect 4036 18464 4100 18468
rect 1426 17980 1490 17984
rect 1426 17924 1430 17980
rect 1430 17924 1486 17980
rect 1486 17924 1490 17980
rect 1426 17920 1490 17924
rect 1506 17980 1570 17984
rect 1506 17924 1510 17980
rect 1510 17924 1566 17980
rect 1566 17924 1570 17980
rect 1506 17920 1570 17924
rect 1586 17980 1650 17984
rect 1586 17924 1590 17980
rect 1590 17924 1646 17980
rect 1646 17924 1650 17980
rect 1586 17920 1650 17924
rect 1666 17980 1730 17984
rect 1666 17924 1670 17980
rect 1670 17924 1726 17980
rect 1726 17924 1730 17980
rect 1666 17920 1730 17924
rect 2374 17980 2438 17984
rect 2374 17924 2378 17980
rect 2378 17924 2434 17980
rect 2434 17924 2438 17980
rect 2374 17920 2438 17924
rect 2454 17980 2518 17984
rect 2454 17924 2458 17980
rect 2458 17924 2514 17980
rect 2514 17924 2518 17980
rect 2454 17920 2518 17924
rect 2534 17980 2598 17984
rect 2534 17924 2538 17980
rect 2538 17924 2594 17980
rect 2594 17924 2598 17980
rect 2534 17920 2598 17924
rect 2614 17980 2678 17984
rect 2614 17924 2618 17980
rect 2618 17924 2674 17980
rect 2674 17924 2678 17980
rect 2614 17920 2678 17924
rect 3322 17980 3386 17984
rect 3322 17924 3326 17980
rect 3326 17924 3382 17980
rect 3382 17924 3386 17980
rect 3322 17920 3386 17924
rect 3402 17980 3466 17984
rect 3402 17924 3406 17980
rect 3406 17924 3462 17980
rect 3462 17924 3466 17980
rect 3402 17920 3466 17924
rect 3482 17980 3546 17984
rect 3482 17924 3486 17980
rect 3486 17924 3542 17980
rect 3542 17924 3546 17980
rect 3482 17920 3546 17924
rect 3562 17980 3626 17984
rect 3562 17924 3566 17980
rect 3566 17924 3622 17980
rect 3622 17924 3626 17980
rect 3562 17920 3626 17924
rect 4270 17980 4334 17984
rect 4270 17924 4274 17980
rect 4274 17924 4330 17980
rect 4330 17924 4334 17980
rect 4270 17920 4334 17924
rect 4350 17980 4414 17984
rect 4350 17924 4354 17980
rect 4354 17924 4410 17980
rect 4410 17924 4414 17980
rect 4350 17920 4414 17924
rect 4430 17980 4494 17984
rect 4430 17924 4434 17980
rect 4434 17924 4490 17980
rect 4490 17924 4494 17980
rect 4430 17920 4494 17924
rect 4510 17980 4574 17984
rect 4510 17924 4514 17980
rect 4514 17924 4570 17980
rect 4570 17924 4574 17980
rect 4510 17920 4574 17924
rect 1900 17436 1964 17440
rect 1900 17380 1904 17436
rect 1904 17380 1960 17436
rect 1960 17380 1964 17436
rect 1900 17376 1964 17380
rect 1980 17436 2044 17440
rect 1980 17380 1984 17436
rect 1984 17380 2040 17436
rect 2040 17380 2044 17436
rect 1980 17376 2044 17380
rect 2060 17436 2124 17440
rect 2060 17380 2064 17436
rect 2064 17380 2120 17436
rect 2120 17380 2124 17436
rect 2060 17376 2124 17380
rect 2140 17436 2204 17440
rect 2140 17380 2144 17436
rect 2144 17380 2200 17436
rect 2200 17380 2204 17436
rect 2140 17376 2204 17380
rect 2848 17436 2912 17440
rect 2848 17380 2852 17436
rect 2852 17380 2908 17436
rect 2908 17380 2912 17436
rect 2848 17376 2912 17380
rect 2928 17436 2992 17440
rect 2928 17380 2932 17436
rect 2932 17380 2988 17436
rect 2988 17380 2992 17436
rect 2928 17376 2992 17380
rect 3008 17436 3072 17440
rect 3008 17380 3012 17436
rect 3012 17380 3068 17436
rect 3068 17380 3072 17436
rect 3008 17376 3072 17380
rect 3088 17436 3152 17440
rect 3088 17380 3092 17436
rect 3092 17380 3148 17436
rect 3148 17380 3152 17436
rect 3088 17376 3152 17380
rect 3796 17436 3860 17440
rect 3796 17380 3800 17436
rect 3800 17380 3856 17436
rect 3856 17380 3860 17436
rect 3796 17376 3860 17380
rect 3876 17436 3940 17440
rect 3876 17380 3880 17436
rect 3880 17380 3936 17436
rect 3936 17380 3940 17436
rect 3876 17376 3940 17380
rect 3956 17436 4020 17440
rect 3956 17380 3960 17436
rect 3960 17380 4016 17436
rect 4016 17380 4020 17436
rect 3956 17376 4020 17380
rect 4036 17436 4100 17440
rect 4036 17380 4040 17436
rect 4040 17380 4096 17436
rect 4096 17380 4100 17436
rect 4036 17376 4100 17380
rect 1426 16892 1490 16896
rect 1426 16836 1430 16892
rect 1430 16836 1486 16892
rect 1486 16836 1490 16892
rect 1426 16832 1490 16836
rect 1506 16892 1570 16896
rect 1506 16836 1510 16892
rect 1510 16836 1566 16892
rect 1566 16836 1570 16892
rect 1506 16832 1570 16836
rect 1586 16892 1650 16896
rect 1586 16836 1590 16892
rect 1590 16836 1646 16892
rect 1646 16836 1650 16892
rect 1586 16832 1650 16836
rect 1666 16892 1730 16896
rect 1666 16836 1670 16892
rect 1670 16836 1726 16892
rect 1726 16836 1730 16892
rect 1666 16832 1730 16836
rect 2374 16892 2438 16896
rect 2374 16836 2378 16892
rect 2378 16836 2434 16892
rect 2434 16836 2438 16892
rect 2374 16832 2438 16836
rect 2454 16892 2518 16896
rect 2454 16836 2458 16892
rect 2458 16836 2514 16892
rect 2514 16836 2518 16892
rect 2454 16832 2518 16836
rect 2534 16892 2598 16896
rect 2534 16836 2538 16892
rect 2538 16836 2594 16892
rect 2594 16836 2598 16892
rect 2534 16832 2598 16836
rect 2614 16892 2678 16896
rect 2614 16836 2618 16892
rect 2618 16836 2674 16892
rect 2674 16836 2678 16892
rect 2614 16832 2678 16836
rect 3322 16892 3386 16896
rect 3322 16836 3326 16892
rect 3326 16836 3382 16892
rect 3382 16836 3386 16892
rect 3322 16832 3386 16836
rect 3402 16892 3466 16896
rect 3402 16836 3406 16892
rect 3406 16836 3462 16892
rect 3462 16836 3466 16892
rect 3402 16832 3466 16836
rect 3482 16892 3546 16896
rect 3482 16836 3486 16892
rect 3486 16836 3542 16892
rect 3542 16836 3546 16892
rect 3482 16832 3546 16836
rect 3562 16892 3626 16896
rect 3562 16836 3566 16892
rect 3566 16836 3622 16892
rect 3622 16836 3626 16892
rect 3562 16832 3626 16836
rect 4270 16892 4334 16896
rect 4270 16836 4274 16892
rect 4274 16836 4330 16892
rect 4330 16836 4334 16892
rect 4270 16832 4334 16836
rect 4350 16892 4414 16896
rect 4350 16836 4354 16892
rect 4354 16836 4410 16892
rect 4410 16836 4414 16892
rect 4350 16832 4414 16836
rect 4430 16892 4494 16896
rect 4430 16836 4434 16892
rect 4434 16836 4490 16892
rect 4490 16836 4494 16892
rect 4430 16832 4494 16836
rect 4510 16892 4574 16896
rect 4510 16836 4514 16892
rect 4514 16836 4570 16892
rect 4570 16836 4574 16892
rect 4510 16832 4574 16836
rect 1900 16348 1964 16352
rect 1900 16292 1904 16348
rect 1904 16292 1960 16348
rect 1960 16292 1964 16348
rect 1900 16288 1964 16292
rect 1980 16348 2044 16352
rect 1980 16292 1984 16348
rect 1984 16292 2040 16348
rect 2040 16292 2044 16348
rect 1980 16288 2044 16292
rect 2060 16348 2124 16352
rect 2060 16292 2064 16348
rect 2064 16292 2120 16348
rect 2120 16292 2124 16348
rect 2060 16288 2124 16292
rect 2140 16348 2204 16352
rect 2140 16292 2144 16348
rect 2144 16292 2200 16348
rect 2200 16292 2204 16348
rect 2140 16288 2204 16292
rect 2848 16348 2912 16352
rect 2848 16292 2852 16348
rect 2852 16292 2908 16348
rect 2908 16292 2912 16348
rect 2848 16288 2912 16292
rect 2928 16348 2992 16352
rect 2928 16292 2932 16348
rect 2932 16292 2988 16348
rect 2988 16292 2992 16348
rect 2928 16288 2992 16292
rect 3008 16348 3072 16352
rect 3008 16292 3012 16348
rect 3012 16292 3068 16348
rect 3068 16292 3072 16348
rect 3008 16288 3072 16292
rect 3088 16348 3152 16352
rect 3088 16292 3092 16348
rect 3092 16292 3148 16348
rect 3148 16292 3152 16348
rect 3088 16288 3152 16292
rect 3796 16348 3860 16352
rect 3796 16292 3800 16348
rect 3800 16292 3856 16348
rect 3856 16292 3860 16348
rect 3796 16288 3860 16292
rect 3876 16348 3940 16352
rect 3876 16292 3880 16348
rect 3880 16292 3936 16348
rect 3936 16292 3940 16348
rect 3876 16288 3940 16292
rect 3956 16348 4020 16352
rect 3956 16292 3960 16348
rect 3960 16292 4016 16348
rect 4016 16292 4020 16348
rect 3956 16288 4020 16292
rect 4036 16348 4100 16352
rect 4036 16292 4040 16348
rect 4040 16292 4096 16348
rect 4096 16292 4100 16348
rect 4036 16288 4100 16292
rect 1426 15804 1490 15808
rect 1426 15748 1430 15804
rect 1430 15748 1486 15804
rect 1486 15748 1490 15804
rect 1426 15744 1490 15748
rect 1506 15804 1570 15808
rect 1506 15748 1510 15804
rect 1510 15748 1566 15804
rect 1566 15748 1570 15804
rect 1506 15744 1570 15748
rect 1586 15804 1650 15808
rect 1586 15748 1590 15804
rect 1590 15748 1646 15804
rect 1646 15748 1650 15804
rect 1586 15744 1650 15748
rect 1666 15804 1730 15808
rect 1666 15748 1670 15804
rect 1670 15748 1726 15804
rect 1726 15748 1730 15804
rect 1666 15744 1730 15748
rect 2374 15804 2438 15808
rect 2374 15748 2378 15804
rect 2378 15748 2434 15804
rect 2434 15748 2438 15804
rect 2374 15744 2438 15748
rect 2454 15804 2518 15808
rect 2454 15748 2458 15804
rect 2458 15748 2514 15804
rect 2514 15748 2518 15804
rect 2454 15744 2518 15748
rect 2534 15804 2598 15808
rect 2534 15748 2538 15804
rect 2538 15748 2594 15804
rect 2594 15748 2598 15804
rect 2534 15744 2598 15748
rect 2614 15804 2678 15808
rect 2614 15748 2618 15804
rect 2618 15748 2674 15804
rect 2674 15748 2678 15804
rect 2614 15744 2678 15748
rect 3322 15804 3386 15808
rect 3322 15748 3326 15804
rect 3326 15748 3382 15804
rect 3382 15748 3386 15804
rect 3322 15744 3386 15748
rect 3402 15804 3466 15808
rect 3402 15748 3406 15804
rect 3406 15748 3462 15804
rect 3462 15748 3466 15804
rect 3402 15744 3466 15748
rect 3482 15804 3546 15808
rect 3482 15748 3486 15804
rect 3486 15748 3542 15804
rect 3542 15748 3546 15804
rect 3482 15744 3546 15748
rect 3562 15804 3626 15808
rect 3562 15748 3566 15804
rect 3566 15748 3622 15804
rect 3622 15748 3626 15804
rect 3562 15744 3626 15748
rect 4270 15804 4334 15808
rect 4270 15748 4274 15804
rect 4274 15748 4330 15804
rect 4330 15748 4334 15804
rect 4270 15744 4334 15748
rect 4350 15804 4414 15808
rect 4350 15748 4354 15804
rect 4354 15748 4410 15804
rect 4410 15748 4414 15804
rect 4350 15744 4414 15748
rect 4430 15804 4494 15808
rect 4430 15748 4434 15804
rect 4434 15748 4490 15804
rect 4490 15748 4494 15804
rect 4430 15744 4494 15748
rect 4510 15804 4574 15808
rect 4510 15748 4514 15804
rect 4514 15748 4570 15804
rect 4570 15748 4574 15804
rect 4510 15744 4574 15748
rect 1900 15260 1964 15264
rect 1900 15204 1904 15260
rect 1904 15204 1960 15260
rect 1960 15204 1964 15260
rect 1900 15200 1964 15204
rect 1980 15260 2044 15264
rect 1980 15204 1984 15260
rect 1984 15204 2040 15260
rect 2040 15204 2044 15260
rect 1980 15200 2044 15204
rect 2060 15260 2124 15264
rect 2060 15204 2064 15260
rect 2064 15204 2120 15260
rect 2120 15204 2124 15260
rect 2060 15200 2124 15204
rect 2140 15260 2204 15264
rect 2140 15204 2144 15260
rect 2144 15204 2200 15260
rect 2200 15204 2204 15260
rect 2140 15200 2204 15204
rect 2848 15260 2912 15264
rect 2848 15204 2852 15260
rect 2852 15204 2908 15260
rect 2908 15204 2912 15260
rect 2848 15200 2912 15204
rect 2928 15260 2992 15264
rect 2928 15204 2932 15260
rect 2932 15204 2988 15260
rect 2988 15204 2992 15260
rect 2928 15200 2992 15204
rect 3008 15260 3072 15264
rect 3008 15204 3012 15260
rect 3012 15204 3068 15260
rect 3068 15204 3072 15260
rect 3008 15200 3072 15204
rect 3088 15260 3152 15264
rect 3088 15204 3092 15260
rect 3092 15204 3148 15260
rect 3148 15204 3152 15260
rect 3088 15200 3152 15204
rect 3796 15260 3860 15264
rect 3796 15204 3800 15260
rect 3800 15204 3856 15260
rect 3856 15204 3860 15260
rect 3796 15200 3860 15204
rect 3876 15260 3940 15264
rect 3876 15204 3880 15260
rect 3880 15204 3936 15260
rect 3936 15204 3940 15260
rect 3876 15200 3940 15204
rect 3956 15260 4020 15264
rect 3956 15204 3960 15260
rect 3960 15204 4016 15260
rect 4016 15204 4020 15260
rect 3956 15200 4020 15204
rect 4036 15260 4100 15264
rect 4036 15204 4040 15260
rect 4040 15204 4096 15260
rect 4096 15204 4100 15260
rect 4036 15200 4100 15204
rect 1426 14716 1490 14720
rect 1426 14660 1430 14716
rect 1430 14660 1486 14716
rect 1486 14660 1490 14716
rect 1426 14656 1490 14660
rect 1506 14716 1570 14720
rect 1506 14660 1510 14716
rect 1510 14660 1566 14716
rect 1566 14660 1570 14716
rect 1506 14656 1570 14660
rect 1586 14716 1650 14720
rect 1586 14660 1590 14716
rect 1590 14660 1646 14716
rect 1646 14660 1650 14716
rect 1586 14656 1650 14660
rect 1666 14716 1730 14720
rect 1666 14660 1670 14716
rect 1670 14660 1726 14716
rect 1726 14660 1730 14716
rect 1666 14656 1730 14660
rect 2374 14716 2438 14720
rect 2374 14660 2378 14716
rect 2378 14660 2434 14716
rect 2434 14660 2438 14716
rect 2374 14656 2438 14660
rect 2454 14716 2518 14720
rect 2454 14660 2458 14716
rect 2458 14660 2514 14716
rect 2514 14660 2518 14716
rect 2454 14656 2518 14660
rect 2534 14716 2598 14720
rect 2534 14660 2538 14716
rect 2538 14660 2594 14716
rect 2594 14660 2598 14716
rect 2534 14656 2598 14660
rect 2614 14716 2678 14720
rect 2614 14660 2618 14716
rect 2618 14660 2674 14716
rect 2674 14660 2678 14716
rect 2614 14656 2678 14660
rect 3322 14716 3386 14720
rect 3322 14660 3326 14716
rect 3326 14660 3382 14716
rect 3382 14660 3386 14716
rect 3322 14656 3386 14660
rect 3402 14716 3466 14720
rect 3402 14660 3406 14716
rect 3406 14660 3462 14716
rect 3462 14660 3466 14716
rect 3402 14656 3466 14660
rect 3482 14716 3546 14720
rect 3482 14660 3486 14716
rect 3486 14660 3542 14716
rect 3542 14660 3546 14716
rect 3482 14656 3546 14660
rect 3562 14716 3626 14720
rect 3562 14660 3566 14716
rect 3566 14660 3622 14716
rect 3622 14660 3626 14716
rect 3562 14656 3626 14660
rect 4270 14716 4334 14720
rect 4270 14660 4274 14716
rect 4274 14660 4330 14716
rect 4330 14660 4334 14716
rect 4270 14656 4334 14660
rect 4350 14716 4414 14720
rect 4350 14660 4354 14716
rect 4354 14660 4410 14716
rect 4410 14660 4414 14716
rect 4350 14656 4414 14660
rect 4430 14716 4494 14720
rect 4430 14660 4434 14716
rect 4434 14660 4490 14716
rect 4490 14660 4494 14716
rect 4430 14656 4494 14660
rect 4510 14716 4574 14720
rect 4510 14660 4514 14716
rect 4514 14660 4570 14716
rect 4570 14660 4574 14716
rect 4510 14656 4574 14660
rect 1900 14172 1964 14176
rect 1900 14116 1904 14172
rect 1904 14116 1960 14172
rect 1960 14116 1964 14172
rect 1900 14112 1964 14116
rect 1980 14172 2044 14176
rect 1980 14116 1984 14172
rect 1984 14116 2040 14172
rect 2040 14116 2044 14172
rect 1980 14112 2044 14116
rect 2060 14172 2124 14176
rect 2060 14116 2064 14172
rect 2064 14116 2120 14172
rect 2120 14116 2124 14172
rect 2060 14112 2124 14116
rect 2140 14172 2204 14176
rect 2140 14116 2144 14172
rect 2144 14116 2200 14172
rect 2200 14116 2204 14172
rect 2140 14112 2204 14116
rect 2848 14172 2912 14176
rect 2848 14116 2852 14172
rect 2852 14116 2908 14172
rect 2908 14116 2912 14172
rect 2848 14112 2912 14116
rect 2928 14172 2992 14176
rect 2928 14116 2932 14172
rect 2932 14116 2988 14172
rect 2988 14116 2992 14172
rect 2928 14112 2992 14116
rect 3008 14172 3072 14176
rect 3008 14116 3012 14172
rect 3012 14116 3068 14172
rect 3068 14116 3072 14172
rect 3008 14112 3072 14116
rect 3088 14172 3152 14176
rect 3088 14116 3092 14172
rect 3092 14116 3148 14172
rect 3148 14116 3152 14172
rect 3088 14112 3152 14116
rect 3796 14172 3860 14176
rect 3796 14116 3800 14172
rect 3800 14116 3856 14172
rect 3856 14116 3860 14172
rect 3796 14112 3860 14116
rect 3876 14172 3940 14176
rect 3876 14116 3880 14172
rect 3880 14116 3936 14172
rect 3936 14116 3940 14172
rect 3876 14112 3940 14116
rect 3956 14172 4020 14176
rect 3956 14116 3960 14172
rect 3960 14116 4016 14172
rect 4016 14116 4020 14172
rect 3956 14112 4020 14116
rect 4036 14172 4100 14176
rect 4036 14116 4040 14172
rect 4040 14116 4096 14172
rect 4096 14116 4100 14172
rect 4036 14112 4100 14116
rect 1426 13628 1490 13632
rect 1426 13572 1430 13628
rect 1430 13572 1486 13628
rect 1486 13572 1490 13628
rect 1426 13568 1490 13572
rect 1506 13628 1570 13632
rect 1506 13572 1510 13628
rect 1510 13572 1566 13628
rect 1566 13572 1570 13628
rect 1506 13568 1570 13572
rect 1586 13628 1650 13632
rect 1586 13572 1590 13628
rect 1590 13572 1646 13628
rect 1646 13572 1650 13628
rect 1586 13568 1650 13572
rect 1666 13628 1730 13632
rect 1666 13572 1670 13628
rect 1670 13572 1726 13628
rect 1726 13572 1730 13628
rect 1666 13568 1730 13572
rect 2374 13628 2438 13632
rect 2374 13572 2378 13628
rect 2378 13572 2434 13628
rect 2434 13572 2438 13628
rect 2374 13568 2438 13572
rect 2454 13628 2518 13632
rect 2454 13572 2458 13628
rect 2458 13572 2514 13628
rect 2514 13572 2518 13628
rect 2454 13568 2518 13572
rect 2534 13628 2598 13632
rect 2534 13572 2538 13628
rect 2538 13572 2594 13628
rect 2594 13572 2598 13628
rect 2534 13568 2598 13572
rect 2614 13628 2678 13632
rect 2614 13572 2618 13628
rect 2618 13572 2674 13628
rect 2674 13572 2678 13628
rect 2614 13568 2678 13572
rect 3322 13628 3386 13632
rect 3322 13572 3326 13628
rect 3326 13572 3382 13628
rect 3382 13572 3386 13628
rect 3322 13568 3386 13572
rect 3402 13628 3466 13632
rect 3402 13572 3406 13628
rect 3406 13572 3462 13628
rect 3462 13572 3466 13628
rect 3402 13568 3466 13572
rect 3482 13628 3546 13632
rect 3482 13572 3486 13628
rect 3486 13572 3542 13628
rect 3542 13572 3546 13628
rect 3482 13568 3546 13572
rect 3562 13628 3626 13632
rect 3562 13572 3566 13628
rect 3566 13572 3622 13628
rect 3622 13572 3626 13628
rect 3562 13568 3626 13572
rect 4270 13628 4334 13632
rect 4270 13572 4274 13628
rect 4274 13572 4330 13628
rect 4330 13572 4334 13628
rect 4270 13568 4334 13572
rect 4350 13628 4414 13632
rect 4350 13572 4354 13628
rect 4354 13572 4410 13628
rect 4410 13572 4414 13628
rect 4350 13568 4414 13572
rect 4430 13628 4494 13632
rect 4430 13572 4434 13628
rect 4434 13572 4490 13628
rect 4490 13572 4494 13628
rect 4430 13568 4494 13572
rect 4510 13628 4574 13632
rect 4510 13572 4514 13628
rect 4514 13572 4570 13628
rect 4570 13572 4574 13628
rect 4510 13568 4574 13572
rect 1900 13084 1964 13088
rect 1900 13028 1904 13084
rect 1904 13028 1960 13084
rect 1960 13028 1964 13084
rect 1900 13024 1964 13028
rect 1980 13084 2044 13088
rect 1980 13028 1984 13084
rect 1984 13028 2040 13084
rect 2040 13028 2044 13084
rect 1980 13024 2044 13028
rect 2060 13084 2124 13088
rect 2060 13028 2064 13084
rect 2064 13028 2120 13084
rect 2120 13028 2124 13084
rect 2060 13024 2124 13028
rect 2140 13084 2204 13088
rect 2140 13028 2144 13084
rect 2144 13028 2200 13084
rect 2200 13028 2204 13084
rect 2140 13024 2204 13028
rect 2848 13084 2912 13088
rect 2848 13028 2852 13084
rect 2852 13028 2908 13084
rect 2908 13028 2912 13084
rect 2848 13024 2912 13028
rect 2928 13084 2992 13088
rect 2928 13028 2932 13084
rect 2932 13028 2988 13084
rect 2988 13028 2992 13084
rect 2928 13024 2992 13028
rect 3008 13084 3072 13088
rect 3008 13028 3012 13084
rect 3012 13028 3068 13084
rect 3068 13028 3072 13084
rect 3008 13024 3072 13028
rect 3088 13084 3152 13088
rect 3088 13028 3092 13084
rect 3092 13028 3148 13084
rect 3148 13028 3152 13084
rect 3088 13024 3152 13028
rect 3796 13084 3860 13088
rect 3796 13028 3800 13084
rect 3800 13028 3856 13084
rect 3856 13028 3860 13084
rect 3796 13024 3860 13028
rect 3876 13084 3940 13088
rect 3876 13028 3880 13084
rect 3880 13028 3936 13084
rect 3936 13028 3940 13084
rect 3876 13024 3940 13028
rect 3956 13084 4020 13088
rect 3956 13028 3960 13084
rect 3960 13028 4016 13084
rect 4016 13028 4020 13084
rect 3956 13024 4020 13028
rect 4036 13084 4100 13088
rect 4036 13028 4040 13084
rect 4040 13028 4096 13084
rect 4096 13028 4100 13084
rect 4036 13024 4100 13028
rect 1426 12540 1490 12544
rect 1426 12484 1430 12540
rect 1430 12484 1486 12540
rect 1486 12484 1490 12540
rect 1426 12480 1490 12484
rect 1506 12540 1570 12544
rect 1506 12484 1510 12540
rect 1510 12484 1566 12540
rect 1566 12484 1570 12540
rect 1506 12480 1570 12484
rect 1586 12540 1650 12544
rect 1586 12484 1590 12540
rect 1590 12484 1646 12540
rect 1646 12484 1650 12540
rect 1586 12480 1650 12484
rect 1666 12540 1730 12544
rect 1666 12484 1670 12540
rect 1670 12484 1726 12540
rect 1726 12484 1730 12540
rect 1666 12480 1730 12484
rect 2374 12540 2438 12544
rect 2374 12484 2378 12540
rect 2378 12484 2434 12540
rect 2434 12484 2438 12540
rect 2374 12480 2438 12484
rect 2454 12540 2518 12544
rect 2454 12484 2458 12540
rect 2458 12484 2514 12540
rect 2514 12484 2518 12540
rect 2454 12480 2518 12484
rect 2534 12540 2598 12544
rect 2534 12484 2538 12540
rect 2538 12484 2594 12540
rect 2594 12484 2598 12540
rect 2534 12480 2598 12484
rect 2614 12540 2678 12544
rect 2614 12484 2618 12540
rect 2618 12484 2674 12540
rect 2674 12484 2678 12540
rect 2614 12480 2678 12484
rect 3322 12540 3386 12544
rect 3322 12484 3326 12540
rect 3326 12484 3382 12540
rect 3382 12484 3386 12540
rect 3322 12480 3386 12484
rect 3402 12540 3466 12544
rect 3402 12484 3406 12540
rect 3406 12484 3462 12540
rect 3462 12484 3466 12540
rect 3402 12480 3466 12484
rect 3482 12540 3546 12544
rect 3482 12484 3486 12540
rect 3486 12484 3542 12540
rect 3542 12484 3546 12540
rect 3482 12480 3546 12484
rect 3562 12540 3626 12544
rect 3562 12484 3566 12540
rect 3566 12484 3622 12540
rect 3622 12484 3626 12540
rect 3562 12480 3626 12484
rect 4270 12540 4334 12544
rect 4270 12484 4274 12540
rect 4274 12484 4330 12540
rect 4330 12484 4334 12540
rect 4270 12480 4334 12484
rect 4350 12540 4414 12544
rect 4350 12484 4354 12540
rect 4354 12484 4410 12540
rect 4410 12484 4414 12540
rect 4350 12480 4414 12484
rect 4430 12540 4494 12544
rect 4430 12484 4434 12540
rect 4434 12484 4490 12540
rect 4490 12484 4494 12540
rect 4430 12480 4494 12484
rect 4510 12540 4574 12544
rect 4510 12484 4514 12540
rect 4514 12484 4570 12540
rect 4570 12484 4574 12540
rect 4510 12480 4574 12484
rect 1900 11996 1964 12000
rect 1900 11940 1904 11996
rect 1904 11940 1960 11996
rect 1960 11940 1964 11996
rect 1900 11936 1964 11940
rect 1980 11996 2044 12000
rect 1980 11940 1984 11996
rect 1984 11940 2040 11996
rect 2040 11940 2044 11996
rect 1980 11936 2044 11940
rect 2060 11996 2124 12000
rect 2060 11940 2064 11996
rect 2064 11940 2120 11996
rect 2120 11940 2124 11996
rect 2060 11936 2124 11940
rect 2140 11996 2204 12000
rect 2140 11940 2144 11996
rect 2144 11940 2200 11996
rect 2200 11940 2204 11996
rect 2140 11936 2204 11940
rect 2848 11996 2912 12000
rect 2848 11940 2852 11996
rect 2852 11940 2908 11996
rect 2908 11940 2912 11996
rect 2848 11936 2912 11940
rect 2928 11996 2992 12000
rect 2928 11940 2932 11996
rect 2932 11940 2988 11996
rect 2988 11940 2992 11996
rect 2928 11936 2992 11940
rect 3008 11996 3072 12000
rect 3008 11940 3012 11996
rect 3012 11940 3068 11996
rect 3068 11940 3072 11996
rect 3008 11936 3072 11940
rect 3088 11996 3152 12000
rect 3088 11940 3092 11996
rect 3092 11940 3148 11996
rect 3148 11940 3152 11996
rect 3088 11936 3152 11940
rect 3796 11996 3860 12000
rect 3796 11940 3800 11996
rect 3800 11940 3856 11996
rect 3856 11940 3860 11996
rect 3796 11936 3860 11940
rect 3876 11996 3940 12000
rect 3876 11940 3880 11996
rect 3880 11940 3936 11996
rect 3936 11940 3940 11996
rect 3876 11936 3940 11940
rect 3956 11996 4020 12000
rect 3956 11940 3960 11996
rect 3960 11940 4016 11996
rect 4016 11940 4020 11996
rect 3956 11936 4020 11940
rect 4036 11996 4100 12000
rect 4036 11940 4040 11996
rect 4040 11940 4096 11996
rect 4096 11940 4100 11996
rect 4036 11936 4100 11940
rect 1426 11452 1490 11456
rect 1426 11396 1430 11452
rect 1430 11396 1486 11452
rect 1486 11396 1490 11452
rect 1426 11392 1490 11396
rect 1506 11452 1570 11456
rect 1506 11396 1510 11452
rect 1510 11396 1566 11452
rect 1566 11396 1570 11452
rect 1506 11392 1570 11396
rect 1586 11452 1650 11456
rect 1586 11396 1590 11452
rect 1590 11396 1646 11452
rect 1646 11396 1650 11452
rect 1586 11392 1650 11396
rect 1666 11452 1730 11456
rect 1666 11396 1670 11452
rect 1670 11396 1726 11452
rect 1726 11396 1730 11452
rect 1666 11392 1730 11396
rect 2374 11452 2438 11456
rect 2374 11396 2378 11452
rect 2378 11396 2434 11452
rect 2434 11396 2438 11452
rect 2374 11392 2438 11396
rect 2454 11452 2518 11456
rect 2454 11396 2458 11452
rect 2458 11396 2514 11452
rect 2514 11396 2518 11452
rect 2454 11392 2518 11396
rect 2534 11452 2598 11456
rect 2534 11396 2538 11452
rect 2538 11396 2594 11452
rect 2594 11396 2598 11452
rect 2534 11392 2598 11396
rect 2614 11452 2678 11456
rect 2614 11396 2618 11452
rect 2618 11396 2674 11452
rect 2674 11396 2678 11452
rect 2614 11392 2678 11396
rect 3322 11452 3386 11456
rect 3322 11396 3326 11452
rect 3326 11396 3382 11452
rect 3382 11396 3386 11452
rect 3322 11392 3386 11396
rect 3402 11452 3466 11456
rect 3402 11396 3406 11452
rect 3406 11396 3462 11452
rect 3462 11396 3466 11452
rect 3402 11392 3466 11396
rect 3482 11452 3546 11456
rect 3482 11396 3486 11452
rect 3486 11396 3542 11452
rect 3542 11396 3546 11452
rect 3482 11392 3546 11396
rect 3562 11452 3626 11456
rect 3562 11396 3566 11452
rect 3566 11396 3622 11452
rect 3622 11396 3626 11452
rect 3562 11392 3626 11396
rect 4270 11452 4334 11456
rect 4270 11396 4274 11452
rect 4274 11396 4330 11452
rect 4330 11396 4334 11452
rect 4270 11392 4334 11396
rect 4350 11452 4414 11456
rect 4350 11396 4354 11452
rect 4354 11396 4410 11452
rect 4410 11396 4414 11452
rect 4350 11392 4414 11396
rect 4430 11452 4494 11456
rect 4430 11396 4434 11452
rect 4434 11396 4490 11452
rect 4490 11396 4494 11452
rect 4430 11392 4494 11396
rect 4510 11452 4574 11456
rect 4510 11396 4514 11452
rect 4514 11396 4570 11452
rect 4570 11396 4574 11452
rect 4510 11392 4574 11396
rect 1900 10908 1964 10912
rect 1900 10852 1904 10908
rect 1904 10852 1960 10908
rect 1960 10852 1964 10908
rect 1900 10848 1964 10852
rect 1980 10908 2044 10912
rect 1980 10852 1984 10908
rect 1984 10852 2040 10908
rect 2040 10852 2044 10908
rect 1980 10848 2044 10852
rect 2060 10908 2124 10912
rect 2060 10852 2064 10908
rect 2064 10852 2120 10908
rect 2120 10852 2124 10908
rect 2060 10848 2124 10852
rect 2140 10908 2204 10912
rect 2140 10852 2144 10908
rect 2144 10852 2200 10908
rect 2200 10852 2204 10908
rect 2140 10848 2204 10852
rect 2848 10908 2912 10912
rect 2848 10852 2852 10908
rect 2852 10852 2908 10908
rect 2908 10852 2912 10908
rect 2848 10848 2912 10852
rect 2928 10908 2992 10912
rect 2928 10852 2932 10908
rect 2932 10852 2988 10908
rect 2988 10852 2992 10908
rect 2928 10848 2992 10852
rect 3008 10908 3072 10912
rect 3008 10852 3012 10908
rect 3012 10852 3068 10908
rect 3068 10852 3072 10908
rect 3008 10848 3072 10852
rect 3088 10908 3152 10912
rect 3088 10852 3092 10908
rect 3092 10852 3148 10908
rect 3148 10852 3152 10908
rect 3088 10848 3152 10852
rect 3796 10908 3860 10912
rect 3796 10852 3800 10908
rect 3800 10852 3856 10908
rect 3856 10852 3860 10908
rect 3796 10848 3860 10852
rect 3876 10908 3940 10912
rect 3876 10852 3880 10908
rect 3880 10852 3936 10908
rect 3936 10852 3940 10908
rect 3876 10848 3940 10852
rect 3956 10908 4020 10912
rect 3956 10852 3960 10908
rect 3960 10852 4016 10908
rect 4016 10852 4020 10908
rect 3956 10848 4020 10852
rect 4036 10908 4100 10912
rect 4036 10852 4040 10908
rect 4040 10852 4096 10908
rect 4096 10852 4100 10908
rect 4036 10848 4100 10852
rect 1426 10364 1490 10368
rect 1426 10308 1430 10364
rect 1430 10308 1486 10364
rect 1486 10308 1490 10364
rect 1426 10304 1490 10308
rect 1506 10364 1570 10368
rect 1506 10308 1510 10364
rect 1510 10308 1566 10364
rect 1566 10308 1570 10364
rect 1506 10304 1570 10308
rect 1586 10364 1650 10368
rect 1586 10308 1590 10364
rect 1590 10308 1646 10364
rect 1646 10308 1650 10364
rect 1586 10304 1650 10308
rect 1666 10364 1730 10368
rect 1666 10308 1670 10364
rect 1670 10308 1726 10364
rect 1726 10308 1730 10364
rect 1666 10304 1730 10308
rect 2374 10364 2438 10368
rect 2374 10308 2378 10364
rect 2378 10308 2434 10364
rect 2434 10308 2438 10364
rect 2374 10304 2438 10308
rect 2454 10364 2518 10368
rect 2454 10308 2458 10364
rect 2458 10308 2514 10364
rect 2514 10308 2518 10364
rect 2454 10304 2518 10308
rect 2534 10364 2598 10368
rect 2534 10308 2538 10364
rect 2538 10308 2594 10364
rect 2594 10308 2598 10364
rect 2534 10304 2598 10308
rect 2614 10364 2678 10368
rect 2614 10308 2618 10364
rect 2618 10308 2674 10364
rect 2674 10308 2678 10364
rect 2614 10304 2678 10308
rect 3322 10364 3386 10368
rect 3322 10308 3326 10364
rect 3326 10308 3382 10364
rect 3382 10308 3386 10364
rect 3322 10304 3386 10308
rect 3402 10364 3466 10368
rect 3402 10308 3406 10364
rect 3406 10308 3462 10364
rect 3462 10308 3466 10364
rect 3402 10304 3466 10308
rect 3482 10364 3546 10368
rect 3482 10308 3486 10364
rect 3486 10308 3542 10364
rect 3542 10308 3546 10364
rect 3482 10304 3546 10308
rect 3562 10364 3626 10368
rect 3562 10308 3566 10364
rect 3566 10308 3622 10364
rect 3622 10308 3626 10364
rect 3562 10304 3626 10308
rect 4270 10364 4334 10368
rect 4270 10308 4274 10364
rect 4274 10308 4330 10364
rect 4330 10308 4334 10364
rect 4270 10304 4334 10308
rect 4350 10364 4414 10368
rect 4350 10308 4354 10364
rect 4354 10308 4410 10364
rect 4410 10308 4414 10364
rect 4350 10304 4414 10308
rect 4430 10364 4494 10368
rect 4430 10308 4434 10364
rect 4434 10308 4490 10364
rect 4490 10308 4494 10364
rect 4430 10304 4494 10308
rect 4510 10364 4574 10368
rect 4510 10308 4514 10364
rect 4514 10308 4570 10364
rect 4570 10308 4574 10364
rect 4510 10304 4574 10308
rect 1900 9820 1964 9824
rect 1900 9764 1904 9820
rect 1904 9764 1960 9820
rect 1960 9764 1964 9820
rect 1900 9760 1964 9764
rect 1980 9820 2044 9824
rect 1980 9764 1984 9820
rect 1984 9764 2040 9820
rect 2040 9764 2044 9820
rect 1980 9760 2044 9764
rect 2060 9820 2124 9824
rect 2060 9764 2064 9820
rect 2064 9764 2120 9820
rect 2120 9764 2124 9820
rect 2060 9760 2124 9764
rect 2140 9820 2204 9824
rect 2140 9764 2144 9820
rect 2144 9764 2200 9820
rect 2200 9764 2204 9820
rect 2140 9760 2204 9764
rect 2848 9820 2912 9824
rect 2848 9764 2852 9820
rect 2852 9764 2908 9820
rect 2908 9764 2912 9820
rect 2848 9760 2912 9764
rect 2928 9820 2992 9824
rect 2928 9764 2932 9820
rect 2932 9764 2988 9820
rect 2988 9764 2992 9820
rect 2928 9760 2992 9764
rect 3008 9820 3072 9824
rect 3008 9764 3012 9820
rect 3012 9764 3068 9820
rect 3068 9764 3072 9820
rect 3008 9760 3072 9764
rect 3088 9820 3152 9824
rect 3088 9764 3092 9820
rect 3092 9764 3148 9820
rect 3148 9764 3152 9820
rect 3088 9760 3152 9764
rect 3796 9820 3860 9824
rect 3796 9764 3800 9820
rect 3800 9764 3856 9820
rect 3856 9764 3860 9820
rect 3796 9760 3860 9764
rect 3876 9820 3940 9824
rect 3876 9764 3880 9820
rect 3880 9764 3936 9820
rect 3936 9764 3940 9820
rect 3876 9760 3940 9764
rect 3956 9820 4020 9824
rect 3956 9764 3960 9820
rect 3960 9764 4016 9820
rect 4016 9764 4020 9820
rect 3956 9760 4020 9764
rect 4036 9820 4100 9824
rect 4036 9764 4040 9820
rect 4040 9764 4096 9820
rect 4096 9764 4100 9820
rect 4036 9760 4100 9764
rect 1426 9276 1490 9280
rect 1426 9220 1430 9276
rect 1430 9220 1486 9276
rect 1486 9220 1490 9276
rect 1426 9216 1490 9220
rect 1506 9276 1570 9280
rect 1506 9220 1510 9276
rect 1510 9220 1566 9276
rect 1566 9220 1570 9276
rect 1506 9216 1570 9220
rect 1586 9276 1650 9280
rect 1586 9220 1590 9276
rect 1590 9220 1646 9276
rect 1646 9220 1650 9276
rect 1586 9216 1650 9220
rect 1666 9276 1730 9280
rect 1666 9220 1670 9276
rect 1670 9220 1726 9276
rect 1726 9220 1730 9276
rect 1666 9216 1730 9220
rect 2374 9276 2438 9280
rect 2374 9220 2378 9276
rect 2378 9220 2434 9276
rect 2434 9220 2438 9276
rect 2374 9216 2438 9220
rect 2454 9276 2518 9280
rect 2454 9220 2458 9276
rect 2458 9220 2514 9276
rect 2514 9220 2518 9276
rect 2454 9216 2518 9220
rect 2534 9276 2598 9280
rect 2534 9220 2538 9276
rect 2538 9220 2594 9276
rect 2594 9220 2598 9276
rect 2534 9216 2598 9220
rect 2614 9276 2678 9280
rect 2614 9220 2618 9276
rect 2618 9220 2674 9276
rect 2674 9220 2678 9276
rect 2614 9216 2678 9220
rect 3322 9276 3386 9280
rect 3322 9220 3326 9276
rect 3326 9220 3382 9276
rect 3382 9220 3386 9276
rect 3322 9216 3386 9220
rect 3402 9276 3466 9280
rect 3402 9220 3406 9276
rect 3406 9220 3462 9276
rect 3462 9220 3466 9276
rect 3402 9216 3466 9220
rect 3482 9276 3546 9280
rect 3482 9220 3486 9276
rect 3486 9220 3542 9276
rect 3542 9220 3546 9276
rect 3482 9216 3546 9220
rect 3562 9276 3626 9280
rect 3562 9220 3566 9276
rect 3566 9220 3622 9276
rect 3622 9220 3626 9276
rect 3562 9216 3626 9220
rect 4270 9276 4334 9280
rect 4270 9220 4274 9276
rect 4274 9220 4330 9276
rect 4330 9220 4334 9276
rect 4270 9216 4334 9220
rect 4350 9276 4414 9280
rect 4350 9220 4354 9276
rect 4354 9220 4410 9276
rect 4410 9220 4414 9276
rect 4350 9216 4414 9220
rect 4430 9276 4494 9280
rect 4430 9220 4434 9276
rect 4434 9220 4490 9276
rect 4490 9220 4494 9276
rect 4430 9216 4494 9220
rect 4510 9276 4574 9280
rect 4510 9220 4514 9276
rect 4514 9220 4570 9276
rect 4570 9220 4574 9276
rect 4510 9216 4574 9220
rect 1900 8732 1964 8736
rect 1900 8676 1904 8732
rect 1904 8676 1960 8732
rect 1960 8676 1964 8732
rect 1900 8672 1964 8676
rect 1980 8732 2044 8736
rect 1980 8676 1984 8732
rect 1984 8676 2040 8732
rect 2040 8676 2044 8732
rect 1980 8672 2044 8676
rect 2060 8732 2124 8736
rect 2060 8676 2064 8732
rect 2064 8676 2120 8732
rect 2120 8676 2124 8732
rect 2060 8672 2124 8676
rect 2140 8732 2204 8736
rect 2140 8676 2144 8732
rect 2144 8676 2200 8732
rect 2200 8676 2204 8732
rect 2140 8672 2204 8676
rect 2848 8732 2912 8736
rect 2848 8676 2852 8732
rect 2852 8676 2908 8732
rect 2908 8676 2912 8732
rect 2848 8672 2912 8676
rect 2928 8732 2992 8736
rect 2928 8676 2932 8732
rect 2932 8676 2988 8732
rect 2988 8676 2992 8732
rect 2928 8672 2992 8676
rect 3008 8732 3072 8736
rect 3008 8676 3012 8732
rect 3012 8676 3068 8732
rect 3068 8676 3072 8732
rect 3008 8672 3072 8676
rect 3088 8732 3152 8736
rect 3088 8676 3092 8732
rect 3092 8676 3148 8732
rect 3148 8676 3152 8732
rect 3088 8672 3152 8676
rect 3796 8732 3860 8736
rect 3796 8676 3800 8732
rect 3800 8676 3856 8732
rect 3856 8676 3860 8732
rect 3796 8672 3860 8676
rect 3876 8732 3940 8736
rect 3876 8676 3880 8732
rect 3880 8676 3936 8732
rect 3936 8676 3940 8732
rect 3876 8672 3940 8676
rect 3956 8732 4020 8736
rect 3956 8676 3960 8732
rect 3960 8676 4016 8732
rect 4016 8676 4020 8732
rect 3956 8672 4020 8676
rect 4036 8732 4100 8736
rect 4036 8676 4040 8732
rect 4040 8676 4096 8732
rect 4096 8676 4100 8732
rect 4036 8672 4100 8676
rect 1426 8188 1490 8192
rect 1426 8132 1430 8188
rect 1430 8132 1486 8188
rect 1486 8132 1490 8188
rect 1426 8128 1490 8132
rect 1506 8188 1570 8192
rect 1506 8132 1510 8188
rect 1510 8132 1566 8188
rect 1566 8132 1570 8188
rect 1506 8128 1570 8132
rect 1586 8188 1650 8192
rect 1586 8132 1590 8188
rect 1590 8132 1646 8188
rect 1646 8132 1650 8188
rect 1586 8128 1650 8132
rect 1666 8188 1730 8192
rect 1666 8132 1670 8188
rect 1670 8132 1726 8188
rect 1726 8132 1730 8188
rect 1666 8128 1730 8132
rect 2374 8188 2438 8192
rect 2374 8132 2378 8188
rect 2378 8132 2434 8188
rect 2434 8132 2438 8188
rect 2374 8128 2438 8132
rect 2454 8188 2518 8192
rect 2454 8132 2458 8188
rect 2458 8132 2514 8188
rect 2514 8132 2518 8188
rect 2454 8128 2518 8132
rect 2534 8188 2598 8192
rect 2534 8132 2538 8188
rect 2538 8132 2594 8188
rect 2594 8132 2598 8188
rect 2534 8128 2598 8132
rect 2614 8188 2678 8192
rect 2614 8132 2618 8188
rect 2618 8132 2674 8188
rect 2674 8132 2678 8188
rect 2614 8128 2678 8132
rect 3322 8188 3386 8192
rect 3322 8132 3326 8188
rect 3326 8132 3382 8188
rect 3382 8132 3386 8188
rect 3322 8128 3386 8132
rect 3402 8188 3466 8192
rect 3402 8132 3406 8188
rect 3406 8132 3462 8188
rect 3462 8132 3466 8188
rect 3402 8128 3466 8132
rect 3482 8188 3546 8192
rect 3482 8132 3486 8188
rect 3486 8132 3542 8188
rect 3542 8132 3546 8188
rect 3482 8128 3546 8132
rect 3562 8188 3626 8192
rect 3562 8132 3566 8188
rect 3566 8132 3622 8188
rect 3622 8132 3626 8188
rect 3562 8128 3626 8132
rect 4270 8188 4334 8192
rect 4270 8132 4274 8188
rect 4274 8132 4330 8188
rect 4330 8132 4334 8188
rect 4270 8128 4334 8132
rect 4350 8188 4414 8192
rect 4350 8132 4354 8188
rect 4354 8132 4410 8188
rect 4410 8132 4414 8188
rect 4350 8128 4414 8132
rect 4430 8188 4494 8192
rect 4430 8132 4434 8188
rect 4434 8132 4490 8188
rect 4490 8132 4494 8188
rect 4430 8128 4494 8132
rect 4510 8188 4574 8192
rect 4510 8132 4514 8188
rect 4514 8132 4570 8188
rect 4570 8132 4574 8188
rect 4510 8128 4574 8132
rect 1900 7644 1964 7648
rect 1900 7588 1904 7644
rect 1904 7588 1960 7644
rect 1960 7588 1964 7644
rect 1900 7584 1964 7588
rect 1980 7644 2044 7648
rect 1980 7588 1984 7644
rect 1984 7588 2040 7644
rect 2040 7588 2044 7644
rect 1980 7584 2044 7588
rect 2060 7644 2124 7648
rect 2060 7588 2064 7644
rect 2064 7588 2120 7644
rect 2120 7588 2124 7644
rect 2060 7584 2124 7588
rect 2140 7644 2204 7648
rect 2140 7588 2144 7644
rect 2144 7588 2200 7644
rect 2200 7588 2204 7644
rect 2140 7584 2204 7588
rect 2848 7644 2912 7648
rect 2848 7588 2852 7644
rect 2852 7588 2908 7644
rect 2908 7588 2912 7644
rect 2848 7584 2912 7588
rect 2928 7644 2992 7648
rect 2928 7588 2932 7644
rect 2932 7588 2988 7644
rect 2988 7588 2992 7644
rect 2928 7584 2992 7588
rect 3008 7644 3072 7648
rect 3008 7588 3012 7644
rect 3012 7588 3068 7644
rect 3068 7588 3072 7644
rect 3008 7584 3072 7588
rect 3088 7644 3152 7648
rect 3088 7588 3092 7644
rect 3092 7588 3148 7644
rect 3148 7588 3152 7644
rect 3088 7584 3152 7588
rect 3796 7644 3860 7648
rect 3796 7588 3800 7644
rect 3800 7588 3856 7644
rect 3856 7588 3860 7644
rect 3796 7584 3860 7588
rect 3876 7644 3940 7648
rect 3876 7588 3880 7644
rect 3880 7588 3936 7644
rect 3936 7588 3940 7644
rect 3876 7584 3940 7588
rect 3956 7644 4020 7648
rect 3956 7588 3960 7644
rect 3960 7588 4016 7644
rect 4016 7588 4020 7644
rect 3956 7584 4020 7588
rect 4036 7644 4100 7648
rect 4036 7588 4040 7644
rect 4040 7588 4096 7644
rect 4096 7588 4100 7644
rect 4036 7584 4100 7588
rect 1426 7100 1490 7104
rect 1426 7044 1430 7100
rect 1430 7044 1486 7100
rect 1486 7044 1490 7100
rect 1426 7040 1490 7044
rect 1506 7100 1570 7104
rect 1506 7044 1510 7100
rect 1510 7044 1566 7100
rect 1566 7044 1570 7100
rect 1506 7040 1570 7044
rect 1586 7100 1650 7104
rect 1586 7044 1590 7100
rect 1590 7044 1646 7100
rect 1646 7044 1650 7100
rect 1586 7040 1650 7044
rect 1666 7100 1730 7104
rect 1666 7044 1670 7100
rect 1670 7044 1726 7100
rect 1726 7044 1730 7100
rect 1666 7040 1730 7044
rect 2374 7100 2438 7104
rect 2374 7044 2378 7100
rect 2378 7044 2434 7100
rect 2434 7044 2438 7100
rect 2374 7040 2438 7044
rect 2454 7100 2518 7104
rect 2454 7044 2458 7100
rect 2458 7044 2514 7100
rect 2514 7044 2518 7100
rect 2454 7040 2518 7044
rect 2534 7100 2598 7104
rect 2534 7044 2538 7100
rect 2538 7044 2594 7100
rect 2594 7044 2598 7100
rect 2534 7040 2598 7044
rect 2614 7100 2678 7104
rect 2614 7044 2618 7100
rect 2618 7044 2674 7100
rect 2674 7044 2678 7100
rect 2614 7040 2678 7044
rect 3322 7100 3386 7104
rect 3322 7044 3326 7100
rect 3326 7044 3382 7100
rect 3382 7044 3386 7100
rect 3322 7040 3386 7044
rect 3402 7100 3466 7104
rect 3402 7044 3406 7100
rect 3406 7044 3462 7100
rect 3462 7044 3466 7100
rect 3402 7040 3466 7044
rect 3482 7100 3546 7104
rect 3482 7044 3486 7100
rect 3486 7044 3542 7100
rect 3542 7044 3546 7100
rect 3482 7040 3546 7044
rect 3562 7100 3626 7104
rect 3562 7044 3566 7100
rect 3566 7044 3622 7100
rect 3622 7044 3626 7100
rect 3562 7040 3626 7044
rect 4270 7100 4334 7104
rect 4270 7044 4274 7100
rect 4274 7044 4330 7100
rect 4330 7044 4334 7100
rect 4270 7040 4334 7044
rect 4350 7100 4414 7104
rect 4350 7044 4354 7100
rect 4354 7044 4410 7100
rect 4410 7044 4414 7100
rect 4350 7040 4414 7044
rect 4430 7100 4494 7104
rect 4430 7044 4434 7100
rect 4434 7044 4490 7100
rect 4490 7044 4494 7100
rect 4430 7040 4494 7044
rect 4510 7100 4574 7104
rect 4510 7044 4514 7100
rect 4514 7044 4570 7100
rect 4570 7044 4574 7100
rect 4510 7040 4574 7044
rect 1900 6556 1964 6560
rect 1900 6500 1904 6556
rect 1904 6500 1960 6556
rect 1960 6500 1964 6556
rect 1900 6496 1964 6500
rect 1980 6556 2044 6560
rect 1980 6500 1984 6556
rect 1984 6500 2040 6556
rect 2040 6500 2044 6556
rect 1980 6496 2044 6500
rect 2060 6556 2124 6560
rect 2060 6500 2064 6556
rect 2064 6500 2120 6556
rect 2120 6500 2124 6556
rect 2060 6496 2124 6500
rect 2140 6556 2204 6560
rect 2140 6500 2144 6556
rect 2144 6500 2200 6556
rect 2200 6500 2204 6556
rect 2140 6496 2204 6500
rect 2848 6556 2912 6560
rect 2848 6500 2852 6556
rect 2852 6500 2908 6556
rect 2908 6500 2912 6556
rect 2848 6496 2912 6500
rect 2928 6556 2992 6560
rect 2928 6500 2932 6556
rect 2932 6500 2988 6556
rect 2988 6500 2992 6556
rect 2928 6496 2992 6500
rect 3008 6556 3072 6560
rect 3008 6500 3012 6556
rect 3012 6500 3068 6556
rect 3068 6500 3072 6556
rect 3008 6496 3072 6500
rect 3088 6556 3152 6560
rect 3088 6500 3092 6556
rect 3092 6500 3148 6556
rect 3148 6500 3152 6556
rect 3088 6496 3152 6500
rect 3796 6556 3860 6560
rect 3796 6500 3800 6556
rect 3800 6500 3856 6556
rect 3856 6500 3860 6556
rect 3796 6496 3860 6500
rect 3876 6556 3940 6560
rect 3876 6500 3880 6556
rect 3880 6500 3936 6556
rect 3936 6500 3940 6556
rect 3876 6496 3940 6500
rect 3956 6556 4020 6560
rect 3956 6500 3960 6556
rect 3960 6500 4016 6556
rect 4016 6500 4020 6556
rect 3956 6496 4020 6500
rect 4036 6556 4100 6560
rect 4036 6500 4040 6556
rect 4040 6500 4096 6556
rect 4096 6500 4100 6556
rect 4036 6496 4100 6500
rect 1426 6012 1490 6016
rect 1426 5956 1430 6012
rect 1430 5956 1486 6012
rect 1486 5956 1490 6012
rect 1426 5952 1490 5956
rect 1506 6012 1570 6016
rect 1506 5956 1510 6012
rect 1510 5956 1566 6012
rect 1566 5956 1570 6012
rect 1506 5952 1570 5956
rect 1586 6012 1650 6016
rect 1586 5956 1590 6012
rect 1590 5956 1646 6012
rect 1646 5956 1650 6012
rect 1586 5952 1650 5956
rect 1666 6012 1730 6016
rect 1666 5956 1670 6012
rect 1670 5956 1726 6012
rect 1726 5956 1730 6012
rect 1666 5952 1730 5956
rect 2374 6012 2438 6016
rect 2374 5956 2378 6012
rect 2378 5956 2434 6012
rect 2434 5956 2438 6012
rect 2374 5952 2438 5956
rect 2454 6012 2518 6016
rect 2454 5956 2458 6012
rect 2458 5956 2514 6012
rect 2514 5956 2518 6012
rect 2454 5952 2518 5956
rect 2534 6012 2598 6016
rect 2534 5956 2538 6012
rect 2538 5956 2594 6012
rect 2594 5956 2598 6012
rect 2534 5952 2598 5956
rect 2614 6012 2678 6016
rect 2614 5956 2618 6012
rect 2618 5956 2674 6012
rect 2674 5956 2678 6012
rect 2614 5952 2678 5956
rect 3322 6012 3386 6016
rect 3322 5956 3326 6012
rect 3326 5956 3382 6012
rect 3382 5956 3386 6012
rect 3322 5952 3386 5956
rect 3402 6012 3466 6016
rect 3402 5956 3406 6012
rect 3406 5956 3462 6012
rect 3462 5956 3466 6012
rect 3402 5952 3466 5956
rect 3482 6012 3546 6016
rect 3482 5956 3486 6012
rect 3486 5956 3542 6012
rect 3542 5956 3546 6012
rect 3482 5952 3546 5956
rect 3562 6012 3626 6016
rect 3562 5956 3566 6012
rect 3566 5956 3622 6012
rect 3622 5956 3626 6012
rect 3562 5952 3626 5956
rect 4270 6012 4334 6016
rect 4270 5956 4274 6012
rect 4274 5956 4330 6012
rect 4330 5956 4334 6012
rect 4270 5952 4334 5956
rect 4350 6012 4414 6016
rect 4350 5956 4354 6012
rect 4354 5956 4410 6012
rect 4410 5956 4414 6012
rect 4350 5952 4414 5956
rect 4430 6012 4494 6016
rect 4430 5956 4434 6012
rect 4434 5956 4490 6012
rect 4490 5956 4494 6012
rect 4430 5952 4494 5956
rect 4510 6012 4574 6016
rect 4510 5956 4514 6012
rect 4514 5956 4570 6012
rect 4570 5956 4574 6012
rect 4510 5952 4574 5956
rect 1900 5468 1964 5472
rect 1900 5412 1904 5468
rect 1904 5412 1960 5468
rect 1960 5412 1964 5468
rect 1900 5408 1964 5412
rect 1980 5468 2044 5472
rect 1980 5412 1984 5468
rect 1984 5412 2040 5468
rect 2040 5412 2044 5468
rect 1980 5408 2044 5412
rect 2060 5468 2124 5472
rect 2060 5412 2064 5468
rect 2064 5412 2120 5468
rect 2120 5412 2124 5468
rect 2060 5408 2124 5412
rect 2140 5468 2204 5472
rect 2140 5412 2144 5468
rect 2144 5412 2200 5468
rect 2200 5412 2204 5468
rect 2140 5408 2204 5412
rect 2848 5468 2912 5472
rect 2848 5412 2852 5468
rect 2852 5412 2908 5468
rect 2908 5412 2912 5468
rect 2848 5408 2912 5412
rect 2928 5468 2992 5472
rect 2928 5412 2932 5468
rect 2932 5412 2988 5468
rect 2988 5412 2992 5468
rect 2928 5408 2992 5412
rect 3008 5468 3072 5472
rect 3008 5412 3012 5468
rect 3012 5412 3068 5468
rect 3068 5412 3072 5468
rect 3008 5408 3072 5412
rect 3088 5468 3152 5472
rect 3088 5412 3092 5468
rect 3092 5412 3148 5468
rect 3148 5412 3152 5468
rect 3088 5408 3152 5412
rect 3796 5468 3860 5472
rect 3796 5412 3800 5468
rect 3800 5412 3856 5468
rect 3856 5412 3860 5468
rect 3796 5408 3860 5412
rect 3876 5468 3940 5472
rect 3876 5412 3880 5468
rect 3880 5412 3936 5468
rect 3936 5412 3940 5468
rect 3876 5408 3940 5412
rect 3956 5468 4020 5472
rect 3956 5412 3960 5468
rect 3960 5412 4016 5468
rect 4016 5412 4020 5468
rect 3956 5408 4020 5412
rect 4036 5468 4100 5472
rect 4036 5412 4040 5468
rect 4040 5412 4096 5468
rect 4096 5412 4100 5468
rect 4036 5408 4100 5412
rect 1426 4924 1490 4928
rect 1426 4868 1430 4924
rect 1430 4868 1486 4924
rect 1486 4868 1490 4924
rect 1426 4864 1490 4868
rect 1506 4924 1570 4928
rect 1506 4868 1510 4924
rect 1510 4868 1566 4924
rect 1566 4868 1570 4924
rect 1506 4864 1570 4868
rect 1586 4924 1650 4928
rect 1586 4868 1590 4924
rect 1590 4868 1646 4924
rect 1646 4868 1650 4924
rect 1586 4864 1650 4868
rect 1666 4924 1730 4928
rect 1666 4868 1670 4924
rect 1670 4868 1726 4924
rect 1726 4868 1730 4924
rect 1666 4864 1730 4868
rect 2374 4924 2438 4928
rect 2374 4868 2378 4924
rect 2378 4868 2434 4924
rect 2434 4868 2438 4924
rect 2374 4864 2438 4868
rect 2454 4924 2518 4928
rect 2454 4868 2458 4924
rect 2458 4868 2514 4924
rect 2514 4868 2518 4924
rect 2454 4864 2518 4868
rect 2534 4924 2598 4928
rect 2534 4868 2538 4924
rect 2538 4868 2594 4924
rect 2594 4868 2598 4924
rect 2534 4864 2598 4868
rect 2614 4924 2678 4928
rect 2614 4868 2618 4924
rect 2618 4868 2674 4924
rect 2674 4868 2678 4924
rect 2614 4864 2678 4868
rect 3322 4924 3386 4928
rect 3322 4868 3326 4924
rect 3326 4868 3382 4924
rect 3382 4868 3386 4924
rect 3322 4864 3386 4868
rect 3402 4924 3466 4928
rect 3402 4868 3406 4924
rect 3406 4868 3462 4924
rect 3462 4868 3466 4924
rect 3402 4864 3466 4868
rect 3482 4924 3546 4928
rect 3482 4868 3486 4924
rect 3486 4868 3542 4924
rect 3542 4868 3546 4924
rect 3482 4864 3546 4868
rect 3562 4924 3626 4928
rect 3562 4868 3566 4924
rect 3566 4868 3622 4924
rect 3622 4868 3626 4924
rect 3562 4864 3626 4868
rect 4270 4924 4334 4928
rect 4270 4868 4274 4924
rect 4274 4868 4330 4924
rect 4330 4868 4334 4924
rect 4270 4864 4334 4868
rect 4350 4924 4414 4928
rect 4350 4868 4354 4924
rect 4354 4868 4410 4924
rect 4410 4868 4414 4924
rect 4350 4864 4414 4868
rect 4430 4924 4494 4928
rect 4430 4868 4434 4924
rect 4434 4868 4490 4924
rect 4490 4868 4494 4924
rect 4430 4864 4494 4868
rect 4510 4924 4574 4928
rect 4510 4868 4514 4924
rect 4514 4868 4570 4924
rect 4570 4868 4574 4924
rect 4510 4864 4574 4868
rect 1900 4380 1964 4384
rect 1900 4324 1904 4380
rect 1904 4324 1960 4380
rect 1960 4324 1964 4380
rect 1900 4320 1964 4324
rect 1980 4380 2044 4384
rect 1980 4324 1984 4380
rect 1984 4324 2040 4380
rect 2040 4324 2044 4380
rect 1980 4320 2044 4324
rect 2060 4380 2124 4384
rect 2060 4324 2064 4380
rect 2064 4324 2120 4380
rect 2120 4324 2124 4380
rect 2060 4320 2124 4324
rect 2140 4380 2204 4384
rect 2140 4324 2144 4380
rect 2144 4324 2200 4380
rect 2200 4324 2204 4380
rect 2140 4320 2204 4324
rect 2848 4380 2912 4384
rect 2848 4324 2852 4380
rect 2852 4324 2908 4380
rect 2908 4324 2912 4380
rect 2848 4320 2912 4324
rect 2928 4380 2992 4384
rect 2928 4324 2932 4380
rect 2932 4324 2988 4380
rect 2988 4324 2992 4380
rect 2928 4320 2992 4324
rect 3008 4380 3072 4384
rect 3008 4324 3012 4380
rect 3012 4324 3068 4380
rect 3068 4324 3072 4380
rect 3008 4320 3072 4324
rect 3088 4380 3152 4384
rect 3088 4324 3092 4380
rect 3092 4324 3148 4380
rect 3148 4324 3152 4380
rect 3088 4320 3152 4324
rect 3796 4380 3860 4384
rect 3796 4324 3800 4380
rect 3800 4324 3856 4380
rect 3856 4324 3860 4380
rect 3796 4320 3860 4324
rect 3876 4380 3940 4384
rect 3876 4324 3880 4380
rect 3880 4324 3936 4380
rect 3936 4324 3940 4380
rect 3876 4320 3940 4324
rect 3956 4380 4020 4384
rect 3956 4324 3960 4380
rect 3960 4324 4016 4380
rect 4016 4324 4020 4380
rect 3956 4320 4020 4324
rect 4036 4380 4100 4384
rect 4036 4324 4040 4380
rect 4040 4324 4096 4380
rect 4096 4324 4100 4380
rect 4036 4320 4100 4324
rect 1426 3836 1490 3840
rect 1426 3780 1430 3836
rect 1430 3780 1486 3836
rect 1486 3780 1490 3836
rect 1426 3776 1490 3780
rect 1506 3836 1570 3840
rect 1506 3780 1510 3836
rect 1510 3780 1566 3836
rect 1566 3780 1570 3836
rect 1506 3776 1570 3780
rect 1586 3836 1650 3840
rect 1586 3780 1590 3836
rect 1590 3780 1646 3836
rect 1646 3780 1650 3836
rect 1586 3776 1650 3780
rect 1666 3836 1730 3840
rect 1666 3780 1670 3836
rect 1670 3780 1726 3836
rect 1726 3780 1730 3836
rect 1666 3776 1730 3780
rect 2374 3836 2438 3840
rect 2374 3780 2378 3836
rect 2378 3780 2434 3836
rect 2434 3780 2438 3836
rect 2374 3776 2438 3780
rect 2454 3836 2518 3840
rect 2454 3780 2458 3836
rect 2458 3780 2514 3836
rect 2514 3780 2518 3836
rect 2454 3776 2518 3780
rect 2534 3836 2598 3840
rect 2534 3780 2538 3836
rect 2538 3780 2594 3836
rect 2594 3780 2598 3836
rect 2534 3776 2598 3780
rect 2614 3836 2678 3840
rect 2614 3780 2618 3836
rect 2618 3780 2674 3836
rect 2674 3780 2678 3836
rect 2614 3776 2678 3780
rect 3322 3836 3386 3840
rect 3322 3780 3326 3836
rect 3326 3780 3382 3836
rect 3382 3780 3386 3836
rect 3322 3776 3386 3780
rect 3402 3836 3466 3840
rect 3402 3780 3406 3836
rect 3406 3780 3462 3836
rect 3462 3780 3466 3836
rect 3402 3776 3466 3780
rect 3482 3836 3546 3840
rect 3482 3780 3486 3836
rect 3486 3780 3542 3836
rect 3542 3780 3546 3836
rect 3482 3776 3546 3780
rect 3562 3836 3626 3840
rect 3562 3780 3566 3836
rect 3566 3780 3622 3836
rect 3622 3780 3626 3836
rect 3562 3776 3626 3780
rect 4270 3836 4334 3840
rect 4270 3780 4274 3836
rect 4274 3780 4330 3836
rect 4330 3780 4334 3836
rect 4270 3776 4334 3780
rect 4350 3836 4414 3840
rect 4350 3780 4354 3836
rect 4354 3780 4410 3836
rect 4410 3780 4414 3836
rect 4350 3776 4414 3780
rect 4430 3836 4494 3840
rect 4430 3780 4434 3836
rect 4434 3780 4490 3836
rect 4490 3780 4494 3836
rect 4430 3776 4494 3780
rect 4510 3836 4574 3840
rect 4510 3780 4514 3836
rect 4514 3780 4570 3836
rect 4570 3780 4574 3836
rect 4510 3776 4574 3780
rect 1900 3292 1964 3296
rect 1900 3236 1904 3292
rect 1904 3236 1960 3292
rect 1960 3236 1964 3292
rect 1900 3232 1964 3236
rect 1980 3292 2044 3296
rect 1980 3236 1984 3292
rect 1984 3236 2040 3292
rect 2040 3236 2044 3292
rect 1980 3232 2044 3236
rect 2060 3292 2124 3296
rect 2060 3236 2064 3292
rect 2064 3236 2120 3292
rect 2120 3236 2124 3292
rect 2060 3232 2124 3236
rect 2140 3292 2204 3296
rect 2140 3236 2144 3292
rect 2144 3236 2200 3292
rect 2200 3236 2204 3292
rect 2140 3232 2204 3236
rect 2848 3292 2912 3296
rect 2848 3236 2852 3292
rect 2852 3236 2908 3292
rect 2908 3236 2912 3292
rect 2848 3232 2912 3236
rect 2928 3292 2992 3296
rect 2928 3236 2932 3292
rect 2932 3236 2988 3292
rect 2988 3236 2992 3292
rect 2928 3232 2992 3236
rect 3008 3292 3072 3296
rect 3008 3236 3012 3292
rect 3012 3236 3068 3292
rect 3068 3236 3072 3292
rect 3008 3232 3072 3236
rect 3088 3292 3152 3296
rect 3088 3236 3092 3292
rect 3092 3236 3148 3292
rect 3148 3236 3152 3292
rect 3088 3232 3152 3236
rect 3796 3292 3860 3296
rect 3796 3236 3800 3292
rect 3800 3236 3856 3292
rect 3856 3236 3860 3292
rect 3796 3232 3860 3236
rect 3876 3292 3940 3296
rect 3876 3236 3880 3292
rect 3880 3236 3936 3292
rect 3936 3236 3940 3292
rect 3876 3232 3940 3236
rect 3956 3292 4020 3296
rect 3956 3236 3960 3292
rect 3960 3236 4016 3292
rect 4016 3236 4020 3292
rect 3956 3232 4020 3236
rect 4036 3292 4100 3296
rect 4036 3236 4040 3292
rect 4040 3236 4096 3292
rect 4096 3236 4100 3292
rect 4036 3232 4100 3236
rect 1426 2748 1490 2752
rect 1426 2692 1430 2748
rect 1430 2692 1486 2748
rect 1486 2692 1490 2748
rect 1426 2688 1490 2692
rect 1506 2748 1570 2752
rect 1506 2692 1510 2748
rect 1510 2692 1566 2748
rect 1566 2692 1570 2748
rect 1506 2688 1570 2692
rect 1586 2748 1650 2752
rect 1586 2692 1590 2748
rect 1590 2692 1646 2748
rect 1646 2692 1650 2748
rect 1586 2688 1650 2692
rect 1666 2748 1730 2752
rect 1666 2692 1670 2748
rect 1670 2692 1726 2748
rect 1726 2692 1730 2748
rect 1666 2688 1730 2692
rect 2374 2748 2438 2752
rect 2374 2692 2378 2748
rect 2378 2692 2434 2748
rect 2434 2692 2438 2748
rect 2374 2688 2438 2692
rect 2454 2748 2518 2752
rect 2454 2692 2458 2748
rect 2458 2692 2514 2748
rect 2514 2692 2518 2748
rect 2454 2688 2518 2692
rect 2534 2748 2598 2752
rect 2534 2692 2538 2748
rect 2538 2692 2594 2748
rect 2594 2692 2598 2748
rect 2534 2688 2598 2692
rect 2614 2748 2678 2752
rect 2614 2692 2618 2748
rect 2618 2692 2674 2748
rect 2674 2692 2678 2748
rect 2614 2688 2678 2692
rect 3322 2748 3386 2752
rect 3322 2692 3326 2748
rect 3326 2692 3382 2748
rect 3382 2692 3386 2748
rect 3322 2688 3386 2692
rect 3402 2748 3466 2752
rect 3402 2692 3406 2748
rect 3406 2692 3462 2748
rect 3462 2692 3466 2748
rect 3402 2688 3466 2692
rect 3482 2748 3546 2752
rect 3482 2692 3486 2748
rect 3486 2692 3542 2748
rect 3542 2692 3546 2748
rect 3482 2688 3546 2692
rect 3562 2748 3626 2752
rect 3562 2692 3566 2748
rect 3566 2692 3622 2748
rect 3622 2692 3626 2748
rect 3562 2688 3626 2692
rect 4270 2748 4334 2752
rect 4270 2692 4274 2748
rect 4274 2692 4330 2748
rect 4330 2692 4334 2748
rect 4270 2688 4334 2692
rect 4350 2748 4414 2752
rect 4350 2692 4354 2748
rect 4354 2692 4410 2748
rect 4410 2692 4414 2748
rect 4350 2688 4414 2692
rect 4430 2748 4494 2752
rect 4430 2692 4434 2748
rect 4434 2692 4490 2748
rect 4490 2692 4494 2748
rect 4430 2688 4494 2692
rect 4510 2748 4574 2752
rect 4510 2692 4514 2748
rect 4514 2692 4570 2748
rect 4570 2692 4574 2748
rect 4510 2688 4574 2692
rect 1900 2204 1964 2208
rect 1900 2148 1904 2204
rect 1904 2148 1960 2204
rect 1960 2148 1964 2204
rect 1900 2144 1964 2148
rect 1980 2204 2044 2208
rect 1980 2148 1984 2204
rect 1984 2148 2040 2204
rect 2040 2148 2044 2204
rect 1980 2144 2044 2148
rect 2060 2204 2124 2208
rect 2060 2148 2064 2204
rect 2064 2148 2120 2204
rect 2120 2148 2124 2204
rect 2060 2144 2124 2148
rect 2140 2204 2204 2208
rect 2140 2148 2144 2204
rect 2144 2148 2200 2204
rect 2200 2148 2204 2204
rect 2140 2144 2204 2148
rect 2848 2204 2912 2208
rect 2848 2148 2852 2204
rect 2852 2148 2908 2204
rect 2908 2148 2912 2204
rect 2848 2144 2912 2148
rect 2928 2204 2992 2208
rect 2928 2148 2932 2204
rect 2932 2148 2988 2204
rect 2988 2148 2992 2204
rect 2928 2144 2992 2148
rect 3008 2204 3072 2208
rect 3008 2148 3012 2204
rect 3012 2148 3068 2204
rect 3068 2148 3072 2204
rect 3008 2144 3072 2148
rect 3088 2204 3152 2208
rect 3088 2148 3092 2204
rect 3092 2148 3148 2204
rect 3148 2148 3152 2204
rect 3088 2144 3152 2148
rect 3796 2204 3860 2208
rect 3796 2148 3800 2204
rect 3800 2148 3856 2204
rect 3856 2148 3860 2204
rect 3796 2144 3860 2148
rect 3876 2204 3940 2208
rect 3876 2148 3880 2204
rect 3880 2148 3936 2204
rect 3936 2148 3940 2204
rect 3876 2144 3940 2148
rect 3956 2204 4020 2208
rect 3956 2148 3960 2204
rect 3960 2148 4016 2204
rect 4016 2148 4020 2204
rect 3956 2144 4020 2148
rect 4036 2204 4100 2208
rect 4036 2148 4040 2204
rect 4040 2148 4096 2204
rect 4096 2148 4100 2204
rect 4036 2144 4100 2148
rect 1426 1660 1490 1664
rect 1426 1604 1430 1660
rect 1430 1604 1486 1660
rect 1486 1604 1490 1660
rect 1426 1600 1490 1604
rect 1506 1660 1570 1664
rect 1506 1604 1510 1660
rect 1510 1604 1566 1660
rect 1566 1604 1570 1660
rect 1506 1600 1570 1604
rect 1586 1660 1650 1664
rect 1586 1604 1590 1660
rect 1590 1604 1646 1660
rect 1646 1604 1650 1660
rect 1586 1600 1650 1604
rect 1666 1660 1730 1664
rect 1666 1604 1670 1660
rect 1670 1604 1726 1660
rect 1726 1604 1730 1660
rect 1666 1600 1730 1604
rect 2374 1660 2438 1664
rect 2374 1604 2378 1660
rect 2378 1604 2434 1660
rect 2434 1604 2438 1660
rect 2374 1600 2438 1604
rect 2454 1660 2518 1664
rect 2454 1604 2458 1660
rect 2458 1604 2514 1660
rect 2514 1604 2518 1660
rect 2454 1600 2518 1604
rect 2534 1660 2598 1664
rect 2534 1604 2538 1660
rect 2538 1604 2594 1660
rect 2594 1604 2598 1660
rect 2534 1600 2598 1604
rect 2614 1660 2678 1664
rect 2614 1604 2618 1660
rect 2618 1604 2674 1660
rect 2674 1604 2678 1660
rect 2614 1600 2678 1604
rect 3322 1660 3386 1664
rect 3322 1604 3326 1660
rect 3326 1604 3382 1660
rect 3382 1604 3386 1660
rect 3322 1600 3386 1604
rect 3402 1660 3466 1664
rect 3402 1604 3406 1660
rect 3406 1604 3462 1660
rect 3462 1604 3466 1660
rect 3402 1600 3466 1604
rect 3482 1660 3546 1664
rect 3482 1604 3486 1660
rect 3486 1604 3542 1660
rect 3542 1604 3546 1660
rect 3482 1600 3546 1604
rect 3562 1660 3626 1664
rect 3562 1604 3566 1660
rect 3566 1604 3622 1660
rect 3622 1604 3626 1660
rect 3562 1600 3626 1604
rect 4270 1660 4334 1664
rect 4270 1604 4274 1660
rect 4274 1604 4330 1660
rect 4330 1604 4334 1660
rect 4270 1600 4334 1604
rect 4350 1660 4414 1664
rect 4350 1604 4354 1660
rect 4354 1604 4410 1660
rect 4410 1604 4414 1660
rect 4350 1600 4414 1604
rect 4430 1660 4494 1664
rect 4430 1604 4434 1660
rect 4434 1604 4490 1660
rect 4490 1604 4494 1660
rect 4430 1600 4494 1604
rect 4510 1660 4574 1664
rect 4510 1604 4514 1660
rect 4514 1604 4570 1660
rect 4570 1604 4574 1660
rect 4510 1600 4574 1604
rect 1900 1116 1964 1120
rect 1900 1060 1904 1116
rect 1904 1060 1960 1116
rect 1960 1060 1964 1116
rect 1900 1056 1964 1060
rect 1980 1116 2044 1120
rect 1980 1060 1984 1116
rect 1984 1060 2040 1116
rect 2040 1060 2044 1116
rect 1980 1056 2044 1060
rect 2060 1116 2124 1120
rect 2060 1060 2064 1116
rect 2064 1060 2120 1116
rect 2120 1060 2124 1116
rect 2060 1056 2124 1060
rect 2140 1116 2204 1120
rect 2140 1060 2144 1116
rect 2144 1060 2200 1116
rect 2200 1060 2204 1116
rect 2140 1056 2204 1060
rect 2848 1116 2912 1120
rect 2848 1060 2852 1116
rect 2852 1060 2908 1116
rect 2908 1060 2912 1116
rect 2848 1056 2912 1060
rect 2928 1116 2992 1120
rect 2928 1060 2932 1116
rect 2932 1060 2988 1116
rect 2988 1060 2992 1116
rect 2928 1056 2992 1060
rect 3008 1116 3072 1120
rect 3008 1060 3012 1116
rect 3012 1060 3068 1116
rect 3068 1060 3072 1116
rect 3008 1056 3072 1060
rect 3088 1116 3152 1120
rect 3088 1060 3092 1116
rect 3092 1060 3148 1116
rect 3148 1060 3152 1116
rect 3088 1056 3152 1060
rect 3796 1116 3860 1120
rect 3796 1060 3800 1116
rect 3800 1060 3856 1116
rect 3856 1060 3860 1116
rect 3796 1056 3860 1060
rect 3876 1116 3940 1120
rect 3876 1060 3880 1116
rect 3880 1060 3936 1116
rect 3936 1060 3940 1116
rect 3876 1056 3940 1060
rect 3956 1116 4020 1120
rect 3956 1060 3960 1116
rect 3960 1060 4016 1116
rect 4016 1060 4020 1116
rect 3956 1056 4020 1060
rect 4036 1116 4100 1120
rect 4036 1060 4040 1116
rect 4040 1060 4096 1116
rect 4096 1060 4100 1116
rect 4036 1056 4100 1060
<< metal4 >>
rect 1418 22336 1738 22896
rect 1418 22272 1426 22336
rect 1490 22272 1506 22336
rect 1570 22272 1586 22336
rect 1650 22272 1666 22336
rect 1730 22272 1738 22336
rect 1418 21248 1738 22272
rect 1418 21184 1426 21248
rect 1490 21184 1506 21248
rect 1570 21184 1586 21248
rect 1650 21184 1666 21248
rect 1730 21184 1738 21248
rect 1418 20160 1738 21184
rect 1418 20096 1426 20160
rect 1490 20096 1506 20160
rect 1570 20096 1586 20160
rect 1650 20096 1666 20160
rect 1730 20096 1738 20160
rect 1418 19072 1738 20096
rect 1418 19008 1426 19072
rect 1490 19008 1506 19072
rect 1570 19008 1586 19072
rect 1650 19008 1666 19072
rect 1730 19008 1738 19072
rect 1418 17984 1738 19008
rect 1418 17920 1426 17984
rect 1490 17920 1506 17984
rect 1570 17920 1586 17984
rect 1650 17920 1666 17984
rect 1730 17920 1738 17984
rect 1418 16896 1738 17920
rect 1418 16832 1426 16896
rect 1490 16832 1506 16896
rect 1570 16832 1586 16896
rect 1650 16832 1666 16896
rect 1730 16832 1738 16896
rect 1418 15808 1738 16832
rect 1418 15744 1426 15808
rect 1490 15744 1506 15808
rect 1570 15744 1586 15808
rect 1650 15744 1666 15808
rect 1730 15744 1738 15808
rect 1418 14720 1738 15744
rect 1418 14656 1426 14720
rect 1490 14656 1506 14720
rect 1570 14656 1586 14720
rect 1650 14656 1666 14720
rect 1730 14656 1738 14720
rect 1418 13632 1738 14656
rect 1418 13568 1426 13632
rect 1490 13568 1506 13632
rect 1570 13568 1586 13632
rect 1650 13568 1666 13632
rect 1730 13568 1738 13632
rect 1418 12544 1738 13568
rect 1418 12480 1426 12544
rect 1490 12480 1506 12544
rect 1570 12480 1586 12544
rect 1650 12480 1666 12544
rect 1730 12480 1738 12544
rect 1418 11456 1738 12480
rect 1418 11392 1426 11456
rect 1490 11392 1506 11456
rect 1570 11392 1586 11456
rect 1650 11392 1666 11456
rect 1730 11392 1738 11456
rect 1418 10368 1738 11392
rect 1418 10304 1426 10368
rect 1490 10304 1506 10368
rect 1570 10304 1586 10368
rect 1650 10304 1666 10368
rect 1730 10304 1738 10368
rect 1418 9280 1738 10304
rect 1418 9216 1426 9280
rect 1490 9216 1506 9280
rect 1570 9216 1586 9280
rect 1650 9216 1666 9280
rect 1730 9216 1738 9280
rect 1418 8192 1738 9216
rect 1418 8128 1426 8192
rect 1490 8128 1506 8192
rect 1570 8128 1586 8192
rect 1650 8128 1666 8192
rect 1730 8128 1738 8192
rect 1418 7104 1738 8128
rect 1418 7040 1426 7104
rect 1490 7040 1506 7104
rect 1570 7040 1586 7104
rect 1650 7040 1666 7104
rect 1730 7040 1738 7104
rect 1418 6016 1738 7040
rect 1418 5952 1426 6016
rect 1490 5952 1506 6016
rect 1570 5952 1586 6016
rect 1650 5952 1666 6016
rect 1730 5952 1738 6016
rect 1418 4928 1738 5952
rect 1418 4864 1426 4928
rect 1490 4864 1506 4928
rect 1570 4864 1586 4928
rect 1650 4864 1666 4928
rect 1730 4864 1738 4928
rect 1418 3840 1738 4864
rect 1418 3776 1426 3840
rect 1490 3776 1506 3840
rect 1570 3776 1586 3840
rect 1650 3776 1666 3840
rect 1730 3776 1738 3840
rect 1418 2752 1738 3776
rect 1418 2688 1426 2752
rect 1490 2688 1506 2752
rect 1570 2688 1586 2752
rect 1650 2688 1666 2752
rect 1730 2688 1738 2752
rect 1418 1664 1738 2688
rect 1418 1600 1426 1664
rect 1490 1600 1506 1664
rect 1570 1600 1586 1664
rect 1650 1600 1666 1664
rect 1730 1600 1738 1664
rect 1418 1040 1738 1600
rect 1892 22880 2212 22896
rect 1892 22816 1900 22880
rect 1964 22816 1980 22880
rect 2044 22816 2060 22880
rect 2124 22816 2140 22880
rect 2204 22816 2212 22880
rect 1892 21792 2212 22816
rect 1892 21728 1900 21792
rect 1964 21728 1980 21792
rect 2044 21728 2060 21792
rect 2124 21728 2140 21792
rect 2204 21728 2212 21792
rect 1892 20704 2212 21728
rect 1892 20640 1900 20704
rect 1964 20640 1980 20704
rect 2044 20640 2060 20704
rect 2124 20640 2140 20704
rect 2204 20640 2212 20704
rect 1892 19616 2212 20640
rect 1892 19552 1900 19616
rect 1964 19552 1980 19616
rect 2044 19552 2060 19616
rect 2124 19552 2140 19616
rect 2204 19552 2212 19616
rect 1892 18528 2212 19552
rect 1892 18464 1900 18528
rect 1964 18464 1980 18528
rect 2044 18464 2060 18528
rect 2124 18464 2140 18528
rect 2204 18464 2212 18528
rect 1892 17440 2212 18464
rect 1892 17376 1900 17440
rect 1964 17376 1980 17440
rect 2044 17376 2060 17440
rect 2124 17376 2140 17440
rect 2204 17376 2212 17440
rect 1892 16352 2212 17376
rect 1892 16288 1900 16352
rect 1964 16288 1980 16352
rect 2044 16288 2060 16352
rect 2124 16288 2140 16352
rect 2204 16288 2212 16352
rect 1892 15264 2212 16288
rect 1892 15200 1900 15264
rect 1964 15200 1980 15264
rect 2044 15200 2060 15264
rect 2124 15200 2140 15264
rect 2204 15200 2212 15264
rect 1892 14176 2212 15200
rect 1892 14112 1900 14176
rect 1964 14112 1980 14176
rect 2044 14112 2060 14176
rect 2124 14112 2140 14176
rect 2204 14112 2212 14176
rect 1892 13088 2212 14112
rect 1892 13024 1900 13088
rect 1964 13024 1980 13088
rect 2044 13024 2060 13088
rect 2124 13024 2140 13088
rect 2204 13024 2212 13088
rect 1892 12000 2212 13024
rect 1892 11936 1900 12000
rect 1964 11936 1980 12000
rect 2044 11936 2060 12000
rect 2124 11936 2140 12000
rect 2204 11936 2212 12000
rect 1892 10912 2212 11936
rect 1892 10848 1900 10912
rect 1964 10848 1980 10912
rect 2044 10848 2060 10912
rect 2124 10848 2140 10912
rect 2204 10848 2212 10912
rect 1892 9824 2212 10848
rect 1892 9760 1900 9824
rect 1964 9760 1980 9824
rect 2044 9760 2060 9824
rect 2124 9760 2140 9824
rect 2204 9760 2212 9824
rect 1892 8736 2212 9760
rect 1892 8672 1900 8736
rect 1964 8672 1980 8736
rect 2044 8672 2060 8736
rect 2124 8672 2140 8736
rect 2204 8672 2212 8736
rect 1892 7648 2212 8672
rect 1892 7584 1900 7648
rect 1964 7584 1980 7648
rect 2044 7584 2060 7648
rect 2124 7584 2140 7648
rect 2204 7584 2212 7648
rect 1892 6560 2212 7584
rect 1892 6496 1900 6560
rect 1964 6496 1980 6560
rect 2044 6496 2060 6560
rect 2124 6496 2140 6560
rect 2204 6496 2212 6560
rect 1892 5472 2212 6496
rect 1892 5408 1900 5472
rect 1964 5408 1980 5472
rect 2044 5408 2060 5472
rect 2124 5408 2140 5472
rect 2204 5408 2212 5472
rect 1892 4384 2212 5408
rect 1892 4320 1900 4384
rect 1964 4320 1980 4384
rect 2044 4320 2060 4384
rect 2124 4320 2140 4384
rect 2204 4320 2212 4384
rect 1892 3296 2212 4320
rect 1892 3232 1900 3296
rect 1964 3232 1980 3296
rect 2044 3232 2060 3296
rect 2124 3232 2140 3296
rect 2204 3232 2212 3296
rect 1892 2208 2212 3232
rect 1892 2144 1900 2208
rect 1964 2144 1980 2208
rect 2044 2144 2060 2208
rect 2124 2144 2140 2208
rect 2204 2144 2212 2208
rect 1892 1120 2212 2144
rect 1892 1056 1900 1120
rect 1964 1056 1980 1120
rect 2044 1056 2060 1120
rect 2124 1056 2140 1120
rect 2204 1056 2212 1120
rect 1892 1040 2212 1056
rect 2366 22336 2686 22896
rect 2366 22272 2374 22336
rect 2438 22272 2454 22336
rect 2518 22272 2534 22336
rect 2598 22272 2614 22336
rect 2678 22272 2686 22336
rect 2366 21248 2686 22272
rect 2366 21184 2374 21248
rect 2438 21184 2454 21248
rect 2518 21184 2534 21248
rect 2598 21184 2614 21248
rect 2678 21184 2686 21248
rect 2366 20160 2686 21184
rect 2366 20096 2374 20160
rect 2438 20096 2454 20160
rect 2518 20096 2534 20160
rect 2598 20096 2614 20160
rect 2678 20096 2686 20160
rect 2366 19072 2686 20096
rect 2366 19008 2374 19072
rect 2438 19008 2454 19072
rect 2518 19008 2534 19072
rect 2598 19008 2614 19072
rect 2678 19008 2686 19072
rect 2366 17984 2686 19008
rect 2366 17920 2374 17984
rect 2438 17920 2454 17984
rect 2518 17920 2534 17984
rect 2598 17920 2614 17984
rect 2678 17920 2686 17984
rect 2366 16896 2686 17920
rect 2366 16832 2374 16896
rect 2438 16832 2454 16896
rect 2518 16832 2534 16896
rect 2598 16832 2614 16896
rect 2678 16832 2686 16896
rect 2366 15808 2686 16832
rect 2366 15744 2374 15808
rect 2438 15744 2454 15808
rect 2518 15744 2534 15808
rect 2598 15744 2614 15808
rect 2678 15744 2686 15808
rect 2366 14720 2686 15744
rect 2366 14656 2374 14720
rect 2438 14656 2454 14720
rect 2518 14656 2534 14720
rect 2598 14656 2614 14720
rect 2678 14656 2686 14720
rect 2366 13632 2686 14656
rect 2366 13568 2374 13632
rect 2438 13568 2454 13632
rect 2518 13568 2534 13632
rect 2598 13568 2614 13632
rect 2678 13568 2686 13632
rect 2366 12544 2686 13568
rect 2366 12480 2374 12544
rect 2438 12480 2454 12544
rect 2518 12480 2534 12544
rect 2598 12480 2614 12544
rect 2678 12480 2686 12544
rect 2366 11456 2686 12480
rect 2366 11392 2374 11456
rect 2438 11392 2454 11456
rect 2518 11392 2534 11456
rect 2598 11392 2614 11456
rect 2678 11392 2686 11456
rect 2366 10368 2686 11392
rect 2366 10304 2374 10368
rect 2438 10304 2454 10368
rect 2518 10304 2534 10368
rect 2598 10304 2614 10368
rect 2678 10304 2686 10368
rect 2366 9280 2686 10304
rect 2366 9216 2374 9280
rect 2438 9216 2454 9280
rect 2518 9216 2534 9280
rect 2598 9216 2614 9280
rect 2678 9216 2686 9280
rect 2366 8192 2686 9216
rect 2366 8128 2374 8192
rect 2438 8128 2454 8192
rect 2518 8128 2534 8192
rect 2598 8128 2614 8192
rect 2678 8128 2686 8192
rect 2366 7104 2686 8128
rect 2366 7040 2374 7104
rect 2438 7040 2454 7104
rect 2518 7040 2534 7104
rect 2598 7040 2614 7104
rect 2678 7040 2686 7104
rect 2366 6016 2686 7040
rect 2366 5952 2374 6016
rect 2438 5952 2454 6016
rect 2518 5952 2534 6016
rect 2598 5952 2614 6016
rect 2678 5952 2686 6016
rect 2366 4928 2686 5952
rect 2366 4864 2374 4928
rect 2438 4864 2454 4928
rect 2518 4864 2534 4928
rect 2598 4864 2614 4928
rect 2678 4864 2686 4928
rect 2366 3840 2686 4864
rect 2366 3776 2374 3840
rect 2438 3776 2454 3840
rect 2518 3776 2534 3840
rect 2598 3776 2614 3840
rect 2678 3776 2686 3840
rect 2366 2752 2686 3776
rect 2366 2688 2374 2752
rect 2438 2688 2454 2752
rect 2518 2688 2534 2752
rect 2598 2688 2614 2752
rect 2678 2688 2686 2752
rect 2366 1664 2686 2688
rect 2366 1600 2374 1664
rect 2438 1600 2454 1664
rect 2518 1600 2534 1664
rect 2598 1600 2614 1664
rect 2678 1600 2686 1664
rect 2366 1040 2686 1600
rect 2840 22880 3160 22896
rect 2840 22816 2848 22880
rect 2912 22816 2928 22880
rect 2992 22816 3008 22880
rect 3072 22816 3088 22880
rect 3152 22816 3160 22880
rect 2840 21792 3160 22816
rect 2840 21728 2848 21792
rect 2912 21728 2928 21792
rect 2992 21728 3008 21792
rect 3072 21728 3088 21792
rect 3152 21728 3160 21792
rect 2840 20704 3160 21728
rect 2840 20640 2848 20704
rect 2912 20640 2928 20704
rect 2992 20640 3008 20704
rect 3072 20640 3088 20704
rect 3152 20640 3160 20704
rect 2840 19616 3160 20640
rect 2840 19552 2848 19616
rect 2912 19552 2928 19616
rect 2992 19552 3008 19616
rect 3072 19552 3088 19616
rect 3152 19552 3160 19616
rect 2840 18528 3160 19552
rect 2840 18464 2848 18528
rect 2912 18464 2928 18528
rect 2992 18464 3008 18528
rect 3072 18464 3088 18528
rect 3152 18464 3160 18528
rect 2840 17440 3160 18464
rect 2840 17376 2848 17440
rect 2912 17376 2928 17440
rect 2992 17376 3008 17440
rect 3072 17376 3088 17440
rect 3152 17376 3160 17440
rect 2840 16352 3160 17376
rect 2840 16288 2848 16352
rect 2912 16288 2928 16352
rect 2992 16288 3008 16352
rect 3072 16288 3088 16352
rect 3152 16288 3160 16352
rect 2840 15264 3160 16288
rect 2840 15200 2848 15264
rect 2912 15200 2928 15264
rect 2992 15200 3008 15264
rect 3072 15200 3088 15264
rect 3152 15200 3160 15264
rect 2840 14176 3160 15200
rect 2840 14112 2848 14176
rect 2912 14112 2928 14176
rect 2992 14112 3008 14176
rect 3072 14112 3088 14176
rect 3152 14112 3160 14176
rect 2840 13088 3160 14112
rect 2840 13024 2848 13088
rect 2912 13024 2928 13088
rect 2992 13024 3008 13088
rect 3072 13024 3088 13088
rect 3152 13024 3160 13088
rect 2840 12000 3160 13024
rect 2840 11936 2848 12000
rect 2912 11936 2928 12000
rect 2992 11936 3008 12000
rect 3072 11936 3088 12000
rect 3152 11936 3160 12000
rect 2840 10912 3160 11936
rect 2840 10848 2848 10912
rect 2912 10848 2928 10912
rect 2992 10848 3008 10912
rect 3072 10848 3088 10912
rect 3152 10848 3160 10912
rect 2840 9824 3160 10848
rect 2840 9760 2848 9824
rect 2912 9760 2928 9824
rect 2992 9760 3008 9824
rect 3072 9760 3088 9824
rect 3152 9760 3160 9824
rect 2840 8736 3160 9760
rect 2840 8672 2848 8736
rect 2912 8672 2928 8736
rect 2992 8672 3008 8736
rect 3072 8672 3088 8736
rect 3152 8672 3160 8736
rect 2840 7648 3160 8672
rect 2840 7584 2848 7648
rect 2912 7584 2928 7648
rect 2992 7584 3008 7648
rect 3072 7584 3088 7648
rect 3152 7584 3160 7648
rect 2840 6560 3160 7584
rect 2840 6496 2848 6560
rect 2912 6496 2928 6560
rect 2992 6496 3008 6560
rect 3072 6496 3088 6560
rect 3152 6496 3160 6560
rect 2840 5472 3160 6496
rect 2840 5408 2848 5472
rect 2912 5408 2928 5472
rect 2992 5408 3008 5472
rect 3072 5408 3088 5472
rect 3152 5408 3160 5472
rect 2840 4384 3160 5408
rect 2840 4320 2848 4384
rect 2912 4320 2928 4384
rect 2992 4320 3008 4384
rect 3072 4320 3088 4384
rect 3152 4320 3160 4384
rect 2840 3296 3160 4320
rect 2840 3232 2848 3296
rect 2912 3232 2928 3296
rect 2992 3232 3008 3296
rect 3072 3232 3088 3296
rect 3152 3232 3160 3296
rect 2840 2208 3160 3232
rect 2840 2144 2848 2208
rect 2912 2144 2928 2208
rect 2992 2144 3008 2208
rect 3072 2144 3088 2208
rect 3152 2144 3160 2208
rect 2840 1120 3160 2144
rect 2840 1056 2848 1120
rect 2912 1056 2928 1120
rect 2992 1056 3008 1120
rect 3072 1056 3088 1120
rect 3152 1056 3160 1120
rect 2840 1040 3160 1056
rect 3314 22336 3634 22896
rect 3314 22272 3322 22336
rect 3386 22272 3402 22336
rect 3466 22272 3482 22336
rect 3546 22272 3562 22336
rect 3626 22272 3634 22336
rect 3314 21248 3634 22272
rect 3314 21184 3322 21248
rect 3386 21184 3402 21248
rect 3466 21184 3482 21248
rect 3546 21184 3562 21248
rect 3626 21184 3634 21248
rect 3314 20160 3634 21184
rect 3314 20096 3322 20160
rect 3386 20096 3402 20160
rect 3466 20096 3482 20160
rect 3546 20096 3562 20160
rect 3626 20096 3634 20160
rect 3314 19072 3634 20096
rect 3314 19008 3322 19072
rect 3386 19008 3402 19072
rect 3466 19008 3482 19072
rect 3546 19008 3562 19072
rect 3626 19008 3634 19072
rect 3314 17984 3634 19008
rect 3314 17920 3322 17984
rect 3386 17920 3402 17984
rect 3466 17920 3482 17984
rect 3546 17920 3562 17984
rect 3626 17920 3634 17984
rect 3314 16896 3634 17920
rect 3314 16832 3322 16896
rect 3386 16832 3402 16896
rect 3466 16832 3482 16896
rect 3546 16832 3562 16896
rect 3626 16832 3634 16896
rect 3314 15808 3634 16832
rect 3314 15744 3322 15808
rect 3386 15744 3402 15808
rect 3466 15744 3482 15808
rect 3546 15744 3562 15808
rect 3626 15744 3634 15808
rect 3314 14720 3634 15744
rect 3314 14656 3322 14720
rect 3386 14656 3402 14720
rect 3466 14656 3482 14720
rect 3546 14656 3562 14720
rect 3626 14656 3634 14720
rect 3314 13632 3634 14656
rect 3314 13568 3322 13632
rect 3386 13568 3402 13632
rect 3466 13568 3482 13632
rect 3546 13568 3562 13632
rect 3626 13568 3634 13632
rect 3314 12544 3634 13568
rect 3314 12480 3322 12544
rect 3386 12480 3402 12544
rect 3466 12480 3482 12544
rect 3546 12480 3562 12544
rect 3626 12480 3634 12544
rect 3314 11456 3634 12480
rect 3314 11392 3322 11456
rect 3386 11392 3402 11456
rect 3466 11392 3482 11456
rect 3546 11392 3562 11456
rect 3626 11392 3634 11456
rect 3314 10368 3634 11392
rect 3314 10304 3322 10368
rect 3386 10304 3402 10368
rect 3466 10304 3482 10368
rect 3546 10304 3562 10368
rect 3626 10304 3634 10368
rect 3314 9280 3634 10304
rect 3314 9216 3322 9280
rect 3386 9216 3402 9280
rect 3466 9216 3482 9280
rect 3546 9216 3562 9280
rect 3626 9216 3634 9280
rect 3314 8192 3634 9216
rect 3314 8128 3322 8192
rect 3386 8128 3402 8192
rect 3466 8128 3482 8192
rect 3546 8128 3562 8192
rect 3626 8128 3634 8192
rect 3314 7104 3634 8128
rect 3314 7040 3322 7104
rect 3386 7040 3402 7104
rect 3466 7040 3482 7104
rect 3546 7040 3562 7104
rect 3626 7040 3634 7104
rect 3314 6016 3634 7040
rect 3314 5952 3322 6016
rect 3386 5952 3402 6016
rect 3466 5952 3482 6016
rect 3546 5952 3562 6016
rect 3626 5952 3634 6016
rect 3314 4928 3634 5952
rect 3314 4864 3322 4928
rect 3386 4864 3402 4928
rect 3466 4864 3482 4928
rect 3546 4864 3562 4928
rect 3626 4864 3634 4928
rect 3314 3840 3634 4864
rect 3314 3776 3322 3840
rect 3386 3776 3402 3840
rect 3466 3776 3482 3840
rect 3546 3776 3562 3840
rect 3626 3776 3634 3840
rect 3314 2752 3634 3776
rect 3314 2688 3322 2752
rect 3386 2688 3402 2752
rect 3466 2688 3482 2752
rect 3546 2688 3562 2752
rect 3626 2688 3634 2752
rect 3314 1664 3634 2688
rect 3314 1600 3322 1664
rect 3386 1600 3402 1664
rect 3466 1600 3482 1664
rect 3546 1600 3562 1664
rect 3626 1600 3634 1664
rect 3314 1040 3634 1600
rect 3788 22880 4108 22896
rect 3788 22816 3796 22880
rect 3860 22816 3876 22880
rect 3940 22816 3956 22880
rect 4020 22816 4036 22880
rect 4100 22816 4108 22880
rect 3788 21792 4108 22816
rect 3788 21728 3796 21792
rect 3860 21728 3876 21792
rect 3940 21728 3956 21792
rect 4020 21728 4036 21792
rect 4100 21728 4108 21792
rect 3788 20704 4108 21728
rect 3788 20640 3796 20704
rect 3860 20640 3876 20704
rect 3940 20640 3956 20704
rect 4020 20640 4036 20704
rect 4100 20640 4108 20704
rect 3788 19616 4108 20640
rect 3788 19552 3796 19616
rect 3860 19552 3876 19616
rect 3940 19552 3956 19616
rect 4020 19552 4036 19616
rect 4100 19552 4108 19616
rect 3788 18528 4108 19552
rect 3788 18464 3796 18528
rect 3860 18464 3876 18528
rect 3940 18464 3956 18528
rect 4020 18464 4036 18528
rect 4100 18464 4108 18528
rect 3788 17440 4108 18464
rect 3788 17376 3796 17440
rect 3860 17376 3876 17440
rect 3940 17376 3956 17440
rect 4020 17376 4036 17440
rect 4100 17376 4108 17440
rect 3788 16352 4108 17376
rect 3788 16288 3796 16352
rect 3860 16288 3876 16352
rect 3940 16288 3956 16352
rect 4020 16288 4036 16352
rect 4100 16288 4108 16352
rect 3788 15264 4108 16288
rect 3788 15200 3796 15264
rect 3860 15200 3876 15264
rect 3940 15200 3956 15264
rect 4020 15200 4036 15264
rect 4100 15200 4108 15264
rect 3788 14176 4108 15200
rect 3788 14112 3796 14176
rect 3860 14112 3876 14176
rect 3940 14112 3956 14176
rect 4020 14112 4036 14176
rect 4100 14112 4108 14176
rect 3788 13088 4108 14112
rect 3788 13024 3796 13088
rect 3860 13024 3876 13088
rect 3940 13024 3956 13088
rect 4020 13024 4036 13088
rect 4100 13024 4108 13088
rect 3788 12000 4108 13024
rect 3788 11936 3796 12000
rect 3860 11936 3876 12000
rect 3940 11936 3956 12000
rect 4020 11936 4036 12000
rect 4100 11936 4108 12000
rect 3788 10912 4108 11936
rect 3788 10848 3796 10912
rect 3860 10848 3876 10912
rect 3940 10848 3956 10912
rect 4020 10848 4036 10912
rect 4100 10848 4108 10912
rect 3788 9824 4108 10848
rect 3788 9760 3796 9824
rect 3860 9760 3876 9824
rect 3940 9760 3956 9824
rect 4020 9760 4036 9824
rect 4100 9760 4108 9824
rect 3788 8736 4108 9760
rect 3788 8672 3796 8736
rect 3860 8672 3876 8736
rect 3940 8672 3956 8736
rect 4020 8672 4036 8736
rect 4100 8672 4108 8736
rect 3788 7648 4108 8672
rect 3788 7584 3796 7648
rect 3860 7584 3876 7648
rect 3940 7584 3956 7648
rect 4020 7584 4036 7648
rect 4100 7584 4108 7648
rect 3788 6560 4108 7584
rect 3788 6496 3796 6560
rect 3860 6496 3876 6560
rect 3940 6496 3956 6560
rect 4020 6496 4036 6560
rect 4100 6496 4108 6560
rect 3788 5472 4108 6496
rect 3788 5408 3796 5472
rect 3860 5408 3876 5472
rect 3940 5408 3956 5472
rect 4020 5408 4036 5472
rect 4100 5408 4108 5472
rect 3788 4384 4108 5408
rect 3788 4320 3796 4384
rect 3860 4320 3876 4384
rect 3940 4320 3956 4384
rect 4020 4320 4036 4384
rect 4100 4320 4108 4384
rect 3788 3296 4108 4320
rect 3788 3232 3796 3296
rect 3860 3232 3876 3296
rect 3940 3232 3956 3296
rect 4020 3232 4036 3296
rect 4100 3232 4108 3296
rect 3788 2208 4108 3232
rect 3788 2144 3796 2208
rect 3860 2144 3876 2208
rect 3940 2144 3956 2208
rect 4020 2144 4036 2208
rect 4100 2144 4108 2208
rect 3788 1120 4108 2144
rect 3788 1056 3796 1120
rect 3860 1056 3876 1120
rect 3940 1056 3956 1120
rect 4020 1056 4036 1120
rect 4100 1056 4108 1120
rect 3788 1040 4108 1056
rect 4262 22336 4582 22896
rect 4262 22272 4270 22336
rect 4334 22272 4350 22336
rect 4414 22272 4430 22336
rect 4494 22272 4510 22336
rect 4574 22272 4582 22336
rect 4262 21248 4582 22272
rect 4262 21184 4270 21248
rect 4334 21184 4350 21248
rect 4414 21184 4430 21248
rect 4494 21184 4510 21248
rect 4574 21184 4582 21248
rect 4262 20160 4582 21184
rect 4262 20096 4270 20160
rect 4334 20096 4350 20160
rect 4414 20096 4430 20160
rect 4494 20096 4510 20160
rect 4574 20096 4582 20160
rect 4262 19072 4582 20096
rect 4262 19008 4270 19072
rect 4334 19008 4350 19072
rect 4414 19008 4430 19072
rect 4494 19008 4510 19072
rect 4574 19008 4582 19072
rect 4262 17984 4582 19008
rect 4262 17920 4270 17984
rect 4334 17920 4350 17984
rect 4414 17920 4430 17984
rect 4494 17920 4510 17984
rect 4574 17920 4582 17984
rect 4262 16896 4582 17920
rect 4262 16832 4270 16896
rect 4334 16832 4350 16896
rect 4414 16832 4430 16896
rect 4494 16832 4510 16896
rect 4574 16832 4582 16896
rect 4262 15808 4582 16832
rect 4262 15744 4270 15808
rect 4334 15744 4350 15808
rect 4414 15744 4430 15808
rect 4494 15744 4510 15808
rect 4574 15744 4582 15808
rect 4262 14720 4582 15744
rect 4262 14656 4270 14720
rect 4334 14656 4350 14720
rect 4414 14656 4430 14720
rect 4494 14656 4510 14720
rect 4574 14656 4582 14720
rect 4262 13632 4582 14656
rect 4262 13568 4270 13632
rect 4334 13568 4350 13632
rect 4414 13568 4430 13632
rect 4494 13568 4510 13632
rect 4574 13568 4582 13632
rect 4262 12544 4582 13568
rect 4262 12480 4270 12544
rect 4334 12480 4350 12544
rect 4414 12480 4430 12544
rect 4494 12480 4510 12544
rect 4574 12480 4582 12544
rect 4262 11456 4582 12480
rect 4262 11392 4270 11456
rect 4334 11392 4350 11456
rect 4414 11392 4430 11456
rect 4494 11392 4510 11456
rect 4574 11392 4582 11456
rect 4262 10368 4582 11392
rect 4262 10304 4270 10368
rect 4334 10304 4350 10368
rect 4414 10304 4430 10368
rect 4494 10304 4510 10368
rect 4574 10304 4582 10368
rect 4262 9280 4582 10304
rect 4262 9216 4270 9280
rect 4334 9216 4350 9280
rect 4414 9216 4430 9280
rect 4494 9216 4510 9280
rect 4574 9216 4582 9280
rect 4262 8192 4582 9216
rect 4262 8128 4270 8192
rect 4334 8128 4350 8192
rect 4414 8128 4430 8192
rect 4494 8128 4510 8192
rect 4574 8128 4582 8192
rect 4262 7104 4582 8128
rect 4262 7040 4270 7104
rect 4334 7040 4350 7104
rect 4414 7040 4430 7104
rect 4494 7040 4510 7104
rect 4574 7040 4582 7104
rect 4262 6016 4582 7040
rect 4262 5952 4270 6016
rect 4334 5952 4350 6016
rect 4414 5952 4430 6016
rect 4494 5952 4510 6016
rect 4574 5952 4582 6016
rect 4262 4928 4582 5952
rect 4262 4864 4270 4928
rect 4334 4864 4350 4928
rect 4414 4864 4430 4928
rect 4494 4864 4510 4928
rect 4574 4864 4582 4928
rect 4262 3840 4582 4864
rect 4262 3776 4270 3840
rect 4334 3776 4350 3840
rect 4414 3776 4430 3840
rect 4494 3776 4510 3840
rect 4574 3776 4582 3840
rect 4262 2752 4582 3776
rect 4262 2688 4270 2752
rect 4334 2688 4350 2752
rect 4414 2688 4430 2752
rect 4494 2688 4510 2752
rect 4574 2688 4582 2752
rect 4262 1664 4582 2688
rect 4262 1600 4270 1664
rect 4334 1600 4350 1664
rect 4414 1600 4430 1664
rect 4494 1600 4510 1664
rect 4574 1600 4582 1664
rect 4262 1040 4582 1600
use sky130_ef_sc_hd__decap_12  FILLER_0_3 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp 1649977179
transform 1 0 4508 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_35 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4324 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_37
timestamp 1649977179
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_35
timestamp 1649977179
transform 1 0 4324 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_37
timestamp 1649977179
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_35
timestamp 1649977179
transform 1 0 4324 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6
timestamp 1649977179
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_18
timestamp 1649977179
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_37
timestamp 1649977179
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_35
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_37
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_11
timestamp 1649977179
transform 1 0 2116 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_19
timestamp 1649977179
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_34
timestamp 1649977179
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_37
timestamp 1649977179
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_15 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_21
timestamp 1649977179
transform 1 0 3036 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 1649977179
transform 1 0 4232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_6
timestamp 1649977179
transform 1 0 1656 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_37
timestamp 1649977179
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_18
timestamp 1649977179
transform 1 0 2760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_34
timestamp 1649977179
transform 1 0 4232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1649977179
transform 1 0 2116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_32
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_11
timestamp 1649977179
transform 1 0 2116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_33
timestamp 1649977179
transform 1 0 4140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_37
timestamp 1649977179
transform 1 0 4508 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_32
timestamp 1649977179
transform 1 0 4048 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_6
timestamp 1649977179
transform 1 0 1656 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_34
timestamp 1649977179
transform 1 0 4232 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1649977179
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_34
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1649977179
transform 1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_34
timestamp 1649977179
transform 1 0 4232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_34
timestamp 1649977179
transform 1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_9
timestamp 1649977179
transform 1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_34
timestamp 1649977179
transform 1 0 4232 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1649977179
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_34
timestamp 1649977179
transform 1 0 4232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1649977179
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_34
timestamp 1649977179
transform 1 0 4232 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_34
timestamp 1649977179
transform 1 0 4232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_9
timestamp 1649977179
transform 1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_34
timestamp 1649977179
transform 1 0 4232 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_34
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_23
timestamp 1649977179
transform 1 0 3220 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_34
timestamp 1649977179
transform 1 0 4232 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_37
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_12
timestamp 1649977179
transform 1 0 2208 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_24
timestamp 1649977179
transform 1 0 3312 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1649977179
transform 1 0 4416 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_9
timestamp 1649977179
transform 1 0 1932 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1649977179
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_34
timestamp 1649977179
transform 1 0 4232 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_35
timestamp 1649977179
transform 1 0 4324 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_34
timestamp 1649977179
transform 1 0 4232 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_35
timestamp 1649977179
transform 1 0 4324 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_37
timestamp 1649977179
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1649977179
transform 1 0 4232 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_37
timestamp 1649977179
transform 1 0 4508 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_35
timestamp 1649977179
transform 1 0 4324 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_34
timestamp 1649977179
transform 1 0 4232 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_29
timestamp 1649977179
transform 1 0 3772 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1649977179
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 4876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 4876 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 4876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 4876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 4876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 4876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 4876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 4876 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 4876 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 4876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 4876 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 4876 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 4876 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 4876 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 4876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 4876 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 4876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 4876 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 4876 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 3680 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 3956 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 3956 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform 1 0 3956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 3956 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 3956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input_buf_clk shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlxtp_1  latch\[0\] shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3128 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[1\]
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[2\]
timestamp 1649977179
transform 1 0 2208 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[3\]
timestamp 1649977179
transform 1 0 3128 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[4\]
timestamp 1649977179
transform 1 0 2208 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[5\]
timestamp 1649977179
transform 1 0 3128 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[6\]
timestamp 1649977179
transform 1 0 2208 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  latch\[7\]
timestamp 1649977179
transform 1 0 2208 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  out_flop_16 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  out_flop shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2392 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  output_buffers\[0\] shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output_buffers\[1\]
timestamp 1649977179
transform -1 0 1932 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output_buffers\[2\]
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output_buffers\[3\]
timestamp 1649977179
transform -1 0 1932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  repeater12
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater13
timestamp 1649977179
transform -1 0 4048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater14
timestamp 1649977179
transform -1 0 4232 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater15 shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[0\] shuttle7/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2208 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[1\]
timestamp 1649977179
transform -1 0 3312 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[2\]
timestamp 1649977179
transform -1 0 4232 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[3\]
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[4\]
timestamp 1649977179
transform -1 0 4232 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[5\]
timestamp 1649977179
transform 1 0 2300 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[6\]
timestamp 1649977179
transform -1 0 3312 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  scan_flop\[7\]
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1970 592
<< labels >>
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 clk_in
port 0 nsew signal input
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 clk_out
port 1 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 data_in
port 2 nsew signal input
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 data_out
port 3 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 latch_enable_in
port 4 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 latch_enable_out
port 5 nsew signal tristate
flabel metal3 s 5200 688 6000 808 0 FreeSans 480 0 0 0 module_data_in[0]
port 6 nsew signal tristate
flabel metal3 s 5200 2184 6000 2304 0 FreeSans 480 0 0 0 module_data_in[1]
port 7 nsew signal tristate
flabel metal3 s 5200 3680 6000 3800 0 FreeSans 480 0 0 0 module_data_in[2]
port 8 nsew signal tristate
flabel metal3 s 5200 5176 6000 5296 0 FreeSans 480 0 0 0 module_data_in[3]
port 9 nsew signal tristate
flabel metal3 s 5200 6672 6000 6792 0 FreeSans 480 0 0 0 module_data_in[4]
port 10 nsew signal tristate
flabel metal3 s 5200 8168 6000 8288 0 FreeSans 480 0 0 0 module_data_in[5]
port 11 nsew signal tristate
flabel metal3 s 5200 9664 6000 9784 0 FreeSans 480 0 0 0 module_data_in[6]
port 12 nsew signal tristate
flabel metal3 s 5200 11160 6000 11280 0 FreeSans 480 0 0 0 module_data_in[7]
port 13 nsew signal tristate
flabel metal3 s 5200 12656 6000 12776 0 FreeSans 480 0 0 0 module_data_out[0]
port 14 nsew signal input
flabel metal3 s 5200 14152 6000 14272 0 FreeSans 480 0 0 0 module_data_out[1]
port 15 nsew signal input
flabel metal3 s 5200 15648 6000 15768 0 FreeSans 480 0 0 0 module_data_out[2]
port 16 nsew signal input
flabel metal3 s 5200 17144 6000 17264 0 FreeSans 480 0 0 0 module_data_out[3]
port 17 nsew signal input
flabel metal3 s 5200 18640 6000 18760 0 FreeSans 480 0 0 0 module_data_out[4]
port 18 nsew signal input
flabel metal3 s 5200 20136 6000 20256 0 FreeSans 480 0 0 0 module_data_out[5]
port 19 nsew signal input
flabel metal3 s 5200 21632 6000 21752 0 FreeSans 480 0 0 0 module_data_out[6]
port 20 nsew signal input
flabel metal3 s 5200 23128 6000 23248 0 FreeSans 480 0 0 0 module_data_out[7]
port 21 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 scan_select_in
port 22 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 scan_select_out
port 23 nsew signal tristate
flabel metal4 s 1418 1040 1738 22896 0 FreeSans 1920 90 0 0 vccd1
port 24 nsew power bidirectional
flabel metal4 s 2366 1040 2686 22896 0 FreeSans 1920 90 0 0 vccd1
port 24 nsew power bidirectional
flabel metal4 s 3314 1040 3634 22896 0 FreeSans 1920 90 0 0 vccd1
port 24 nsew power bidirectional
flabel metal4 s 4262 1040 4582 22896 0 FreeSans 1920 90 0 0 vccd1
port 24 nsew power bidirectional
flabel metal4 s 1892 1040 2212 22896 0 FreeSans 1920 90 0 0 vssd1
port 25 nsew ground bidirectional
flabel metal4 s 2840 1040 3160 22896 0 FreeSans 1920 90 0 0 vssd1
port 25 nsew ground bidirectional
flabel metal4 s 3788 1040 4108 22896 0 FreeSans 1920 90 0 0 vssd1
port 25 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 6000 24000
<< end >>
