/* Automatically generated from https://wokwi.com/projects/347592305412145748 */

`default_nettype none

module user_module_347592305412145748(
  input [7:0] io_in,
  output [7:0] io_out
);
  wire net1 = io_in[0];
  wire net2 = io_in[1];
  wire net3 = io_in[2];
  wire net4 = io_in[3];
  wire net5 = io_in[4];
  wire net6 = io_in[5];
  wire net7 = io_in[6];
  wire net8 = io_in[7];
  wire net9;
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14 = 1'b0;
  wire net15 = 1'b1;
  wire net16 = 1'b1;
  wire net17;
  wire net18;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138 = 1'b0;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284;
  wire net285;
  wire net286;
  wire net287;
  wire net288;
  wire net289;
  wire net290;
  wire net291;
  wire net292;
  wire net293;
  wire net294;
  wire net295;
  wire net296;
  wire net297;
  wire net298;
  wire net299;
  wire net300;
  wire net301;
  wire net302;
  wire net303;
  wire net304;
  wire net305;
  wire net306;
  wire net307;
  wire net308;
  wire net309;
  wire net310;
  wire net311;
  wire net312;
  wire net313;
  wire net314;
  wire net315;
  wire net316;
  wire net317;
  wire net318;
  wire net319;
  wire net320;
  wire net321;
  wire net322;
  wire net323;
  wire net324;
  wire net325;
  wire net326;
  wire net327;
  wire net328;
  wire net329;
  wire net330;
  wire net331;
  wire net332;
  wire net333;
  wire net334;
  wire net335;
  wire net336;
  wire net337;
  wire net338;
  wire net339;
  wire net340;
  wire net341;
  wire net342;
  wire net343;
  wire net344;
  wire net345;
  wire net346;
  wire net347;
  wire net348;
  wire net349;
  wire net350;
  wire net351;
  wire net352;
  wire net353;
  wire net354;
  wire net355;
  wire net356;
  wire net357;
  wire net358;
  wire net359;
  wire net360;
  wire net361;
  wire net362;
  wire net363;
  wire net364;
  wire net365;
  wire net366;
  wire net367;
  wire net368;
  wire net369;
  wire net370;
  wire net371;
  wire net372;
  wire net373;
  wire net374;
  wire net375;
  wire net376;
  wire net377;
  wire net378;
  wire net379;
  wire net380;
  wire net381;
  wire net382;
  wire net383;
  wire net384;
  wire net385;
  wire net386;
  wire net387;
  wire net388;
  wire net389;
  wire net390;
  wire net391;
  wire net392;
  wire net393;
  wire net394;
  wire net395;
  wire net396;
  wire net397;
  wire net398;
  wire net399;
  wire net400;
  wire net401;
  wire net402;
  wire net403;
  wire net404;
  wire net405;
  wire net406;
  wire net407;
  wire net408;
  wire net409;
  wire net410;
  wire net411;
  wire net412;
  wire net413;
  wire net414;
  wire net415;
  wire net416;
  wire net417;
  wire net418;
  wire net419;
  wire net420;
  wire net421;
  wire net422;
  wire net423;
  wire net424;
  wire net425;
  wire net426;
  wire net427;
  wire net428;
  wire net429;
  wire net430;
  wire net431;
  wire net432;
  wire net433;
  wire net434;
  wire net435;
  wire net436;
  wire net437;
  wire net438;
  wire net439;
  wire net440;
  wire net441;
  wire net442;
  wire net443;
  wire net444;
  wire net445;
  wire net446;
  wire net447;
  wire net448;
  wire net449;
  wire net450;
  wire net451;
  wire net452;
  wire net453;
  wire net454;
  wire net455;
  wire net456;
  wire net457;
  wire net458;
  wire net459;
  wire net460;
  wire net461;
  wire net462;
  wire net463;
  wire net464;
  wire net465;
  wire net466;
  wire net467;
  wire net468;
  wire net469;
  wire net470;
  wire net471;
  wire net472;
  wire net473;

  assign io_out[0] = net9;
  assign io_out[1] = net10;
  assign io_out[2] = net11;
  assign io_out[3] = net12;
  assign io_out[4] = net6;
  assign io_out[5] = net5;
  assign io_out[7] = net13;

  dff_cell flipflop10 (
    .d (net17),
    .clk (net13),
    .q (net9)
  );
  xor_cell gate18 (
    .a (net9),
    .b (net18),
    .out (net17)
  );
  buffer_cell gate22 (
    .in (net19),
    .out (net20)
  );
  buffer_cell gate23 (
    .in (net21),
    .out (net22)
  );
  and_cell gate24 (
    .a (net23),
    .b (net24),
    .out (net25)
  );
  and_cell gate25 (
    .a (net25),
    .b (net26),
    .out (net27)
  );
  and_cell gate26 (
    .a (net20),
    .b (net28),
    .out (net29)
  );
  and_cell gate27 (
    .a (net29),
    .b (net26),
    .out (net30)
  );
  and_cell gate28 (
    .a (net31),
    .b (net23),
    .out (net32)
  );
  and_cell gate29 (
    .a (net32),
    .b (net28),
    .out (net33)
  );
  and_cell gate30 (
    .a (net33),
    .b (net34),
    .out (net35)
  );
  and_cell gate31 (
    .a (net31),
    .b (net20),
    .out (net36)
  );
  and_cell gate32 (
    .a (net36),
    .b (net24),
    .out (net37)
  );
  and_cell gate33 (
    .a (net37),
    .b (net38),
    .out (net39)
  );
  and_cell gate34 (
    .a (net22),
    .b (net23),
    .out (net40)
  );
  and_cell gate35 (
    .a (net40),
    .b (net28),
    .out (net41)
  );
  and_cell gate36 (
    .a (net41),
    .b (net38),
    .out (net42)
  );
  and_cell gate37 (
    .a (net22),
    .b (net20),
    .out (net43)
  );
  and_cell gate38 (
    .a (net43),
    .b (net24),
    .out (net44)
  );
  and_cell gate39 (
    .a (net44),
    .b (net34),
    .out (net45)
  );
  or_cell gate40 (
    .a (net27),
    .b (net30),
    .out (net46)
  );
  or_cell gate41 (
    .a (net35),
    .b (net39),
    .out (net47)
  );
  or_cell gate42 (
    .a (net42),
    .b (net45),
    .out (net48)
  );
  or_cell gate43 (
    .a (net47),
    .b (net48),
    .out (net49)
  );
  or_cell gate44 (
    .a (net46),
    .b (net49),
    .out (net50)
  );
  not_cell gate45 (
    .in (net21),
    .out (net31)
  );
  not_cell gate46 (
    .in (net19),
    .out (net23)
  );
  buffer_cell gate19 (
    .in (net7),
    .out (net38)
  );
  buffer_cell gate20 (
    .in (net51),
    .out (net24)
  );
  not_cell gate21 (
    .in (net51),
    .out (net28)
  );
  not_cell gate47 (
    .in (net7),
    .out (net34)
  );
  buffer_cell gate48 (
    .in (net8),
    .out (net52)
  );
  not_cell gate49 (
    .in (net8),
    .out (net26)
  );
  and_cell gate50 (
    .a (net23),
    .b (net24),
    .out (net53)
  );
  and_cell gate51 (
    .a (net53),
    .b (net52),
    .out (net54)
  );
  and_cell gate52 (
    .a (net20),
    .b (net28),
    .out (net55)
  );
  and_cell gate53 (
    .a (net55),
    .b (net52),
    .out (net56)
  );
  and_cell gate54 (
    .a (net31),
    .b (net23),
    .out (net57)
  );
  and_cell gate55 (
    .a (net57),
    .b (net38),
    .out (net58)
  );
  and_cell gate56 (
    .a (net58),
    .b (net52),
    .out (net59)
  );
  and_cell gate57 (
    .a (net31),
    .b (net24),
    .out (net60)
  );
  and_cell gate58 (
    .a (net60),
    .b (net34),
    .out (net61)
  );
  and_cell gate59 (
    .a (net61),
    .b (net52),
    .out (net62)
  );
  or_cell gate60 (
    .a (net54),
    .b (net56),
    .out (net63)
  );
  or_cell gate61 (
    .a (net59),
    .b (net62),
    .out (net64)
  );
  or_cell gate62 (
    .a (net63),
    .b (net64),
    .out (net65)
  );
  and_cell gate63 (
    .a (net22),
    .b (net20),
    .out (net66)
  );
  and_cell gate64 (
    .a (net66),
    .b (net24),
    .out (net67)
  );
  and_cell gate65 (
    .a (net67),
    .b (net38),
    .out (net68)
  );
  and_cell gate66 (
    .a (net31),
    .b (net23),
    .out (net69)
  );
  and_cell gate67 (
    .a (net69),
    .b (net28),
    .out (net70)
  );
  and_cell gate68 (
    .a (net70),
    .b (net38),
    .out (net71)
  );
  and_cell gate69 (
    .a (net71),
    .b (net26),
    .out (net72)
  );
  and_cell gate70 (
    .a (net31),
    .b (net20),
    .out (net73)
  );
  and_cell gate71 (
    .a (net73),
    .b (net24),
    .out (net74)
  );
  and_cell gate72 (
    .a (net74),
    .b (net34),
    .out (net75)
  );
  and_cell gate73 (
    .a (net75),
    .b (net26),
    .out (net76)
  );
  and_cell gate74 (
    .a (net22),
    .b (net23),
    .out (net77)
  );
  and_cell gate75 (
    .a (net77),
    .b (net28),
    .out (net78)
  );
  and_cell gate76 (
    .a (net78),
    .b (net34),
    .out (net79)
  );
  and_cell gate77 (
    .a (net79),
    .b (net26),
    .out (net80)
  );
  or_cell gate78 (
    .a (net68),
    .b (net72),
    .out (net81)
  );
  or_cell gate79 (
    .a (net76),
    .b (net80),
    .out (net82)
  );
  or_cell gate80 (
    .a (net81),
    .b (net82),
    .out (net83)
  );
  and_cell gate81 (
    .a (net22),
    .b (net23),
    .out (net84)
  );
  and_cell gate82 (
    .a (net84),
    .b (net28),
    .out (net85)
  );
  and_cell gate83 (
    .a (net85),
    .b (net34),
    .out (net86)
  );
  and_cell gate84 (
    .a (net86),
    .b (net52),
    .out (net87)
  );
  buffer_cell gate85 (
    .in (net2),
    .out (net88)
  );
  buffer_cell gate86 (
    .in (net3),
    .out (net89)
  );
  not_cell gate87 (
    .in (net3),
    .out (net90)
  );
  not_cell gate88 (
    .in (net2),
    .out (net91)
  );
  buffer_cell gate89 (
    .in (net83),
    .out (net92)
  );
  buffer_cell gate90 (
    .in (net87),
    .out (net93)
  );
  not_cell gate91 (
    .in (net87),
    .out (net94)
  );
  not_cell gate92 (
    .in (net83),
    .out (net95)
  );
  buffer_cell gate93 (
    .in (net65),
    .out (net96)
  );
  not_cell gate94 (
    .in (net65),
    .out (net97)
  );
  buffer_cell gate95 (
    .in (net4),
    .out (net98)
  );
  buffer_cell gate97 (
    .in (net50),
    .out (net99)
  );
  not_cell gate152 (
    .in (net100),
    .out (net101)
  );
  and_cell gate153 (
    .a (net101),
    .b (net102),
    .out (net103)
  );
  or_cell gate154 (
    .a (net103),
    .b (net104),
    .out (net105)
  );
  not_cell gate155 (
    .in (net102),
    .out (net106)
  );
  not_cell gate156 (
    .in (net107),
    .out (net108)
  );
  not_cell gate157 (
    .in (net109),
    .out (net110)
  );
  not_cell gate158 (
    .in (net111),
    .out (net112)
  );
  not_cell gate159 (
    .in (net113),
    .out (net114)
  );
  not_cell gate160 (
    .in (net115),
    .out (net116)
  );
  and_cell gate162 (
    .a (net100),
    .b (net106),
    .out (net104)
  );
  and_cell gate163 (
    .a (net108),
    .b (net109),
    .out (net117)
  );
  and_cell gate164 (
    .a (net107),
    .b (net110),
    .out (net118)
  );
  and_cell gate165 (
    .a (net112),
    .b (net113),
    .out (net119)
  );
  and_cell gate166 (
    .a (net111),
    .b (net114),
    .out (net120)
  );
  and_cell gate167 (
    .a (net116),
    .b (net121),
    .out (net122)
  );
  or_cell gate169 (
    .a (net117),
    .b (net118),
    .out (net123)
  );
  or_cell gate170 (
    .a (net119),
    .b (net120),
    .out (net124)
  );
  not_cell gate173 (
    .in (net124),
    .out (net125)
  );
  not_cell gate174 (
    .in (net123),
    .out (net126)
  );
  not_cell gate175 (
    .in (net105),
    .out (net127)
  );
  and_cell gate176 (
    .a (net127),
    .b (net117),
    .out (net128)
  );
  or_cell gate177 (
    .a (net103),
    .b (net128),
    .out (net129)
  );
  or_cell gate178 (
    .a (net129),
    .b (net130),
    .out (net131)
  );
  and_cell gate179 (
    .a (net132),
    .b (net119),
    .out (net130)
  );
  and_cell gate180 (
    .a (net127),
    .b (net126),
    .out (net132)
  );
  or_cell gate181 (
    .a (net131),
    .b (net133),
    .out (net134)
  );
  and_cell gate182 (
    .a (net135),
    .b (net122),
    .out (net133)
  );
  and_cell gate168 (
    .a (net132),
    .b (net125),
    .out (net135)
  );
  or_cell gate184 (
    .a (net136),
    .b (net99),
    .out (net137)
  );
  dff_cell flipflop15 (
    .d (net139),
    .clk (net13),
    .q (net10)
  );
  xor_cell gate161 (
    .a (net10),
    .b (net140),
    .out (net139)
  );
  dff_cell flipflop16 (
    .d (net141),
    .clk (net13),
    .q (net11)
  );
  xor_cell gate186 (
    .a (net11),
    .b (net142),
    .out (net141)
  );
  dff_cell flipflop17 (
    .d (net143),
    .clk (net13),
    .q (net12)
  );
  xor_cell gate187 (
    .a (net12),
    .b (net144),
    .out (net143)
  );
  and_cell gate188 (
    .a (net145),
    .b (net137),
    .out (net18)
  );
  and_cell gate190 (
    .a (net146),
    .b (net137),
    .out (net140)
  );
  and_cell gate191 (
    .a (net147),
    .b (net137),
    .out (net142)
  );
  and_cell gate192 (
    .a (net148),
    .b (net137),
    .out (net144)
  );
  and_cell gate193 (
    .a (net149),
    .b (net150),
    .out (net145)
  );
  and_cell gate194 (
    .a (net149),
    .b (net151),
    .out (net146)
  );
  and_cell gate195 (
    .a (net150),
    .b (net152),
    .out (net147)
  );
  and_cell gate196 (
    .a (net151),
    .b (net152),
    .out (net148)
  );
  not_cell gate197 (
    .in (net152),
    .out (net149)
  );
  not_cell gate198 (
    .in (net151),
    .out (net150)
  );
  or_cell gate7 (
    .a (net153),
    .b (net154),
    .out (net21)
  );
  or_cell gate8 (
    .a (net155),
    .b (net156),
    .out (net154)
  );
  or_cell gate9 (
    .a (net157),
    .b (net158),
    .out (net153)
  );
  and_cell gate10 (
    .a (net9),
    .b (net145),
    .out (net156)
  );
  and_cell gate11 (
    .a (net10),
    .b (net146),
    .out (net155)
  );
  and_cell gate12 (
    .a (net11),
    .b (net147),
    .out (net158)
  );
  and_cell gate13 (
    .a (net12),
    .b (net148),
    .out (net157)
  );
  or_cell gate14 (
    .a (net159),
    .b (net160),
    .out (net51)
  );
  or_cell gate15 (
    .a (net161),
    .b (net162),
    .out (net160)
  );
  or_cell gate16 (
    .a (net163),
    .b (net164),
    .out (net159)
  );
  and_cell gate17 (
    .a (net5),
    .b (net145),
    .out (net162)
  );
  and_cell gate171 (
    .a (net9),
    .b (net146),
    .out (net161)
  );
  and_cell gate172 (
    .a (net10),
    .b (net147),
    .out (net164)
  );
  and_cell gate183 (
    .a (net11),
    .b (net148),
    .out (net163)
  );
  or_cell gate189 (
    .a (net165),
    .b (net166),
    .out (net19)
  );
  or_cell gate199 (
    .a (net167),
    .b (net168),
    .out (net166)
  );
  or_cell gate200 (
    .a (net169),
    .b (net170),
    .out (net165)
  );
  and_cell gate201 (
    .a (net10),
    .b (net145),
    .out (net168)
  );
  and_cell gate202 (
    .a (net11),
    .b (net146),
    .out (net167)
  );
  and_cell gate203 (
    .a (net12),
    .b (net147),
    .out (net170)
  );
  and_cell gate204 (
    .a (net6),
    .b (net148),
    .out (net169)
  );
  dff_cell flipflop2 (
    .d (net171),
    .clk (net1),
    .q (net172),
    .notq (net173)
  );
  dff_cell flipflop3 (
    .d (net172),
    .clk (net1),
    .q (net174),
    .notq (net175)
  );
  dff_cell flipflop4 (
    .d (net174),
    .clk (net1),
    .q (net176),
    .notq (net177)
  );
  dff_cell flipflop5 (
    .d (net176),
    .clk (net1),
    .q (net178),
    .notq (net179)
  );
  or_cell gate205 (
    .a (net180),
    .b (net13),
    .out (net171)
  );
  and_cell gate206 (
    .a (net173),
    .b (net175),
    .out (net181)
  );
  and_cell gate207 (
    .a (net177),
    .b (net179),
    .out (net182)
  );
  and_cell gate208 (
    .a (net181),
    .b (net182),
    .out (net183)
  );
  dff_cell flipflop6 (
    .d (net178),
    .clk (net1),
    .q (net184),
    .notq (net185)
  );
  dff_cell flipflop7 (
    .d (net184),
    .clk (net1),
    .q (net186),
    .notq (net187)
  );
  and_cell gate209 (
    .a (net185),
    .b (net187),
    .out (net188)
  );
  and_cell gate210 (
    .a (net183),
    .b (net189),
    .out (net180)
  );
  dff_cell flipflop8 (
    .d (net190),
    .clk (net1),
    .q (net191),
    .notq (net192)
  );
  dff_cell flipflop9 (
    .d (net193),
    .clk (net1),
    .q (net194),
    .notq (net195)
  );
  and_cell gate211 (
    .a (net192),
    .b (net195),
    .out (net196)
  );
  or_cell gate212 (
    .a (net197),
    .b (net197),
    .out (net190)
  );
  or_cell gate213 (
    .a (net198),
    .b (net191),
    .out (net193)
  );
  dff_cell flipflop11 (
    .d (net199),
    .clk (net1),
    .q (net200),
    .notq (net201)
  );
  dff_cell flipflop12 (
    .d (net202),
    .clk (net1),
    .q (net203),
    .notq (net204)
  );
  and_cell gate214 (
    .a (net201),
    .b (net204),
    .out (net205)
  );
  or_cell gate215 (
    .a (net194),
    .b (net194),
    .out (net199)
  );
  or_cell gate216 (
    .a (net198),
    .b (net200),
    .out (net202)
  );
  dff_cell flipflop13 (
    .d (net206),
    .clk (net1),
    .q (net207),
    .notq (net208)
  );
  dff_cell flipflop14 (
    .d (net209),
    .clk (net1),
    .q (net210),
    .notq (net211)
  );
  and_cell gate217 (
    .a (net208),
    .b (net211),
    .out (net212)
  );
  or_cell gate218 (
    .a (net203),
    .b (net203),
    .out (net206)
  );
  or_cell gate219 (
    .a (net207),
    .b (net207),
    .out (net209)
  );
  dff_cell flipflop18 (
    .d (net213),
    .clk (net1),
    .q (net214),
    .notq (net215)
  );
  dff_cell flipflop19 (
    .d (net216),
    .clk (net1),
    .q (net217),
    .notq (net218)
  );
  and_cell gate220 (
    .a (net215),
    .b (net218),
    .out (net219)
  );
  or_cell gate221 (
    .a (net198),
    .b (net210),
    .out (net213)
  );
  or_cell gate222 (
    .a (net214),
    .b (net214),
    .out (net216)
  );
  dff_cell flipflop20 (
    .d (net220),
    .clk (net1),
    .q (net221),
    .notq (net222)
  );
  dff_cell flipflop21 (
    .d (net223),
    .clk (net1),
    .q (net224),
    .notq (net225)
  );
  and_cell gate223 (
    .a (net222),
    .b (net225),
    .out (net226)
  );
  or_cell gate224 (
    .a (net217),
    .b (net217),
    .out (net220)
  );
  or_cell gate225 (
    .a (net198),
    .b (net221),
    .out (net223)
  );
  dff_cell flipflop22 (
    .d (net227),
    .clk (net1),
    .q (net228),
    .notq (net229)
  );
  dff_cell flipflop23 (
    .d (net230),
    .clk (net1),
    .q (net231),
    .notq (net232)
  );
  and_cell gate226 (
    .a (net229),
    .b (net232),
    .out (net233)
  );
  or_cell gate227 (
    .a (net224),
    .b (net224),
    .out (net227)
  );
  or_cell gate228 (
    .a (net228),
    .b (net228),
    .out (net230)
  );
  dff_cell flipflop24 (
    .d (net234),
    .clk (net1),
    .q (net235),
    .notq (net236)
  );
  dff_cell flipflop25 (
    .d (net237),
    .clk (net1),
    .q (net238),
    .notq (net239)
  );
  and_cell gate229 (
    .a (net236),
    .b (net239),
    .out (net240)
  );
  or_cell gate230 (
    .a (net231),
    .b (net231),
    .out (net234)
  );
  or_cell gate231 (
    .a (net235),
    .b (net235),
    .out (net237)
  );
  dff_cell flipflop26 (
    .d (net241),
    .clk (net1),
    .q (net242),
    .notq (net243)
  );
  dff_cell flipflop27 (
    .d (net244),
    .clk (net1),
    .q (net245),
    .notq (net246)
  );
  and_cell gate232 (
    .a (net243),
    .b (net246),
    .out (net247)
  );
  or_cell gate233 (
    .a (net238),
    .b (net238),
    .out (net241)
  );
  or_cell gate234 (
    .a (net198),
    .b (net242),
    .out (net244)
  );
  dff_cell flipflop28 (
    .d (net248),
    .clk (net1),
    .q (net249),
    .notq (net250)
  );
  dff_cell flipflop29 (
    .d (net251),
    .clk (net1),
    .q (net252),
    .notq (net253)
  );
  and_cell gate235 (
    .a (net250),
    .b (net253),
    .out (net254)
  );
  or_cell gate236 (
    .a (net245),
    .b (net245),
    .out (net248)
  );
  or_cell gate237 (
    .a (net198),
    .b (net249),
    .out (net251)
  );
  dff_cell flipflop30 (
    .d (net255),
    .clk (net1),
    .q (net256),
    .notq (net257)
  );
  dff_cell flipflop31 (
    .d (net258),
    .clk (net1),
    .q (net259),
    .notq (net260)
  );
  and_cell gate238 (
    .a (net257),
    .b (net260),
    .out (net261)
  );
  or_cell gate239 (
    .a (net252),
    .b (net252),
    .out (net255)
  );
  or_cell gate240 (
    .a (net256),
    .b (net256),
    .out (net258)
  );
  dff_cell flipflop32 (
    .d (net262),
    .clk (net1),
    .q (net263),
    .notq (net264)
  );
  dff_cell flipflop33 (
    .d (net265),
    .clk (net1),
    .q (net266),
    .notq (net267)
  );
  and_cell gate241 (
    .a (net264),
    .b (net267),
    .out (net268)
  );
  or_cell gate242 (
    .a (net198),
    .b (net259),
    .out (net262)
  );
  or_cell gate243 (
    .a (net198),
    .b (net263),
    .out (net265)
  );
  dff_cell flipflop34 (
    .d (net269),
    .clk (net1),
    .q (net270),
    .notq (net271)
  );
  dff_cell flipflop35 (
    .d (net272),
    .clk (net1),
    .q (net273),
    .notq (net274)
  );
  and_cell gate244 (
    .a (net271),
    .b (net274),
    .out (net275)
  );
  or_cell gate245 (
    .a (net198),
    .b (net266),
    .out (net269)
  );
  or_cell gate246 (
    .a (net270),
    .b (net270),
    .out (net272)
  );
  dff_cell flipflop36 (
    .d (net276),
    .clk (net1),
    .q (net277),
    .notq (net278)
  );
  dff_cell flipflop37 (
    .d (net279),
    .clk (net1),
    .q (net280),
    .notq (net281)
  );
  and_cell gate247 (
    .a (net278),
    .b (net281),
    .out (net282)
  );
  or_cell gate248 (
    .a (net273),
    .b (net273),
    .out (net276)
  );
  or_cell gate249 (
    .a (net198),
    .b (net277),
    .out (net279)
  );
  dff_cell flipflop38 (
    .d (net283),
    .clk (net1),
    .q (net115),
    .notq (net284)
  );
  dff_cell flipflop39 (
    .d (net285),
    .clk (net1),
    .q (net111),
    .notq (net286)
  );
  and_cell gate250 (
    .a (net284),
    .b (net286),
    .out (net287)
  );
  or_cell gate251 (
    .a (net280),
    .b (net280),
    .out (net283)
  );
  or_cell gate252 (
    .a (net115),
    .b (net115),
    .out (net285)
  );
  dff_cell flipflop40 (
    .d (net288),
    .clk (net1),
    .q (net107),
    .notq (net289)
  );
  dff_cell flipflop41 (
    .d (net290),
    .clk (net1),
    .q (net100),
    .notq (net291)
  );
  and_cell gate253 (
    .a (net289),
    .b (net291),
    .out (net292)
  );
  or_cell gate254 (
    .a (net111),
    .b (net111),
    .out (net288)
  );
  or_cell gate255 (
    .a (net198),
    .b (net107),
    .out (net290)
  );
  dff_cell flipflop42 (
    .d (net293),
    .clk (net1),
    .q (net151),
    .notq (net294)
  );
  dff_cell flipflop43 (
    .d (net295),
    .clk (net1),
    .q (net152),
    .notq (net296)
  );
  and_cell gate256 (
    .a (net294),
    .b (net296),
    .out (net297)
  );
  or_cell gate257 (
    .a (net100),
    .b (net100),
    .out (net293)
  );
  or_cell gate258 (
    .a (net151),
    .b (net151),
    .out (net295)
  );
  and_cell gate259 (
    .a (net254),
    .b (net298),
    .out (net299)
  );
  and_cell gate260 (
    .a (net300),
    .b (net299),
    .out (net198)
  );
  and_cell gate261 (
    .a (net196),
    .b (net301),
    .out (net300)
  );
  and_cell gate262 (
    .a (net261),
    .b (net302),
    .out (net298)
  );
  and_cell gate263 (
    .a (net268),
    .b (net303),
    .out (net302)
  );
  and_cell gate264 (
    .a (net275),
    .b (net304),
    .out (net303)
  );
  and_cell gate265 (
    .a (net282),
    .b (net305),
    .out (net304)
  );
  and_cell gate266 (
    .a (net287),
    .b (net306),
    .out (net305)
  );
  and_cell gate267 (
    .a (net292),
    .b (net297),
    .out (net306)
  );
  and_cell gate268 (
    .a (net205),
    .b (net307),
    .out (net301)
  );
  and_cell gate269 (
    .a (net212),
    .b (net308),
    .out (net307)
  );
  and_cell gate270 (
    .a (net219),
    .b (net309),
    .out (net308)
  );
  and_cell gate271 (
    .a (net226),
    .b (net310),
    .out (net309)
  );
  and_cell gate272 (
    .a (net233),
    .b (net311),
    .out (net310)
  );
  and_cell gate273 (
    .a (net240),
    .b (net247),
    .out (net311)
  );
  xor_cell xor1 (
    .a (net312),
    .b (net194),
    .out (net313)
  );
  xor_cell xor2 (
    .a (net152),
    .b (net266),
    .out (net312)
  );
  xor_cell xor3 (
    .a (net313),
    .b (net191),
    .out (net197)
  );
  not_cell gate96 (
    .in (net4),
    .out (net314)
  );
  and_cell gate100 (
    .a (net88),
    .b (net97),
    .out (net315)
  );
  and_cell gate101 (
    .a (net314),
    .b (net88),
    .out (net316)
  );
  and_cell gate102 (
    .a (net89),
    .b (net92),
    .out (net317)
  );
  and_cell gate103 (
    .a (net314),
    .b (net89),
    .out (net318)
  );
  and_cell gate104 (
    .a (net318),
    .b (net97),
    .out (net319)
  );
  and_cell gate105 (
    .a (net98),
    .b (net90),
    .out (net320)
  );
  and_cell gate106 (
    .a (net320),
    .b (net93),
    .out (net321)
  );
  and_cell gate107 (
    .a (net98),
    .b (net91),
    .out (net322)
  );
  and_cell gate108 (
    .a (net322),
    .b (net96),
    .out (net323)
  );
  or_cell gate109 (
    .a (net315),
    .b (net316),
    .out (net324)
  );
  or_cell gate110 (
    .a (net324),
    .b (net325),
    .out (net326)
  );
  or_cell gate111 (
    .a (net317),
    .b (net319),
    .out (net325)
  );
  or_cell gate112 (
    .a (net321),
    .b (net323),
    .out (net327)
  );
  or_cell gate113 (
    .a (net326),
    .b (net327),
    .out (net328)
  );
  and_cell gate114 (
    .a (net98),
    .b (net91),
    .out (net329)
  );
  and_cell gate115 (
    .a (net329),
    .b (net94),
    .out (net330)
  );
  and_cell gate116 (
    .a (net89),
    .b (net91),
    .out (net331)
  );
  and_cell gate117 (
    .a (net331),
    .b (net94),
    .out (net332)
  );
  or_cell gate118 (
    .a (net330),
    .b (net332),
    .out (net333)
  );
  and_cell gate119 (
    .a (net98),
    .b (net89),
    .out (net334)
  );
  and_cell gate120 (
    .a (net334),
    .b (net91),
    .out (net335)
  );
  and_cell gate121 (
    .a (net314),
    .b (net89),
    .out (net336)
  );
  and_cell gate122 (
    .a (net336),
    .b (net88),
    .out (net337)
  );
  or_cell gate123 (
    .a (net335),
    .b (net337),
    .out (net338)
  );
  and_cell gate124 (
    .a (net98),
    .b (net90),
    .out (net339)
  );
  and_cell gate125 (
    .a (net339),
    .b (net92),
    .out (net340)
  );
  and_cell gate126 (
    .a (net314),
    .b (net88),
    .out (net341)
  );
  and_cell gate127 (
    .a (net341),
    .b (net96),
    .out (net342)
  );
  or_cell gate128 (
    .a (net340),
    .b (net342),
    .out (net343)
  );
  or_cell gate129 (
    .a (net333),
    .b (net344),
    .out (net345)
  );
  or_cell gate130 (
    .a (net338),
    .b (net343),
    .out (net344)
  );
  and_cell gate131 (
    .a (net89),
    .b (net91),
    .out (net346)
  );
  and_cell gate132 (
    .a (net346),
    .b (net95),
    .out (net347)
  );
  and_cell gate133 (
    .a (net98),
    .b (net89),
    .out (net348)
  );
  and_cell gate134 (
    .a (net348),
    .b (net93),
    .out (net349)
  );
  or_cell gate135 (
    .a (net347),
    .b (net349),
    .out (net350)
  );
  and_cell gate136 (
    .a (net351),
    .b (net88),
    .out (net352)
  );
  and_cell gate137 (
    .a (net352),
    .b (net95),
    .out (net353)
  );
  and_cell gate138 (
    .a (net354),
    .b (net91),
    .out (net355)
  );
  and_cell gate139 (
    .a (net355),
    .b (net92),
    .out (net356)
  );
  or_cell gate140 (
    .a (net353),
    .b (net356),
    .out (net357)
  );
  and_cell gate141 (
    .a (net98),
    .b (net90),
    .out (net351)
  );
  and_cell gate142 (
    .a (net98),
    .b (net90),
    .out (net354)
  );
  and_cell gate143 (
    .a (net358),
    .b (net88),
    .out (net359)
  );
  and_cell gate144 (
    .a (net359),
    .b (net92),
    .out (net360)
  );
  and_cell gate145 (
    .a (net314),
    .b (net90),
    .out (net358)
  );
  or_cell gate146 (
    .a (net361),
    .b (net357),
    .out (net362)
  );
  or_cell gate147 (
    .a (net350),
    .b (net360),
    .out (net361)
  );
  and_cell gate148 (
    .a (net98),
    .b (net90),
    .out (net363)
  );
  and_cell gate149 (
    .a (net363),
    .b (net95),
    .out (net364)
  );
  and_cell gate150 (
    .a (net98),
    .b (net90),
    .out (net365)
  );
  and_cell gate151 (
    .a (net365),
    .b (net91),
    .out (net366)
  );
  or_cell gate274 (
    .a (net364),
    .b (net366),
    .out (net367)
  );
  and_cell gate275 (
    .a (net98),
    .b (net93),
    .out (net368)
  );
  and_cell gate276 (
    .a (net369),
    .b (net91),
    .out (net370)
  );
  and_cell gate277 (
    .a (net370),
    .b (net95),
    .out (net371)
  );
  and_cell gate278 (
    .a (net314),
    .b (net89),
    .out (net369)
  );
  or_cell gate279 (
    .a (net368),
    .b (net367),
    .out (net372)
  );
  or_cell gate280 (
    .a (net372),
    .b (net371),
    .out (net373)
  );
  and_cell gate98 (
    .a (net98),
    .b (net91),
    .out (net374)
  );
  and_cell gate99 (
    .a (net374),
    .b (net95),
    .out (net375)
  );
  and_cell gate281 (
    .a (net98),
    .b (net90),
    .out (net376)
  );
  and_cell gate282 (
    .a (net376),
    .b (net91),
    .out (net377)
  );
  or_cell gate283 (
    .a (net375),
    .b (net377),
    .out (net378)
  );
  and_cell gate284 (
    .a (net98),
    .b (net88),
    .out (net379)
  );
  and_cell gate285 (
    .a (net379),
    .b (net92),
    .out (net380)
  );
  and_cell gate286 (
    .a (net89),
    .b (net91),
    .out (net381)
  );
  and_cell gate287 (
    .a (net381),
    .b (net96),
    .out (net382)
  );
  or_cell gate288 (
    .a (net380),
    .b (net382),
    .out (net383)
  );
  or_cell gate289 (
    .a (net378),
    .b (net383),
    .out (net121)
  );
  and_cell gate290 (
    .a (net89),
    .b (net88),
    .out (net384)
  );
  and_cell gate291 (
    .a (net384),
    .b (net93),
    .out (net385)
  );
  and_cell gate292 (
    .a (net90),
    .b (net88),
    .out (net386)
  );
  and_cell gate293 (
    .a (net386),
    .b (net96),
    .out (net387)
  );
  or_cell gate294 (
    .a (net385),
    .b (net387),
    .out (net388)
  );
  and_cell gate295 (
    .a (net389),
    .b (net88),
    .out (net390)
  );
  and_cell gate296 (
    .a (net390),
    .b (net94),
    .out (net391)
  );
  and_cell gate297 (
    .a (net392),
    .b (net91),
    .out (net393)
  );
  and_cell gate298 (
    .a (net393),
    .b (net93),
    .out (net394)
  );
  or_cell gate299 (
    .a (net391),
    .b (net394),
    .out (net395)
  );
  and_cell gate300 (
    .a (net98),
    .b (net90),
    .out (net389)
  );
  and_cell gate301 (
    .a (net98),
    .b (net90),
    .out (net392)
  );
  and_cell gate302 (
    .a (net396),
    .b (net91),
    .out (net397)
  );
  and_cell gate303 (
    .a (net397),
    .b (net92),
    .out (net398)
  );
  and_cell gate304 (
    .a (net399),
    .b (net91),
    .out (net400)
  );
  and_cell gate305 (
    .a (net400),
    .b (net96),
    .out (net401)
  );
  or_cell gate306 (
    .a (net398),
    .b (net401),
    .out (net402)
  );
  and_cell gate307 (
    .a (net314),
    .b (net89),
    .out (net396)
  );
  and_cell gate308 (
    .a (net98),
    .b (net89),
    .out (net399)
  );
  or_cell gate309 (
    .a (net395),
    .b (net402),
    .out (net403)
  );
  or_cell gate310 (
    .a (net388),
    .b (net403),
    .out (net113)
  );
  and_cell gate311 (
    .a (net98),
    .b (net89),
    .out (net404)
  );
  and_cell gate312 (
    .a (net404),
    .b (net93),
    .out (net405)
  );
  and_cell gate313 (
    .a (net98),
    .b (net88),
    .out (net406)
  );
  and_cell gate314 (
    .a (net406),
    .b (net93),
    .out (net407)
  );
  or_cell gate315 (
    .a (net405),
    .b (net407),
    .out (net408)
  );
  and_cell gate316 (
    .a (net98),
    .b (net90),
    .out (net409)
  );
  and_cell gate317 (
    .a (net409),
    .b (net92),
    .out (net410)
  );
  and_cell gate318 (
    .a (net411),
    .b (net88),
    .out (net412)
  );
  and_cell gate319 (
    .a (net412),
    .b (net92),
    .out (net413)
  );
  and_cell gate320 (
    .a (net414),
    .b (net91),
    .out (net415)
  );
  and_cell gate321 (
    .a (net415),
    .b (net96),
    .out (net416)
  );
  or_cell gate322 (
    .a (net413),
    .b (net416),
    .out (net417)
  );
  and_cell gate323 (
    .a (net314),
    .b (net89),
    .out (net411)
  );
  and_cell gate324 (
    .a (net314),
    .b (net89),
    .out (net414)
  );
  and_cell gate325 (
    .a (net418),
    .b (net88),
    .out (net419)
  );
  and_cell gate326 (
    .a (net419),
    .b (net95),
    .out (net420)
  );
  and_cell gate327 (
    .a (net98),
    .b (net89),
    .out (net418)
  );
  or_cell gate328 (
    .a (net410),
    .b (net420),
    .out (net421)
  );
  or_cell gate329 (
    .a (net408),
    .b (net421),
    .out (net422)
  );
  or_cell gate330 (
    .a (net422),
    .b (net417),
    .out (net109)
  );
  and_cell gate331 (
    .a (net98),
    .b (net89),
    .out (net423)
  );
  and_cell gate332 (
    .a (net423),
    .b (net94),
    .out (net424)
  );
  and_cell gate333 (
    .a (net89),
    .b (net88),
    .out (net425)
  );
  and_cell gate334 (
    .a (net425),
    .b (net96),
    .out (net426)
  );
  or_cell gate335 (
    .a (net424),
    .b (net426),
    .out (net427)
  );
  and_cell gate336 (
    .a (net98),
    .b (net96),
    .out (net428)
  );
  or_cell gate337 (
    .a (net428),
    .b (net427),
    .out (net102)
  );
  and_cell gate1 (
    .a (net115),
    .b (net429),
    .out (net430)
  );
  not_cell gate2 (
    .in (net121),
    .out (net429)
  );
  or_cell gate3 (
    .a (net122),
    .b (net430),
    .out (net431)
  );
  not_cell gate4 (
    .in (net431),
    .out (net432)
  );
  and_cell gate5 (
    .a (net135),
    .b (net432),
    .out (net433)
  );
  or_cell gate6 (
    .a (net134),
    .b (net433),
    .out (net434)
  );
  not_cell gate185 (
    .in (net280),
    .out (net435)
  );
  and_cell gate338 (
    .a (net435),
    .b (net373),
    .out (net436)
  );
  or_cell gate339 (
    .a (net436),
    .b (net437),
    .out (net438)
  );
  not_cell gate340 (
    .in (net373),
    .out (net439)
  );
  not_cell gate341 (
    .in (net277),
    .out (net440)
  );
  not_cell gate342 (
    .in (net362),
    .out (net441)
  );
  not_cell gate343 (
    .in (net273),
    .out (net442)
  );
  not_cell gate344 (
    .in (net345),
    .out (net443)
  );
  not_cell gate345 (
    .in (net270),
    .out (net444)
  );
  and_cell gate346 (
    .a (net280),
    .b (net439),
    .out (net437)
  );
  and_cell gate347 (
    .a (net440),
    .b (net362),
    .out (net445)
  );
  and_cell gate348 (
    .a (net277),
    .b (net441),
    .out (net446)
  );
  and_cell gate349 (
    .a (net442),
    .b (net345),
    .out (net447)
  );
  and_cell gate350 (
    .a (net273),
    .b (net443),
    .out (net448)
  );
  and_cell gate351 (
    .a (net444),
    .b (net449),
    .out (net450)
  );
  or_cell gate352 (
    .a (net445),
    .b (net446),
    .out (net451)
  );
  or_cell gate353 (
    .a (net447),
    .b (net448),
    .out (net452)
  );
  not_cell gate354 (
    .in (net452),
    .out (net453)
  );
  not_cell gate355 (
    .in (net451),
    .out (net454)
  );
  not_cell gate356 (
    .in (net438),
    .out (net455)
  );
  and_cell gate357 (
    .a (net455),
    .b (net445),
    .out (net456)
  );
  or_cell gate358 (
    .a (net436),
    .b (net456),
    .out (net457)
  );
  or_cell gate359 (
    .a (net457),
    .b (net458),
    .out (net459)
  );
  and_cell gate360 (
    .a (net460),
    .b (net447),
    .out (net458)
  );
  and_cell gate361 (
    .a (net455),
    .b (net454),
    .out (net460)
  );
  or_cell gate362 (
    .a (net459),
    .b (net461),
    .out (net462)
  );
  and_cell gate363 (
    .a (net463),
    .b (net450),
    .out (net461)
  );
  and_cell gate364 (
    .a (net460),
    .b (net453),
    .out (net463)
  );
  and_cell gate371 (
    .a (net434),
    .b (net462),
    .out (net136)
  );
  buffer_cell gate365 (
    .in (net328),
    .out (net449)
  );
  dff_cell flipflop1 (
    .d (net186),
    .clk (net1),
    .q (net464),
    .notq (net465)
  );
  dff_cell flipflop44 (
    .d (net464),
    .clk (net1),
    .q (net466),
    .notq (net467)
  );
  and_cell gate366 (
    .a (net465),
    .b (net467),
    .out (net468)
  );
  dff_cell flipflop45 (
    .d (net466),
    .clk (net1),
    .q (net469),
    .notq (net470)
  );
  dff_cell flipflop46 (
    .d (net469),
    .clk (net1),
    .q (net13),
    .notq (net471)
  );
  and_cell gate367 (
    .a (net470),
    .b (net471),
    .out (net472)
  );
  and_cell gate368 (
    .a (net188),
    .b (net473),
    .out (net189)
  );
  and_cell gate369 (
    .a (net468),
    .b (net472),
    .out (net473)
  );
endmodule
