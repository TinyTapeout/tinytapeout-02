* NGSPICE file created from user_project_wrapper.ext - technology: sky130B

* Black-box entry subcircuit for user_module_349011320806310484 abstract view
.subckt user_module_349011320806310484 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341589685194195540 abstract view
.subckt user_module_341589685194195540 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for scanchain abstract view
.subckt scanchain clk_in clk_out data_in data_out latch_enable_in latch_enable_out
+ module_data_in[0] module_data_in[1] module_data_in[2] module_data_in[3] module_data_in[4]
+ module_data_in[5] module_data_in[6] module_data_in[7] module_data_out[0] module_data_out[1]
+ module_data_out[2] module_data_out[3] module_data_out[4] module_data_out[5] module_data_out[6]
+ module_data_out[7] scan_select_in scan_select_out vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348255968419643987 abstract view
.subckt user_module_348255968419643987 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341535056611770964 abstract view
.subckt user_module_341535056611770964 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for xor_shift32_quantamhd abstract view
.subckt xor_shift32_quantamhd io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tomkeddie_top_tto abstract view
.subckt tomkeddie_top_tto io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for tholin_avalonsemi_5401 abstract view
.subckt tholin_avalonsemi_5401 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for AidanMedcalf_pid_controller abstract view
.subckt AidanMedcalf_pid_controller io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348381622440034899 abstract view
.subckt user_module_348381622440034899 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for ericsmi_speed_test abstract view
.subckt ericsmi_speed_test io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for aramsey118_freq_counter abstract view
.subckt aramsey118_freq_counter io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341423712597181012 abstract view
.subckt user_module_341423712597181012 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348121131386929746 abstract view
.subckt user_module_348121131386929746 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341620484740219475 abstract view
.subckt user_module_341620484740219475 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347619669052490324 abstract view
.subckt user_module_347619669052490324 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for jar_illegal_logic abstract view
.subckt jar_illegal_logic io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for meriac_tt02_play_tune abstract view
.subckt meriac_tt02_play_tune io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341178154799333971 abstract view
.subckt user_module_341178154799333971 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt2_tholin_namebadge abstract view
.subckt tt2_tholin_namebadge io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341490465660469844 abstract view
.subckt user_module_341490465660469844 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341608574336631379 abstract view
.subckt user_module_341608574336631379 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for krasin_3_bit_8_channel_pwm_driver abstract view
.subckt krasin_3_bit_8_channel_pwm_driver io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for thunderbird_taillight_ctrl abstract view
.subckt thunderbird_taillight_ctrl io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for mbikovitsky_top abstract view
.subckt mbikovitsky_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347592305412145748 abstract view
.subckt user_module_347592305412145748 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for moyes0_top_module abstract view
.subckt moyes0_top_module io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for cpldcpu_MCPU5plus abstract view
.subckt cpldcpu_MCPU5plus io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_342981109408072274 abstract view
.subckt user_module_342981109408072274 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt2_tholin_diceroll abstract view
.subckt tt2_tholin_diceroll io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_nickoe abstract view
.subckt user_module_nickoe io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341541108650607187 abstract view
.subckt user_module_341541108650607187 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_349546262775726676 abstract view
.subckt user_module_349546262775726676 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for github_com_proppy_tt02_xls_popcount abstract view
.subckt github_com_proppy_tt02_xls_popcount io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341614374571475540 abstract view
.subckt user_module_341614374571475540 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for krasin_tt02_verilog_spi_7_channel_pwm_driver abstract view
.subckt krasin_tt02_verilog_spi_7_channel_pwm_driver io_in[0] io_in[1] io_in[2] io_in[3]
+ io_in[4] io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for udxs_sqrt_top abstract view
.subckt udxs_sqrt_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for moonbase_cpu_8bit abstract view
.subckt moonbase_cpu_8bit io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for loxodes_sequencer abstract view
.subckt loxodes_sequencer io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347594509754827347 abstract view
.subckt user_module_347594509754827347 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for yupferris_bitslam abstract view
.subckt yupferris_bitslam io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for phasenoisepon_seven_segment_seconds abstract view
.subckt phasenoisepon_seven_segment_seconds io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348961139276644947 abstract view
.subckt user_module_348961139276644947 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for migcorre_pwm abstract view
.subckt migcorre_pwm io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_346553315158393428 abstract view
.subckt user_module_346553315158393428 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for jar_sram_top abstract view
.subckt jar_sram_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for yubex_egg_timer abstract view
.subckt yubex_egg_timer io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for flygoat_tt02_play_tune abstract view
.subckt flygoat_tt02_play_tune io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for s4ga abstract view
.subckt s4ga io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for rc5_top abstract view
.subckt rc5_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_349228308755382868 abstract view
.subckt user_module_349228308755382868 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for mm21_LEDMatrixTop abstract view
.subckt mm21_LEDMatrixTop io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for cchan_fp8_multiplier abstract view
.subckt cchan_fp8_multiplier io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341516949939814994 abstract view
.subckt user_module_341516949939814994 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tholin_avalonsemi_tbb1143 abstract view
.subckt tholin_avalonsemi_tbb1143 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for wren6991_whisk_tt2_io_wrapper abstract view
.subckt wren6991_whisk_tt2_io_wrapper io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for azdle_binary_clock abstract view
.subckt azdle_binary_clock io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_346916357828248146 abstract view
.subckt user_module_346916357828248146 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tomkeddie_top_tto_a abstract view
.subckt tomkeddie_top_tto_a io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tiny_fft abstract view
.subckt tiny_fft io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for rolfmobile99_alu_fsm_top abstract view
.subckt rolfmobile99_alu_fsm_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348260124451668562 abstract view
.subckt user_module_348260124451668562 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for zoechip abstract view
.subckt zoechip io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for xyz_peppergray_Potato1_top abstract view
.subckt xyz_peppergray_Potato1_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for hex_sr abstract view
.subckt hex_sr io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341277789473735250 abstract view
.subckt user_module_341277789473735250 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347894637149553236 abstract view
.subckt user_module_347894637149553236 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for alu_top abstract view
.subckt alu_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for moonbase_cpu_4bit abstract view
.subckt moonbase_cpu_4bit io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341164910646919762 abstract view
.subckt user_module_341164910646919762 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for fraserbc_simon abstract view
.subckt fraserbc_simon io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for davidsiaw_stackcalc abstract view
.subckt davidsiaw_stackcalc io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt2_tholin_multiplier abstract view
.subckt tt2_tholin_multiplier io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341571228858843732 abstract view
.subckt user_module_341571228858843732 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for xor_shift32_evango abstract view
.subckt xor_shift32_evango io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for github_com_proppy_tt02_xls_counter abstract view
.subckt github_com_proppy_tt02_xls_counter io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for tt2_tholin_multiplexed_counter abstract view
.subckt tt2_tholin_multiplexed_counter io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for asic_multiplier_wrapper abstract view
.subckt asic_multiplier_wrapper io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_349405063877231188 abstract view
.subckt user_module_349405063877231188 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for pwm_gen abstract view
.subckt pwm_gen io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348195845106041428 abstract view
.subckt user_module_348195845106041428 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for aidan_McCoy abstract view
.subckt aidan_McCoy io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_341609034095264340 abstract view
.subckt user_module_341609034095264340 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for scan_controller abstract view
.subckt scan_controller active_select[0] active_select[1] active_select[2] active_select[3]
+ active_select[4] active_select[5] active_select[6] active_select[7] active_select[8]
+ clk driver_sel[0] driver_sel[1] inputs[0] inputs[1] inputs[2] inputs[3] inputs[4]
+ inputs[5] inputs[6] inputs[7] la_scan_clk_in la_scan_data_in la_scan_data_out la_scan_latch_en
+ la_scan_select oeb[0] oeb[10] oeb[11] oeb[12] oeb[13] oeb[14] oeb[15] oeb[16] oeb[17]
+ oeb[18] oeb[19] oeb[1] oeb[20] oeb[21] oeb[22] oeb[23] oeb[24] oeb[25] oeb[26] oeb[27]
+ oeb[28] oeb[29] oeb[2] oeb[30] oeb[31] oeb[32] oeb[33] oeb[34] oeb[35] oeb[36] oeb[37]
+ oeb[3] oeb[4] oeb[5] oeb[6] oeb[7] oeb[8] oeb[9] outputs[0] outputs[1] outputs[2]
+ outputs[3] outputs[4] outputs[5] outputs[6] outputs[7] ready reset scan_clk_in scan_clk_out
+ scan_data_in scan_data_out scan_latch_en scan_select set_clk_div slow_clk vccd1
+ vssd1
.ends

* Black-box entry subcircuit for user_module_347688030570545747 abstract view
.subckt user_module_347688030570545747 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for chase_the_beat abstract view
.subckt chase_the_beat io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_349047610915422802 abstract view
.subckt user_module_349047610915422802 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for navray_top abstract view
.subckt navray_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for gatecat_fpga_top abstract view
.subckt gatecat_fpga_top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for thezoq2_yafpga abstract view
.subckt thezoq2_yafpga io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_340318610245288530 abstract view
.subckt user_module_340318610245288530 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for chrisruk_matrix abstract view
.subckt chrisruk_matrix io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5] io_in[6]
+ io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348540666182107731 abstract view
.subckt user_module_348540666182107731 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347787021138264660 abstract view
.subckt user_module_347787021138264660 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for cpldcpu_TrainLED2top abstract view
.subckt cpldcpu_TrainLED2top io_in[0] io_in[1] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_347690870424732244 abstract view
.subckt user_module_347690870424732244 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348787952842703444 abstract view
.subckt user_module_348787952842703444 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

* Black-box entry subcircuit for user_module_348242239268323922 abstract view
.subckt user_module_348242239268323922 io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] vccd1 vssd1
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xuser_module_349011320806310484_071 scanchain_071/module_data_in[0] scanchain_071/module_data_in[1]
+ scanchain_071/module_data_in[2] scanchain_071/module_data_in[3] scanchain_071/module_data_in[4]
+ scanchain_071/module_data_in[5] scanchain_071/module_data_in[6] scanchain_071/module_data_in[7]
+ scanchain_071/module_data_out[0] scanchain_071/module_data_out[1] scanchain_071/module_data_out[2]
+ scanchain_071/module_data_out[3] scanchain_071/module_data_out[4] scanchain_071/module_data_out[5]
+ scanchain_071/module_data_out[6] scanchain_071/module_data_out[7] vccd1 vssd1 user_module_349011320806310484
Xuser_module_341589685194195540_090 scanchain_090/module_data_in[0] scanchain_090/module_data_in[1]
+ scanchain_090/module_data_in[2] scanchain_090/module_data_in[3] scanchain_090/module_data_in[4]
+ scanchain_090/module_data_in[5] scanchain_090/module_data_in[6] scanchain_090/module_data_in[7]
+ scanchain_090/module_data_out[0] scanchain_090/module_data_out[1] scanchain_090/module_data_out[2]
+ scanchain_090/module_data_out[3] scanchain_090/module_data_out[4] scanchain_090/module_data_out[5]
+ scanchain_090/module_data_out[6] scanchain_090/module_data_out[7] vccd1 vssd1 user_module_341589685194195540
Xscanchain_150 scanchain_150/clk_in scanchain_151/clk_in scanchain_150/data_in scanchain_151/data_in
+ scanchain_150/latch_enable_in scanchain_151/latch_enable_in scanchain_150/module_data_in[0]
+ scanchain_150/module_data_in[1] scanchain_150/module_data_in[2] scanchain_150/module_data_in[3]
+ scanchain_150/module_data_in[4] scanchain_150/module_data_in[5] scanchain_150/module_data_in[6]
+ scanchain_150/module_data_in[7] scanchain_150/module_data_out[0] scanchain_150/module_data_out[1]
+ scanchain_150/module_data_out[2] scanchain_150/module_data_out[3] scanchain_150/module_data_out[4]
+ scanchain_150/module_data_out[5] scanchain_150/module_data_out[6] scanchain_150/module_data_out[7]
+ scanchain_150/scan_select_in scanchain_151/scan_select_in vccd1 vssd1 scanchain
Xscanchain_161 scanchain_161/clk_in scanchain_162/clk_in scanchain_161/data_in scanchain_162/data_in
+ scanchain_161/latch_enable_in scanchain_162/latch_enable_in scanchain_161/module_data_in[0]
+ scanchain_161/module_data_in[1] scanchain_161/module_data_in[2] scanchain_161/module_data_in[3]
+ scanchain_161/module_data_in[4] scanchain_161/module_data_in[5] scanchain_161/module_data_in[6]
+ scanchain_161/module_data_in[7] scanchain_161/module_data_out[0] scanchain_161/module_data_out[1]
+ scanchain_161/module_data_out[2] scanchain_161/module_data_out[3] scanchain_161/module_data_out[4]
+ scanchain_161/module_data_out[5] scanchain_161/module_data_out[6] scanchain_161/module_data_out[7]
+ scanchain_161/scan_select_in scanchain_162/scan_select_in vccd1 vssd1 scanchain
Xscanchain_194 scanchain_194/clk_in scanchain_195/clk_in scanchain_194/data_in scanchain_195/data_in
+ scanchain_194/latch_enable_in scanchain_195/latch_enable_in scanchain_194/module_data_in[0]
+ scanchain_194/module_data_in[1] scanchain_194/module_data_in[2] scanchain_194/module_data_in[3]
+ scanchain_194/module_data_in[4] scanchain_194/module_data_in[5] scanchain_194/module_data_in[6]
+ scanchain_194/module_data_in[7] scanchain_194/module_data_out[0] scanchain_194/module_data_out[1]
+ scanchain_194/module_data_out[2] scanchain_194/module_data_out[3] scanchain_194/module_data_out[4]
+ scanchain_194/module_data_out[5] scanchain_194/module_data_out[6] scanchain_194/module_data_out[7]
+ scanchain_194/scan_select_in scanchain_195/scan_select_in vccd1 vssd1 scanchain
Xscanchain_172 scanchain_172/clk_in scanchain_173/clk_in scanchain_172/data_in scanchain_173/data_in
+ scanchain_172/latch_enable_in scanchain_173/latch_enable_in scanchain_172/module_data_in[0]
+ scanchain_172/module_data_in[1] scanchain_172/module_data_in[2] scanchain_172/module_data_in[3]
+ scanchain_172/module_data_in[4] scanchain_172/module_data_in[5] scanchain_172/module_data_in[6]
+ scanchain_172/module_data_in[7] scanchain_172/module_data_out[0] scanchain_172/module_data_out[1]
+ scanchain_172/module_data_out[2] scanchain_172/module_data_out[3] scanchain_172/module_data_out[4]
+ scanchain_172/module_data_out[5] scanchain_172/module_data_out[6] scanchain_172/module_data_out[7]
+ scanchain_172/scan_select_in scanchain_173/scan_select_in vccd1 vssd1 scanchain
Xscanchain_183 scanchain_183/clk_in scanchain_184/clk_in scanchain_183/data_in scanchain_184/data_in
+ scanchain_183/latch_enable_in scanchain_184/latch_enable_in scanchain_183/module_data_in[0]
+ scanchain_183/module_data_in[1] scanchain_183/module_data_in[2] scanchain_183/module_data_in[3]
+ scanchain_183/module_data_in[4] scanchain_183/module_data_in[5] scanchain_183/module_data_in[6]
+ scanchain_183/module_data_in[7] scanchain_183/module_data_out[0] scanchain_183/module_data_out[1]
+ scanchain_183/module_data_out[2] scanchain_183/module_data_out[3] scanchain_183/module_data_out[4]
+ scanchain_183/module_data_out[5] scanchain_183/module_data_out[6] scanchain_183/module_data_out[7]
+ scanchain_183/scan_select_in scanchain_184/scan_select_in vccd1 vssd1 scanchain
Xuser_module_348255968419643987_032 scanchain_032/module_data_in[0] scanchain_032/module_data_in[1]
+ scanchain_032/module_data_in[2] scanchain_032/module_data_in[3] scanchain_032/module_data_in[4]
+ scanchain_032/module_data_in[5] scanchain_032/module_data_in[6] scanchain_032/module_data_in[7]
+ scanchain_032/module_data_out[0] scanchain_032/module_data_out[1] scanchain_032/module_data_out[2]
+ scanchain_032/module_data_out[3] scanchain_032/module_data_out[4] scanchain_032/module_data_out[5]
+ scanchain_032/module_data_out[6] scanchain_032/module_data_out[7] vccd1 vssd1 user_module_348255968419643987
Xuser_module_341535056611770964_199 scanchain_199/module_data_in[0] scanchain_199/module_data_in[1]
+ scanchain_199/module_data_in[2] scanchain_199/module_data_in[3] scanchain_199/module_data_in[4]
+ scanchain_199/module_data_in[5] scanchain_199/module_data_in[6] scanchain_199/module_data_in[7]
+ scanchain_199/module_data_out[0] scanchain_199/module_data_out[1] scanchain_199/module_data_out[2]
+ scanchain_199/module_data_out[3] scanchain_199/module_data_out[4] scanchain_199/module_data_out[5]
+ scanchain_199/module_data_out[6] scanchain_199/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xxor_shift32_quantamhd_052 scanchain_052/module_data_in[0] scanchain_052/module_data_in[1]
+ scanchain_052/module_data_in[2] scanchain_052/module_data_in[3] scanchain_052/module_data_in[4]
+ scanchain_052/module_data_in[5] scanchain_052/module_data_in[6] scanchain_052/module_data_in[7]
+ scanchain_052/module_data_out[0] scanchain_052/module_data_out[1] scanchain_052/module_data_out[2]
+ scanchain_052/module_data_out[3] scanchain_052/module_data_out[4] scanchain_052/module_data_out[5]
+ scanchain_052/module_data_out[6] scanchain_052/module_data_out[7] vccd1 vssd1 xor_shift32_quantamhd
Xuser_module_341535056611770964_100 scanchain_100/module_data_in[0] scanchain_100/module_data_in[1]
+ scanchain_100/module_data_in[2] scanchain_100/module_data_in[3] scanchain_100/module_data_in[4]
+ scanchain_100/module_data_in[5] scanchain_100/module_data_in[6] scanchain_100/module_data_in[7]
+ scanchain_100/module_data_out[0] scanchain_100/module_data_out[1] scanchain_100/module_data_out[2]
+ scanchain_100/module_data_out[3] scanchain_100/module_data_out[4] scanchain_100/module_data_out[5]
+ scanchain_100/module_data_out[6] scanchain_100/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_111 scanchain_111/module_data_in[0] scanchain_111/module_data_in[1]
+ scanchain_111/module_data_in[2] scanchain_111/module_data_in[3] scanchain_111/module_data_in[4]
+ scanchain_111/module_data_in[5] scanchain_111/module_data_in[6] scanchain_111/module_data_in[7]
+ scanchain_111/module_data_out[0] scanchain_111/module_data_out[1] scanchain_111/module_data_out[2]
+ scanchain_111/module_data_out[3] scanchain_111/module_data_out[4] scanchain_111/module_data_out[5]
+ scanchain_111/module_data_out[6] scanchain_111/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_122 scanchain_122/module_data_in[0] scanchain_122/module_data_in[1]
+ scanchain_122/module_data_in[2] scanchain_122/module_data_in[3] scanchain_122/module_data_in[4]
+ scanchain_122/module_data_in[5] scanchain_122/module_data_in[6] scanchain_122/module_data_in[7]
+ scanchain_122/module_data_out[0] scanchain_122/module_data_out[1] scanchain_122/module_data_out[2]
+ scanchain_122/module_data_out[3] scanchain_122/module_data_out[4] scanchain_122/module_data_out[5]
+ scanchain_122/module_data_out[6] scanchain_122/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_133 scanchain_133/module_data_in[0] scanchain_133/module_data_in[1]
+ scanchain_133/module_data_in[2] scanchain_133/module_data_in[3] scanchain_133/module_data_in[4]
+ scanchain_133/module_data_in[5] scanchain_133/module_data_in[6] scanchain_133/module_data_in[7]
+ scanchain_133/module_data_out[0] scanchain_133/module_data_out[1] scanchain_133/module_data_out[2]
+ scanchain_133/module_data_out[3] scanchain_133/module_data_out[4] scanchain_133/module_data_out[5]
+ scanchain_133/module_data_out[6] scanchain_133/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_144 scanchain_144/module_data_in[0] scanchain_144/module_data_in[1]
+ scanchain_144/module_data_in[2] scanchain_144/module_data_in[3] scanchain_144/module_data_in[4]
+ scanchain_144/module_data_in[5] scanchain_144/module_data_in[6] scanchain_144/module_data_in[7]
+ scanchain_144/module_data_out[0] scanchain_144/module_data_out[1] scanchain_144/module_data_out[2]
+ scanchain_144/module_data_out[3] scanchain_144/module_data_out[4] scanchain_144/module_data_out[5]
+ scanchain_144/module_data_out[6] scanchain_144/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_155 scanchain_155/module_data_in[0] scanchain_155/module_data_in[1]
+ scanchain_155/module_data_in[2] scanchain_155/module_data_in[3] scanchain_155/module_data_in[4]
+ scanchain_155/module_data_in[5] scanchain_155/module_data_in[6] scanchain_155/module_data_in[7]
+ scanchain_155/module_data_out[0] scanchain_155/module_data_out[1] scanchain_155/module_data_out[2]
+ scanchain_155/module_data_out[3] scanchain_155/module_data_out[4] scanchain_155/module_data_out[5]
+ scanchain_155/module_data_out[6] scanchain_155/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_166 scanchain_166/module_data_in[0] scanchain_166/module_data_in[1]
+ scanchain_166/module_data_in[2] scanchain_166/module_data_in[3] scanchain_166/module_data_in[4]
+ scanchain_166/module_data_in[5] scanchain_166/module_data_in[6] scanchain_166/module_data_in[7]
+ scanchain_166/module_data_out[0] scanchain_166/module_data_out[1] scanchain_166/module_data_out[2]
+ scanchain_166/module_data_out[3] scanchain_166/module_data_out[4] scanchain_166/module_data_out[5]
+ scanchain_166/module_data_out[6] scanchain_166/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_177 scanchain_177/module_data_in[0] scanchain_177/module_data_in[1]
+ scanchain_177/module_data_in[2] scanchain_177/module_data_in[3] scanchain_177/module_data_in[4]
+ scanchain_177/module_data_in[5] scanchain_177/module_data_in[6] scanchain_177/module_data_in[7]
+ scanchain_177/module_data_out[0] scanchain_177/module_data_out[1] scanchain_177/module_data_out[2]
+ scanchain_177/module_data_out[3] scanchain_177/module_data_out[4] scanchain_177/module_data_out[5]
+ scanchain_177/module_data_out[6] scanchain_177/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_188 scanchain_188/module_data_in[0] scanchain_188/module_data_in[1]
+ scanchain_188/module_data_in[2] scanchain_188/module_data_in[3] scanchain_188/module_data_in[4]
+ scanchain_188/module_data_in[5] scanchain_188/module_data_in[6] scanchain_188/module_data_in[7]
+ scanchain_188/module_data_out[0] scanchain_188/module_data_out[1] scanchain_188/module_data_out[2]
+ scanchain_188/module_data_out[3] scanchain_188/module_data_out[4] scanchain_188/module_data_out[5]
+ scanchain_188/module_data_out[6] scanchain_188/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xtomkeddie_top_tto_002 tomkeddie_top_tto_002/io_in[0] tomkeddie_top_tto_002/io_in[1]
+ tomkeddie_top_tto_002/io_in[2] tomkeddie_top_tto_002/io_in[3] tomkeddie_top_tto_002/io_in[4]
+ tomkeddie_top_tto_002/io_in[5] tomkeddie_top_tto_002/io_in[6] tomkeddie_top_tto_002/io_in[7]
+ tomkeddie_top_tto_002/io_out[0] tomkeddie_top_tto_002/io_out[1] tomkeddie_top_tto_002/io_out[2]
+ tomkeddie_top_tto_002/io_out[3] tomkeddie_top_tto_002/io_out[4] tomkeddie_top_tto_002/io_out[5]
+ tomkeddie_top_tto_002/io_out[6] tomkeddie_top_tto_002/io_out[7] vccd1 vssd1 tomkeddie_top_tto
Xscanchain_195 scanchain_195/clk_in scanchain_196/clk_in scanchain_195/data_in scanchain_196/data_in
+ scanchain_195/latch_enable_in scanchain_196/latch_enable_in scanchain_195/module_data_in[0]
+ scanchain_195/module_data_in[1] scanchain_195/module_data_in[2] scanchain_195/module_data_in[3]
+ scanchain_195/module_data_in[4] scanchain_195/module_data_in[5] scanchain_195/module_data_in[6]
+ scanchain_195/module_data_in[7] scanchain_195/module_data_out[0] scanchain_195/module_data_out[1]
+ scanchain_195/module_data_out[2] scanchain_195/module_data_out[3] scanchain_195/module_data_out[4]
+ scanchain_195/module_data_out[5] scanchain_195/module_data_out[6] scanchain_195/module_data_out[7]
+ scanchain_195/scan_select_in scanchain_196/scan_select_in vccd1 vssd1 scanchain
Xscanchain_140 scanchain_140/clk_in scanchain_141/clk_in scanchain_140/data_in scanchain_141/data_in
+ scanchain_140/latch_enable_in scanchain_141/latch_enable_in scanchain_140/module_data_in[0]
+ scanchain_140/module_data_in[1] scanchain_140/module_data_in[2] scanchain_140/module_data_in[3]
+ scanchain_140/module_data_in[4] scanchain_140/module_data_in[5] scanchain_140/module_data_in[6]
+ scanchain_140/module_data_in[7] scanchain_140/module_data_out[0] scanchain_140/module_data_out[1]
+ scanchain_140/module_data_out[2] scanchain_140/module_data_out[3] scanchain_140/module_data_out[4]
+ scanchain_140/module_data_out[5] scanchain_140/module_data_out[6] scanchain_140/module_data_out[7]
+ scanchain_140/scan_select_in scanchain_141/scan_select_in vccd1 vssd1 scanchain
Xscanchain_151 scanchain_151/clk_in scanchain_152/clk_in scanchain_151/data_in scanchain_152/data_in
+ scanchain_151/latch_enable_in scanchain_152/latch_enable_in scanchain_151/module_data_in[0]
+ scanchain_151/module_data_in[1] scanchain_151/module_data_in[2] scanchain_151/module_data_in[3]
+ scanchain_151/module_data_in[4] scanchain_151/module_data_in[5] scanchain_151/module_data_in[6]
+ scanchain_151/module_data_in[7] scanchain_151/module_data_out[0] scanchain_151/module_data_out[1]
+ scanchain_151/module_data_out[2] scanchain_151/module_data_out[3] scanchain_151/module_data_out[4]
+ scanchain_151/module_data_out[5] scanchain_151/module_data_out[6] scanchain_151/module_data_out[7]
+ scanchain_151/scan_select_in scanchain_152/scan_select_in vccd1 vssd1 scanchain
Xscanchain_162 scanchain_162/clk_in scanchain_163/clk_in scanchain_162/data_in scanchain_163/data_in
+ scanchain_162/latch_enable_in scanchain_163/latch_enable_in scanchain_162/module_data_in[0]
+ scanchain_162/module_data_in[1] scanchain_162/module_data_in[2] scanchain_162/module_data_in[3]
+ scanchain_162/module_data_in[4] scanchain_162/module_data_in[5] scanchain_162/module_data_in[6]
+ scanchain_162/module_data_in[7] scanchain_162/module_data_out[0] scanchain_162/module_data_out[1]
+ scanchain_162/module_data_out[2] scanchain_162/module_data_out[3] scanchain_162/module_data_out[4]
+ scanchain_162/module_data_out[5] scanchain_162/module_data_out[6] scanchain_162/module_data_out[7]
+ scanchain_162/scan_select_in scanchain_163/scan_select_in vccd1 vssd1 scanchain
Xscanchain_173 scanchain_173/clk_in scanchain_174/clk_in scanchain_173/data_in scanchain_174/data_in
+ scanchain_173/latch_enable_in scanchain_174/latch_enable_in scanchain_173/module_data_in[0]
+ scanchain_173/module_data_in[1] scanchain_173/module_data_in[2] scanchain_173/module_data_in[3]
+ scanchain_173/module_data_in[4] scanchain_173/module_data_in[5] scanchain_173/module_data_in[6]
+ scanchain_173/module_data_in[7] scanchain_173/module_data_out[0] scanchain_173/module_data_out[1]
+ scanchain_173/module_data_out[2] scanchain_173/module_data_out[3] scanchain_173/module_data_out[4]
+ scanchain_173/module_data_out[5] scanchain_173/module_data_out[6] scanchain_173/module_data_out[7]
+ scanchain_173/scan_select_in scanchain_174/scan_select_in vccd1 vssd1 scanchain
Xscanchain_184 scanchain_184/clk_in scanchain_185/clk_in scanchain_184/data_in scanchain_185/data_in
+ scanchain_184/latch_enable_in scanchain_185/latch_enable_in scanchain_184/module_data_in[0]
+ scanchain_184/module_data_in[1] scanchain_184/module_data_in[2] scanchain_184/module_data_in[3]
+ scanchain_184/module_data_in[4] scanchain_184/module_data_in[5] scanchain_184/module_data_in[6]
+ scanchain_184/module_data_in[7] scanchain_184/module_data_out[0] scanchain_184/module_data_out[1]
+ scanchain_184/module_data_out[2] scanchain_184/module_data_out[3] scanchain_184/module_data_out[4]
+ scanchain_184/module_data_out[5] scanchain_184/module_data_out[6] scanchain_184/module_data_out[7]
+ scanchain_184/scan_select_in scanchain_185/scan_select_in vccd1 vssd1 scanchain
Xtholin_avalonsemi_5401_014 scanchain_014/module_data_in[0] scanchain_014/module_data_in[1]
+ scanchain_014/module_data_in[2] scanchain_014/module_data_in[3] scanchain_014/module_data_in[4]
+ scanchain_014/module_data_in[5] scanchain_014/module_data_in[6] scanchain_014/module_data_in[7]
+ scanchain_014/module_data_out[0] scanchain_014/module_data_out[1] scanchain_014/module_data_out[2]
+ scanchain_014/module_data_out[3] scanchain_014/module_data_out[4] scanchain_014/module_data_out[5]
+ scanchain_014/module_data_out[6] scanchain_014/module_data_out[7] vccd1 vssd1 tholin_avalonsemi_5401
XAidanMedcalf_pid_controller_075 scanchain_075/module_data_in[0] scanchain_075/module_data_in[1]
+ scanchain_075/module_data_in[2] scanchain_075/module_data_in[3] scanchain_075/module_data_in[4]
+ scanchain_075/module_data_in[5] scanchain_075/module_data_in[6] scanchain_075/module_data_in[7]
+ scanchain_075/module_data_out[0] scanchain_075/module_data_out[1] scanchain_075/module_data_out[2]
+ scanchain_075/module_data_out[3] scanchain_075/module_data_out[4] scanchain_075/module_data_out[5]
+ scanchain_075/module_data_out[6] scanchain_075/module_data_out[7] vccd1 vssd1 AidanMedcalf_pid_controller
Xuser_module_348381622440034899_083 scanchain_083/module_data_in[0] scanchain_083/module_data_in[1]
+ scanchain_083/module_data_in[2] scanchain_083/module_data_in[3] scanchain_083/module_data_in[4]
+ scanchain_083/module_data_in[5] scanchain_083/module_data_in[6] scanchain_083/module_data_in[7]
+ scanchain_083/module_data_out[0] scanchain_083/module_data_out[1] scanchain_083/module_data_out[2]
+ scanchain_083/module_data_out[3] scanchain_083/module_data_out[4] scanchain_083/module_data_out[5]
+ scanchain_083/module_data_out[6] scanchain_083/module_data_out[7] vccd1 vssd1 user_module_348381622440034899
Xuser_module_341535056611770964_101 scanchain_101/module_data_in[0] scanchain_101/module_data_in[1]
+ scanchain_101/module_data_in[2] scanchain_101/module_data_in[3] scanchain_101/module_data_in[4]
+ scanchain_101/module_data_in[5] scanchain_101/module_data_in[6] scanchain_101/module_data_in[7]
+ scanchain_101/module_data_out[0] scanchain_101/module_data_out[1] scanchain_101/module_data_out[2]
+ scanchain_101/module_data_out[3] scanchain_101/module_data_out[4] scanchain_101/module_data_out[5]
+ scanchain_101/module_data_out[6] scanchain_101/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_112 scanchain_112/module_data_in[0] scanchain_112/module_data_in[1]
+ scanchain_112/module_data_in[2] scanchain_112/module_data_in[3] scanchain_112/module_data_in[4]
+ scanchain_112/module_data_in[5] scanchain_112/module_data_in[6] scanchain_112/module_data_in[7]
+ scanchain_112/module_data_out[0] scanchain_112/module_data_out[1] scanchain_112/module_data_out[2]
+ scanchain_112/module_data_out[3] scanchain_112/module_data_out[4] scanchain_112/module_data_out[5]
+ scanchain_112/module_data_out[6] scanchain_112/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_123 scanchain_123/module_data_in[0] scanchain_123/module_data_in[1]
+ scanchain_123/module_data_in[2] scanchain_123/module_data_in[3] scanchain_123/module_data_in[4]
+ scanchain_123/module_data_in[5] scanchain_123/module_data_in[6] scanchain_123/module_data_in[7]
+ scanchain_123/module_data_out[0] scanchain_123/module_data_out[1] scanchain_123/module_data_out[2]
+ scanchain_123/module_data_out[3] scanchain_123/module_data_out[4] scanchain_123/module_data_out[5]
+ scanchain_123/module_data_out[6] scanchain_123/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_134 scanchain_134/module_data_in[0] scanchain_134/module_data_in[1]
+ scanchain_134/module_data_in[2] scanchain_134/module_data_in[3] scanchain_134/module_data_in[4]
+ scanchain_134/module_data_in[5] scanchain_134/module_data_in[6] scanchain_134/module_data_in[7]
+ scanchain_134/module_data_out[0] scanchain_134/module_data_out[1] scanchain_134/module_data_out[2]
+ scanchain_134/module_data_out[3] scanchain_134/module_data_out[4] scanchain_134/module_data_out[5]
+ scanchain_134/module_data_out[6] scanchain_134/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_145 scanchain_145/module_data_in[0] scanchain_145/module_data_in[1]
+ scanchain_145/module_data_in[2] scanchain_145/module_data_in[3] scanchain_145/module_data_in[4]
+ scanchain_145/module_data_in[5] scanchain_145/module_data_in[6] scanchain_145/module_data_in[7]
+ scanchain_145/module_data_out[0] scanchain_145/module_data_out[1] scanchain_145/module_data_out[2]
+ scanchain_145/module_data_out[3] scanchain_145/module_data_out[4] scanchain_145/module_data_out[5]
+ scanchain_145/module_data_out[6] scanchain_145/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_156 scanchain_156/module_data_in[0] scanchain_156/module_data_in[1]
+ scanchain_156/module_data_in[2] scanchain_156/module_data_in[3] scanchain_156/module_data_in[4]
+ scanchain_156/module_data_in[5] scanchain_156/module_data_in[6] scanchain_156/module_data_in[7]
+ scanchain_156/module_data_out[0] scanchain_156/module_data_out[1] scanchain_156/module_data_out[2]
+ scanchain_156/module_data_out[3] scanchain_156/module_data_out[4] scanchain_156/module_data_out[5]
+ scanchain_156/module_data_out[6] scanchain_156/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_167 scanchain_167/module_data_in[0] scanchain_167/module_data_in[1]
+ scanchain_167/module_data_in[2] scanchain_167/module_data_in[3] scanchain_167/module_data_in[4]
+ scanchain_167/module_data_in[5] scanchain_167/module_data_in[6] scanchain_167/module_data_in[7]
+ scanchain_167/module_data_out[0] scanchain_167/module_data_out[1] scanchain_167/module_data_out[2]
+ scanchain_167/module_data_out[3] scanchain_167/module_data_out[4] scanchain_167/module_data_out[5]
+ scanchain_167/module_data_out[6] scanchain_167/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_178 scanchain_178/module_data_in[0] scanchain_178/module_data_in[1]
+ scanchain_178/module_data_in[2] scanchain_178/module_data_in[3] scanchain_178/module_data_in[4]
+ scanchain_178/module_data_in[5] scanchain_178/module_data_in[6] scanchain_178/module_data_in[7]
+ scanchain_178/module_data_out[0] scanchain_178/module_data_out[1] scanchain_178/module_data_out[2]
+ scanchain_178/module_data_out[3] scanchain_178/module_data_out[4] scanchain_178/module_data_out[5]
+ scanchain_178/module_data_out[6] scanchain_178/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_189 scanchain_189/module_data_in[0] scanchain_189/module_data_in[1]
+ scanchain_189/module_data_in[2] scanchain_189/module_data_in[3] scanchain_189/module_data_in[4]
+ scanchain_189/module_data_in[5] scanchain_189/module_data_in[6] scanchain_189/module_data_in[7]
+ scanchain_189/module_data_out[0] scanchain_189/module_data_out[1] scanchain_189/module_data_out[2]
+ scanchain_189/module_data_out[3] scanchain_189/module_data_out[4] scanchain_189/module_data_out[5]
+ scanchain_189/module_data_out[6] scanchain_189/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_196 scanchain_196/clk_in scanchain_197/clk_in scanchain_196/data_in scanchain_197/data_in
+ scanchain_196/latch_enable_in scanchain_197/latch_enable_in scanchain_196/module_data_in[0]
+ scanchain_196/module_data_in[1] scanchain_196/module_data_in[2] scanchain_196/module_data_in[3]
+ scanchain_196/module_data_in[4] scanchain_196/module_data_in[5] scanchain_196/module_data_in[6]
+ scanchain_196/module_data_in[7] scanchain_196/module_data_out[0] scanchain_196/module_data_out[1]
+ scanchain_196/module_data_out[2] scanchain_196/module_data_out[3] scanchain_196/module_data_out[4]
+ scanchain_196/module_data_out[5] scanchain_196/module_data_out[6] scanchain_196/module_data_out[7]
+ scanchain_196/scan_select_in scanchain_197/scan_select_in vccd1 vssd1 scanchain
Xscanchain_130 scanchain_130/clk_in scanchain_131/clk_in scanchain_130/data_in scanchain_131/data_in
+ scanchain_130/latch_enable_in scanchain_131/latch_enable_in scanchain_130/module_data_in[0]
+ scanchain_130/module_data_in[1] scanchain_130/module_data_in[2] scanchain_130/module_data_in[3]
+ scanchain_130/module_data_in[4] scanchain_130/module_data_in[5] scanchain_130/module_data_in[6]
+ scanchain_130/module_data_in[7] scanchain_130/module_data_out[0] scanchain_130/module_data_out[1]
+ scanchain_130/module_data_out[2] scanchain_130/module_data_out[3] scanchain_130/module_data_out[4]
+ scanchain_130/module_data_out[5] scanchain_130/module_data_out[6] scanchain_130/module_data_out[7]
+ scanchain_130/scan_select_in scanchain_131/scan_select_in vccd1 vssd1 scanchain
Xscanchain_141 scanchain_141/clk_in scanchain_142/clk_in scanchain_141/data_in scanchain_142/data_in
+ scanchain_141/latch_enable_in scanchain_142/latch_enable_in scanchain_141/module_data_in[0]
+ scanchain_141/module_data_in[1] scanchain_141/module_data_in[2] scanchain_141/module_data_in[3]
+ scanchain_141/module_data_in[4] scanchain_141/module_data_in[5] scanchain_141/module_data_in[6]
+ scanchain_141/module_data_in[7] scanchain_141/module_data_out[0] scanchain_141/module_data_out[1]
+ scanchain_141/module_data_out[2] scanchain_141/module_data_out[3] scanchain_141/module_data_out[4]
+ scanchain_141/module_data_out[5] scanchain_141/module_data_out[6] scanchain_141/module_data_out[7]
+ scanchain_141/scan_select_in scanchain_142/scan_select_in vccd1 vssd1 scanchain
Xscanchain_163 scanchain_163/clk_in scanchain_164/clk_in scanchain_163/data_in scanchain_164/data_in
+ scanchain_163/latch_enable_in scanchain_164/latch_enable_in scanchain_163/module_data_in[0]
+ scanchain_163/module_data_in[1] scanchain_163/module_data_in[2] scanchain_163/module_data_in[3]
+ scanchain_163/module_data_in[4] scanchain_163/module_data_in[5] scanchain_163/module_data_in[6]
+ scanchain_163/module_data_in[7] scanchain_163/module_data_out[0] scanchain_163/module_data_out[1]
+ scanchain_163/module_data_out[2] scanchain_163/module_data_out[3] scanchain_163/module_data_out[4]
+ scanchain_163/module_data_out[5] scanchain_163/module_data_out[6] scanchain_163/module_data_out[7]
+ scanchain_163/scan_select_in scanchain_164/scan_select_in vccd1 vssd1 scanchain
Xscanchain_152 scanchain_152/clk_in scanchain_153/clk_in scanchain_152/data_in scanchain_153/data_in
+ scanchain_152/latch_enable_in scanchain_153/latch_enable_in scanchain_152/module_data_in[0]
+ scanchain_152/module_data_in[1] scanchain_152/module_data_in[2] scanchain_152/module_data_in[3]
+ scanchain_152/module_data_in[4] scanchain_152/module_data_in[5] scanchain_152/module_data_in[6]
+ scanchain_152/module_data_in[7] scanchain_152/module_data_out[0] scanchain_152/module_data_out[1]
+ scanchain_152/module_data_out[2] scanchain_152/module_data_out[3] scanchain_152/module_data_out[4]
+ scanchain_152/module_data_out[5] scanchain_152/module_data_out[6] scanchain_152/module_data_out[7]
+ scanchain_152/scan_select_in scanchain_153/scan_select_in vccd1 vssd1 scanchain
Xscanchain_174 scanchain_174/clk_in scanchain_175/clk_in scanchain_174/data_in scanchain_175/data_in
+ scanchain_174/latch_enable_in scanchain_175/latch_enable_in scanchain_174/module_data_in[0]
+ scanchain_174/module_data_in[1] scanchain_174/module_data_in[2] scanchain_174/module_data_in[3]
+ scanchain_174/module_data_in[4] scanchain_174/module_data_in[5] scanchain_174/module_data_in[6]
+ scanchain_174/module_data_in[7] scanchain_174/module_data_out[0] scanchain_174/module_data_out[1]
+ scanchain_174/module_data_out[2] scanchain_174/module_data_out[3] scanchain_174/module_data_out[4]
+ scanchain_174/module_data_out[5] scanchain_174/module_data_out[6] scanchain_174/module_data_out[7]
+ scanchain_174/scan_select_in scanchain_175/scan_select_in vccd1 vssd1 scanchain
Xscanchain_185 scanchain_185/clk_in scanchain_186/clk_in scanchain_185/data_in scanchain_186/data_in
+ scanchain_185/latch_enable_in scanchain_186/latch_enable_in scanchain_185/module_data_in[0]
+ scanchain_185/module_data_in[1] scanchain_185/module_data_in[2] scanchain_185/module_data_in[3]
+ scanchain_185/module_data_in[4] scanchain_185/module_data_in[5] scanchain_185/module_data_in[6]
+ scanchain_185/module_data_in[7] scanchain_185/module_data_out[0] scanchain_185/module_data_out[1]
+ scanchain_185/module_data_out[2] scanchain_185/module_data_out[3] scanchain_185/module_data_out[4]
+ scanchain_185/module_data_out[5] scanchain_185/module_data_out[6] scanchain_185/module_data_out[7]
+ scanchain_185/scan_select_in scanchain_186/scan_select_in vccd1 vssd1 scanchain
Xericsmi_speed_test_074 scanchain_074/module_data_in[0] scanchain_074/module_data_in[1]
+ scanchain_074/module_data_in[2] scanchain_074/module_data_in[3] scanchain_074/module_data_in[4]
+ scanchain_074/module_data_in[5] scanchain_074/module_data_in[6] scanchain_074/module_data_in[7]
+ scanchain_074/module_data_out[0] scanchain_074/module_data_out[1] scanchain_074/module_data_out[2]
+ scanchain_074/module_data_out[3] scanchain_074/module_data_out[4] scanchain_074/module_data_out[5]
+ scanchain_074/module_data_out[6] scanchain_074/module_data_out[7] vccd1 vssd1 ericsmi_speed_test
Xaramsey118_freq_counter_087 scanchain_087/module_data_in[0] scanchain_087/module_data_in[1]
+ scanchain_087/module_data_in[2] scanchain_087/module_data_in[3] scanchain_087/module_data_in[4]
+ scanchain_087/module_data_in[5] scanchain_087/module_data_in[6] scanchain_087/module_data_in[7]
+ scanchain_087/module_data_out[0] scanchain_087/module_data_out[1] scanchain_087/module_data_out[2]
+ scanchain_087/module_data_out[3] scanchain_087/module_data_out[4] scanchain_087/module_data_out[5]
+ scanchain_087/module_data_out[6] scanchain_087/module_data_out[7] vccd1 vssd1 aramsey118_freq_counter
Xuser_module_341423712597181012_093 scanchain_093/module_data_in[0] scanchain_093/module_data_in[1]
+ scanchain_093/module_data_in[2] scanchain_093/module_data_in[3] scanchain_093/module_data_in[4]
+ scanchain_093/module_data_in[5] scanchain_093/module_data_in[6] scanchain_093/module_data_in[7]
+ scanchain_093/module_data_out[0] scanchain_093/module_data_out[1] scanchain_093/module_data_out[2]
+ scanchain_093/module_data_out[3] scanchain_093/module_data_out[4] scanchain_093/module_data_out[5]
+ scanchain_093/module_data_out[6] scanchain_093/module_data_out[7] vccd1 vssd1 user_module_341423712597181012
Xuser_module_341535056611770964_102 scanchain_102/module_data_in[0] scanchain_102/module_data_in[1]
+ scanchain_102/module_data_in[2] scanchain_102/module_data_in[3] scanchain_102/module_data_in[4]
+ scanchain_102/module_data_in[5] scanchain_102/module_data_in[6] scanchain_102/module_data_in[7]
+ scanchain_102/module_data_out[0] scanchain_102/module_data_out[1] scanchain_102/module_data_out[2]
+ scanchain_102/module_data_out[3] scanchain_102/module_data_out[4] scanchain_102/module_data_out[5]
+ scanchain_102/module_data_out[6] scanchain_102/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_113 scanchain_113/module_data_in[0] scanchain_113/module_data_in[1]
+ scanchain_113/module_data_in[2] scanchain_113/module_data_in[3] scanchain_113/module_data_in[4]
+ scanchain_113/module_data_in[5] scanchain_113/module_data_in[6] scanchain_113/module_data_in[7]
+ scanchain_113/module_data_out[0] scanchain_113/module_data_out[1] scanchain_113/module_data_out[2]
+ scanchain_113/module_data_out[3] scanchain_113/module_data_out[4] scanchain_113/module_data_out[5]
+ scanchain_113/module_data_out[6] scanchain_113/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_135 scanchain_135/module_data_in[0] scanchain_135/module_data_in[1]
+ scanchain_135/module_data_in[2] scanchain_135/module_data_in[3] scanchain_135/module_data_in[4]
+ scanchain_135/module_data_in[5] scanchain_135/module_data_in[6] scanchain_135/module_data_in[7]
+ scanchain_135/module_data_out[0] scanchain_135/module_data_out[1] scanchain_135/module_data_out[2]
+ scanchain_135/module_data_out[3] scanchain_135/module_data_out[4] scanchain_135/module_data_out[5]
+ scanchain_135/module_data_out[6] scanchain_135/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_124 scanchain_124/module_data_in[0] scanchain_124/module_data_in[1]
+ scanchain_124/module_data_in[2] scanchain_124/module_data_in[3] scanchain_124/module_data_in[4]
+ scanchain_124/module_data_in[5] scanchain_124/module_data_in[6] scanchain_124/module_data_in[7]
+ scanchain_124/module_data_out[0] scanchain_124/module_data_out[1] scanchain_124/module_data_out[2]
+ scanchain_124/module_data_out[3] scanchain_124/module_data_out[4] scanchain_124/module_data_out[5]
+ scanchain_124/module_data_out[6] scanchain_124/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_146 scanchain_146/module_data_in[0] scanchain_146/module_data_in[1]
+ scanchain_146/module_data_in[2] scanchain_146/module_data_in[3] scanchain_146/module_data_in[4]
+ scanchain_146/module_data_in[5] scanchain_146/module_data_in[6] scanchain_146/module_data_in[7]
+ scanchain_146/module_data_out[0] scanchain_146/module_data_out[1] scanchain_146/module_data_out[2]
+ scanchain_146/module_data_out[3] scanchain_146/module_data_out[4] scanchain_146/module_data_out[5]
+ scanchain_146/module_data_out[6] scanchain_146/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_157 scanchain_157/module_data_in[0] scanchain_157/module_data_in[1]
+ scanchain_157/module_data_in[2] scanchain_157/module_data_in[3] scanchain_157/module_data_in[4]
+ scanchain_157/module_data_in[5] scanchain_157/module_data_in[6] scanchain_157/module_data_in[7]
+ scanchain_157/module_data_out[0] scanchain_157/module_data_out[1] scanchain_157/module_data_out[2]
+ scanchain_157/module_data_out[3] scanchain_157/module_data_out[4] scanchain_157/module_data_out[5]
+ scanchain_157/module_data_out[6] scanchain_157/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_168 scanchain_168/module_data_in[0] scanchain_168/module_data_in[1]
+ scanchain_168/module_data_in[2] scanchain_168/module_data_in[3] scanchain_168/module_data_in[4]
+ scanchain_168/module_data_in[5] scanchain_168/module_data_in[6] scanchain_168/module_data_in[7]
+ scanchain_168/module_data_out[0] scanchain_168/module_data_out[1] scanchain_168/module_data_out[2]
+ scanchain_168/module_data_out[3] scanchain_168/module_data_out[4] scanchain_168/module_data_out[5]
+ scanchain_168/module_data_out[6] scanchain_168/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_179 scanchain_179/module_data_in[0] scanchain_179/module_data_in[1]
+ scanchain_179/module_data_in[2] scanchain_179/module_data_in[3] scanchain_179/module_data_in[4]
+ scanchain_179/module_data_in[5] scanchain_179/module_data_in[6] scanchain_179/module_data_in[7]
+ scanchain_179/module_data_out[0] scanchain_179/module_data_out[1] scanchain_179/module_data_out[2]
+ scanchain_179/module_data_out[3] scanchain_179/module_data_out[4] scanchain_179/module_data_out[5]
+ scanchain_179/module_data_out[6] scanchain_179/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_348121131386929746_028 scanchain_028/module_data_in[0] scanchain_028/module_data_in[1]
+ scanchain_028/module_data_in[2] scanchain_028/module_data_in[3] scanchain_028/module_data_in[4]
+ scanchain_028/module_data_in[5] scanchain_028/module_data_in[6] scanchain_028/module_data_in[7]
+ scanchain_028/module_data_out[0] scanchain_028/module_data_out[1] scanchain_028/module_data_out[2]
+ scanchain_028/module_data_out[3] scanchain_028/module_data_out[4] scanchain_028/module_data_out[5]
+ scanchain_028/module_data_out[6] scanchain_028/module_data_out[7] vccd1 vssd1 user_module_348121131386929746
Xuser_module_341620484740219475_041 scanchain_041/module_data_in[0] scanchain_041/module_data_in[1]
+ scanchain_041/module_data_in[2] scanchain_041/module_data_in[3] scanchain_041/module_data_in[4]
+ scanchain_041/module_data_in[5] scanchain_041/module_data_in[6] scanchain_041/module_data_in[7]
+ scanchain_041/module_data_out[0] scanchain_041/module_data_out[1] scanchain_041/module_data_out[2]
+ scanchain_041/module_data_out[3] scanchain_041/module_data_out[4] scanchain_041/module_data_out[5]
+ scanchain_041/module_data_out[6] scanchain_041/module_data_out[7] vccd1 vssd1 user_module_341620484740219475
Xscanchain_197 scanchain_197/clk_in scanchain_198/clk_in scanchain_197/data_in scanchain_198/data_in
+ scanchain_197/latch_enable_in scanchain_198/latch_enable_in scanchain_197/module_data_in[0]
+ scanchain_197/module_data_in[1] scanchain_197/module_data_in[2] scanchain_197/module_data_in[3]
+ scanchain_197/module_data_in[4] scanchain_197/module_data_in[5] scanchain_197/module_data_in[6]
+ scanchain_197/module_data_in[7] scanchain_197/module_data_out[0] scanchain_197/module_data_out[1]
+ scanchain_197/module_data_out[2] scanchain_197/module_data_out[3] scanchain_197/module_data_out[4]
+ scanchain_197/module_data_out[5] scanchain_197/module_data_out[6] scanchain_197/module_data_out[7]
+ scanchain_197/scan_select_in scanchain_198/scan_select_in vccd1 vssd1 scanchain
Xuser_module_347619669052490324_056 scanchain_056/module_data_in[0] scanchain_056/module_data_in[1]
+ scanchain_056/module_data_in[2] scanchain_056/module_data_in[3] scanchain_056/module_data_in[4]
+ scanchain_056/module_data_in[5] scanchain_056/module_data_in[6] scanchain_056/module_data_in[7]
+ scanchain_056/module_data_out[0] scanchain_056/module_data_out[1] scanchain_056/module_data_out[2]
+ scanchain_056/module_data_out[3] scanchain_056/module_data_out[4] scanchain_056/module_data_out[5]
+ scanchain_056/module_data_out[6] scanchain_056/module_data_out[7] vccd1 vssd1 user_module_347619669052490324
Xscanchain_120 scanchain_120/clk_in scanchain_121/clk_in scanchain_120/data_in scanchain_121/data_in
+ scanchain_120/latch_enable_in scanchain_121/latch_enable_in scanchain_120/module_data_in[0]
+ scanchain_120/module_data_in[1] scanchain_120/module_data_in[2] scanchain_120/module_data_in[3]
+ scanchain_120/module_data_in[4] scanchain_120/module_data_in[5] scanchain_120/module_data_in[6]
+ scanchain_120/module_data_in[7] scanchain_120/module_data_out[0] scanchain_120/module_data_out[1]
+ scanchain_120/module_data_out[2] scanchain_120/module_data_out[3] scanchain_120/module_data_out[4]
+ scanchain_120/module_data_out[5] scanchain_120/module_data_out[6] scanchain_120/module_data_out[7]
+ scanchain_120/scan_select_in scanchain_121/scan_select_in vccd1 vssd1 scanchain
Xscanchain_131 scanchain_131/clk_in scanchain_132/clk_in scanchain_131/data_in scanchain_132/data_in
+ scanchain_131/latch_enable_in scanchain_132/latch_enable_in scanchain_131/module_data_in[0]
+ scanchain_131/module_data_in[1] scanchain_131/module_data_in[2] scanchain_131/module_data_in[3]
+ scanchain_131/module_data_in[4] scanchain_131/module_data_in[5] scanchain_131/module_data_in[6]
+ scanchain_131/module_data_in[7] scanchain_131/module_data_out[0] scanchain_131/module_data_out[1]
+ scanchain_131/module_data_out[2] scanchain_131/module_data_out[3] scanchain_131/module_data_out[4]
+ scanchain_131/module_data_out[5] scanchain_131/module_data_out[6] scanchain_131/module_data_out[7]
+ scanchain_131/scan_select_in scanchain_132/scan_select_in vccd1 vssd1 scanchain
Xscanchain_142 scanchain_142/clk_in scanchain_143/clk_in scanchain_142/data_in scanchain_143/data_in
+ scanchain_142/latch_enable_in scanchain_143/latch_enable_in scanchain_142/module_data_in[0]
+ scanchain_142/module_data_in[1] scanchain_142/module_data_in[2] scanchain_142/module_data_in[3]
+ scanchain_142/module_data_in[4] scanchain_142/module_data_in[5] scanchain_142/module_data_in[6]
+ scanchain_142/module_data_in[7] scanchain_142/module_data_out[0] scanchain_142/module_data_out[1]
+ scanchain_142/module_data_out[2] scanchain_142/module_data_out[3] scanchain_142/module_data_out[4]
+ scanchain_142/module_data_out[5] scanchain_142/module_data_out[6] scanchain_142/module_data_out[7]
+ scanchain_142/scan_select_in scanchain_143/scan_select_in vccd1 vssd1 scanchain
Xscanchain_164 scanchain_164/clk_in scanchain_165/clk_in scanchain_164/data_in scanchain_165/data_in
+ scanchain_164/latch_enable_in scanchain_165/latch_enable_in scanchain_164/module_data_in[0]
+ scanchain_164/module_data_in[1] scanchain_164/module_data_in[2] scanchain_164/module_data_in[3]
+ scanchain_164/module_data_in[4] scanchain_164/module_data_in[5] scanchain_164/module_data_in[6]
+ scanchain_164/module_data_in[7] scanchain_164/module_data_out[0] scanchain_164/module_data_out[1]
+ scanchain_164/module_data_out[2] scanchain_164/module_data_out[3] scanchain_164/module_data_out[4]
+ scanchain_164/module_data_out[5] scanchain_164/module_data_out[6] scanchain_164/module_data_out[7]
+ scanchain_164/scan_select_in scanchain_165/scan_select_in vccd1 vssd1 scanchain
Xscanchain_153 scanchain_153/clk_in scanchain_154/clk_in scanchain_153/data_in scanchain_154/data_in
+ scanchain_153/latch_enable_in scanchain_154/latch_enable_in scanchain_153/module_data_in[0]
+ scanchain_153/module_data_in[1] scanchain_153/module_data_in[2] scanchain_153/module_data_in[3]
+ scanchain_153/module_data_in[4] scanchain_153/module_data_in[5] scanchain_153/module_data_in[6]
+ scanchain_153/module_data_in[7] scanchain_153/module_data_out[0] scanchain_153/module_data_out[1]
+ scanchain_153/module_data_out[2] scanchain_153/module_data_out[3] scanchain_153/module_data_out[4]
+ scanchain_153/module_data_out[5] scanchain_153/module_data_out[6] scanchain_153/module_data_out[7]
+ scanchain_153/scan_select_in scanchain_154/scan_select_in vccd1 vssd1 scanchain
Xscanchain_175 scanchain_175/clk_in scanchain_176/clk_in scanchain_175/data_in scanchain_176/data_in
+ scanchain_175/latch_enable_in scanchain_176/latch_enable_in scanchain_175/module_data_in[0]
+ scanchain_175/module_data_in[1] scanchain_175/module_data_in[2] scanchain_175/module_data_in[3]
+ scanchain_175/module_data_in[4] scanchain_175/module_data_in[5] scanchain_175/module_data_in[6]
+ scanchain_175/module_data_in[7] scanchain_175/module_data_out[0] scanchain_175/module_data_out[1]
+ scanchain_175/module_data_out[2] scanchain_175/module_data_out[3] scanchain_175/module_data_out[4]
+ scanchain_175/module_data_out[5] scanchain_175/module_data_out[6] scanchain_175/module_data_out[7]
+ scanchain_175/scan_select_in scanchain_176/scan_select_in vccd1 vssd1 scanchain
Xscanchain_186 scanchain_186/clk_in scanchain_187/clk_in scanchain_186/data_in scanchain_187/data_in
+ scanchain_186/latch_enable_in scanchain_187/latch_enable_in scanchain_186/module_data_in[0]
+ scanchain_186/module_data_in[1] scanchain_186/module_data_in[2] scanchain_186/module_data_in[3]
+ scanchain_186/module_data_in[4] scanchain_186/module_data_in[5] scanchain_186/module_data_in[6]
+ scanchain_186/module_data_in[7] scanchain_186/module_data_out[0] scanchain_186/module_data_out[1]
+ scanchain_186/module_data_out[2] scanchain_186/module_data_out[3] scanchain_186/module_data_out[4]
+ scanchain_186/module_data_out[5] scanchain_186/module_data_out[6] scanchain_186/module_data_out[7]
+ scanchain_186/scan_select_in scanchain_187/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_103 scanchain_103/module_data_in[0] scanchain_103/module_data_in[1]
+ scanchain_103/module_data_in[2] scanchain_103/module_data_in[3] scanchain_103/module_data_in[4]
+ scanchain_103/module_data_in[5] scanchain_103/module_data_in[6] scanchain_103/module_data_in[7]
+ scanchain_103/module_data_out[0] scanchain_103/module_data_out[1] scanchain_103/module_data_out[2]
+ scanchain_103/module_data_out[3] scanchain_103/module_data_out[4] scanchain_103/module_data_out[5]
+ scanchain_103/module_data_out[6] scanchain_103/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_114 scanchain_114/module_data_in[0] scanchain_114/module_data_in[1]
+ scanchain_114/module_data_in[2] scanchain_114/module_data_in[3] scanchain_114/module_data_in[4]
+ scanchain_114/module_data_in[5] scanchain_114/module_data_in[6] scanchain_114/module_data_in[7]
+ scanchain_114/module_data_out[0] scanchain_114/module_data_out[1] scanchain_114/module_data_out[2]
+ scanchain_114/module_data_out[3] scanchain_114/module_data_out[4] scanchain_114/module_data_out[5]
+ scanchain_114/module_data_out[6] scanchain_114/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_136 scanchain_136/module_data_in[0] scanchain_136/module_data_in[1]
+ scanchain_136/module_data_in[2] scanchain_136/module_data_in[3] scanchain_136/module_data_in[4]
+ scanchain_136/module_data_in[5] scanchain_136/module_data_in[6] scanchain_136/module_data_in[7]
+ scanchain_136/module_data_out[0] scanchain_136/module_data_out[1] scanchain_136/module_data_out[2]
+ scanchain_136/module_data_out[3] scanchain_136/module_data_out[4] scanchain_136/module_data_out[5]
+ scanchain_136/module_data_out[6] scanchain_136/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_125 scanchain_125/module_data_in[0] scanchain_125/module_data_in[1]
+ scanchain_125/module_data_in[2] scanchain_125/module_data_in[3] scanchain_125/module_data_in[4]
+ scanchain_125/module_data_in[5] scanchain_125/module_data_in[6] scanchain_125/module_data_in[7]
+ scanchain_125/module_data_out[0] scanchain_125/module_data_out[1] scanchain_125/module_data_out[2]
+ scanchain_125/module_data_out[3] scanchain_125/module_data_out[4] scanchain_125/module_data_out[5]
+ scanchain_125/module_data_out[6] scanchain_125/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_147 scanchain_147/module_data_in[0] scanchain_147/module_data_in[1]
+ scanchain_147/module_data_in[2] scanchain_147/module_data_in[3] scanchain_147/module_data_in[4]
+ scanchain_147/module_data_in[5] scanchain_147/module_data_in[6] scanchain_147/module_data_in[7]
+ scanchain_147/module_data_out[0] scanchain_147/module_data_out[1] scanchain_147/module_data_out[2]
+ scanchain_147/module_data_out[3] scanchain_147/module_data_out[4] scanchain_147/module_data_out[5]
+ scanchain_147/module_data_out[6] scanchain_147/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_158 scanchain_158/module_data_in[0] scanchain_158/module_data_in[1]
+ scanchain_158/module_data_in[2] scanchain_158/module_data_in[3] scanchain_158/module_data_in[4]
+ scanchain_158/module_data_in[5] scanchain_158/module_data_in[6] scanchain_158/module_data_in[7]
+ scanchain_158/module_data_out[0] scanchain_158/module_data_out[1] scanchain_158/module_data_out[2]
+ scanchain_158/module_data_out[3] scanchain_158/module_data_out[4] scanchain_158/module_data_out[5]
+ scanchain_158/module_data_out[6] scanchain_158/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_169 scanchain_169/module_data_in[0] scanchain_169/module_data_in[1]
+ scanchain_169/module_data_in[2] scanchain_169/module_data_in[3] scanchain_169/module_data_in[4]
+ scanchain_169/module_data_in[5] scanchain_169/module_data_in[6] scanchain_169/module_data_in[7]
+ scanchain_169/module_data_out[0] scanchain_169/module_data_out[1] scanchain_169/module_data_out[2]
+ scanchain_169/module_data_out[3] scanchain_169/module_data_out[4] scanchain_169/module_data_out[5]
+ scanchain_169/module_data_out[6] scanchain_169/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_198 scanchain_198/clk_in scanchain_199/clk_in scanchain_198/data_in scanchain_199/data_in
+ scanchain_198/latch_enable_in scanchain_199/latch_enable_in scanchain_198/module_data_in[0]
+ scanchain_198/module_data_in[1] scanchain_198/module_data_in[2] scanchain_198/module_data_in[3]
+ scanchain_198/module_data_in[4] scanchain_198/module_data_in[5] scanchain_198/module_data_in[6]
+ scanchain_198/module_data_in[7] scanchain_198/module_data_out[0] scanchain_198/module_data_out[1]
+ scanchain_198/module_data_out[2] scanchain_198/module_data_out[3] scanchain_198/module_data_out[4]
+ scanchain_198/module_data_out[5] scanchain_198/module_data_out[6] scanchain_198/module_data_out[7]
+ scanchain_198/scan_select_in scanchain_199/scan_select_in vccd1 vssd1 scanchain
Xscanchain_110 scanchain_110/clk_in scanchain_111/clk_in scanchain_110/data_in scanchain_111/data_in
+ scanchain_110/latch_enable_in scanchain_111/latch_enable_in scanchain_110/module_data_in[0]
+ scanchain_110/module_data_in[1] scanchain_110/module_data_in[2] scanchain_110/module_data_in[3]
+ scanchain_110/module_data_in[4] scanchain_110/module_data_in[5] scanchain_110/module_data_in[6]
+ scanchain_110/module_data_in[7] scanchain_110/module_data_out[0] scanchain_110/module_data_out[1]
+ scanchain_110/module_data_out[2] scanchain_110/module_data_out[3] scanchain_110/module_data_out[4]
+ scanchain_110/module_data_out[5] scanchain_110/module_data_out[6] scanchain_110/module_data_out[7]
+ scanchain_110/scan_select_in scanchain_111/scan_select_in vccd1 vssd1 scanchain
Xscanchain_121 scanchain_121/clk_in scanchain_122/clk_in scanchain_121/data_in scanchain_122/data_in
+ scanchain_121/latch_enable_in scanchain_122/latch_enable_in scanchain_121/module_data_in[0]
+ scanchain_121/module_data_in[1] scanchain_121/module_data_in[2] scanchain_121/module_data_in[3]
+ scanchain_121/module_data_in[4] scanchain_121/module_data_in[5] scanchain_121/module_data_in[6]
+ scanchain_121/module_data_in[7] scanchain_121/module_data_out[0] scanchain_121/module_data_out[1]
+ scanchain_121/module_data_out[2] scanchain_121/module_data_out[3] scanchain_121/module_data_out[4]
+ scanchain_121/module_data_out[5] scanchain_121/module_data_out[6] scanchain_121/module_data_out[7]
+ scanchain_121/scan_select_in scanchain_122/scan_select_in vccd1 vssd1 scanchain
Xscanchain_132 scanchain_132/clk_in scanchain_133/clk_in scanchain_132/data_in scanchain_133/data_in
+ scanchain_132/latch_enable_in scanchain_133/latch_enable_in scanchain_132/module_data_in[0]
+ scanchain_132/module_data_in[1] scanchain_132/module_data_in[2] scanchain_132/module_data_in[3]
+ scanchain_132/module_data_in[4] scanchain_132/module_data_in[5] scanchain_132/module_data_in[6]
+ scanchain_132/module_data_in[7] scanchain_132/module_data_out[0] scanchain_132/module_data_out[1]
+ scanchain_132/module_data_out[2] scanchain_132/module_data_out[3] scanchain_132/module_data_out[4]
+ scanchain_132/module_data_out[5] scanchain_132/module_data_out[6] scanchain_132/module_data_out[7]
+ scanchain_132/scan_select_in scanchain_133/scan_select_in vccd1 vssd1 scanchain
Xscanchain_143 scanchain_143/clk_in scanchain_144/clk_in scanchain_143/data_in scanchain_144/data_in
+ scanchain_143/latch_enable_in scanchain_144/latch_enable_in scanchain_143/module_data_in[0]
+ scanchain_143/module_data_in[1] scanchain_143/module_data_in[2] scanchain_143/module_data_in[3]
+ scanchain_143/module_data_in[4] scanchain_143/module_data_in[5] scanchain_143/module_data_in[6]
+ scanchain_143/module_data_in[7] scanchain_143/module_data_out[0] scanchain_143/module_data_out[1]
+ scanchain_143/module_data_out[2] scanchain_143/module_data_out[3] scanchain_143/module_data_out[4]
+ scanchain_143/module_data_out[5] scanchain_143/module_data_out[6] scanchain_143/module_data_out[7]
+ scanchain_143/scan_select_in scanchain_144/scan_select_in vccd1 vssd1 scanchain
Xscanchain_165 scanchain_165/clk_in scanchain_166/clk_in scanchain_165/data_in scanchain_166/data_in
+ scanchain_165/latch_enable_in scanchain_166/latch_enable_in scanchain_165/module_data_in[0]
+ scanchain_165/module_data_in[1] scanchain_165/module_data_in[2] scanchain_165/module_data_in[3]
+ scanchain_165/module_data_in[4] scanchain_165/module_data_in[5] scanchain_165/module_data_in[6]
+ scanchain_165/module_data_in[7] scanchain_165/module_data_out[0] scanchain_165/module_data_out[1]
+ scanchain_165/module_data_out[2] scanchain_165/module_data_out[3] scanchain_165/module_data_out[4]
+ scanchain_165/module_data_out[5] scanchain_165/module_data_out[6] scanchain_165/module_data_out[7]
+ scanchain_165/scan_select_in scanchain_166/scan_select_in vccd1 vssd1 scanchain
Xscanchain_154 scanchain_154/clk_in scanchain_155/clk_in scanchain_154/data_in scanchain_155/data_in
+ scanchain_154/latch_enable_in scanchain_155/latch_enable_in scanchain_154/module_data_in[0]
+ scanchain_154/module_data_in[1] scanchain_154/module_data_in[2] scanchain_154/module_data_in[3]
+ scanchain_154/module_data_in[4] scanchain_154/module_data_in[5] scanchain_154/module_data_in[6]
+ scanchain_154/module_data_in[7] scanchain_154/module_data_out[0] scanchain_154/module_data_out[1]
+ scanchain_154/module_data_out[2] scanchain_154/module_data_out[3] scanchain_154/module_data_out[4]
+ scanchain_154/module_data_out[5] scanchain_154/module_data_out[6] scanchain_154/module_data_out[7]
+ scanchain_154/scan_select_in scanchain_155/scan_select_in vccd1 vssd1 scanchain
Xscanchain_176 scanchain_176/clk_in scanchain_177/clk_in scanchain_176/data_in scanchain_177/data_in
+ scanchain_176/latch_enable_in scanchain_177/latch_enable_in scanchain_176/module_data_in[0]
+ scanchain_176/module_data_in[1] scanchain_176/module_data_in[2] scanchain_176/module_data_in[3]
+ scanchain_176/module_data_in[4] scanchain_176/module_data_in[5] scanchain_176/module_data_in[6]
+ scanchain_176/module_data_in[7] scanchain_176/module_data_out[0] scanchain_176/module_data_out[1]
+ scanchain_176/module_data_out[2] scanchain_176/module_data_out[3] scanchain_176/module_data_out[4]
+ scanchain_176/module_data_out[5] scanchain_176/module_data_out[6] scanchain_176/module_data_out[7]
+ scanchain_176/scan_select_in scanchain_177/scan_select_in vccd1 vssd1 scanchain
Xscanchain_187 scanchain_187/clk_in scanchain_188/clk_in scanchain_187/data_in scanchain_188/data_in
+ scanchain_187/latch_enable_in scanchain_188/latch_enable_in scanchain_187/module_data_in[0]
+ scanchain_187/module_data_in[1] scanchain_187/module_data_in[2] scanchain_187/module_data_in[3]
+ scanchain_187/module_data_in[4] scanchain_187/module_data_in[5] scanchain_187/module_data_in[6]
+ scanchain_187/module_data_in[7] scanchain_187/module_data_out[0] scanchain_187/module_data_out[1]
+ scanchain_187/module_data_out[2] scanchain_187/module_data_out[3] scanchain_187/module_data_out[4]
+ scanchain_187/module_data_out[5] scanchain_187/module_data_out[6] scanchain_187/module_data_out[7]
+ scanchain_187/scan_select_in scanchain_188/scan_select_in vccd1 vssd1 scanchain
Xjar_illegal_logic_036 jar_illegal_logic_036/io_in[0] jar_illegal_logic_036/io_in[1]
+ jar_illegal_logic_036/io_in[2] jar_illegal_logic_036/io_in[3] jar_illegal_logic_036/io_in[4]
+ jar_illegal_logic_036/io_in[5] jar_illegal_logic_036/io_in[6] jar_illegal_logic_036/io_in[7]
+ jar_illegal_logic_036/io_out[0] jar_illegal_logic_036/io_out[1] jar_illegal_logic_036/io_out[2]
+ jar_illegal_logic_036/io_out[3] jar_illegal_logic_036/io_out[4] jar_illegal_logic_036/io_out[5]
+ jar_illegal_logic_036/io_out[6] jar_illegal_logic_036/io_out[7] vccd1 vssd1 jar_illegal_logic
Xmeriac_tt02_play_tune_045 scanchain_045/module_data_in[0] scanchain_045/module_data_in[1]
+ scanchain_045/module_data_in[2] scanchain_045/module_data_in[3] scanchain_045/module_data_in[4]
+ scanchain_045/module_data_in[5] scanchain_045/module_data_in[6] scanchain_045/module_data_in[7]
+ scanchain_045/module_data_out[0] scanchain_045/module_data_out[1] scanchain_045/module_data_out[2]
+ scanchain_045/module_data_out[3] scanchain_045/module_data_out[4] scanchain_045/module_data_out[5]
+ scanchain_045/module_data_out[6] scanchain_045/module_data_out[7] vccd1 vssd1 meriac_tt02_play_tune
Xuser_module_341535056611770964_104 scanchain_104/module_data_in[0] scanchain_104/module_data_in[1]
+ scanchain_104/module_data_in[2] scanchain_104/module_data_in[3] scanchain_104/module_data_in[4]
+ scanchain_104/module_data_in[5] scanchain_104/module_data_in[6] scanchain_104/module_data_in[7]
+ scanchain_104/module_data_out[0] scanchain_104/module_data_out[1] scanchain_104/module_data_out[2]
+ scanchain_104/module_data_out[3] scanchain_104/module_data_out[4] scanchain_104/module_data_out[5]
+ scanchain_104/module_data_out[6] scanchain_104/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_115 scanchain_115/module_data_in[0] scanchain_115/module_data_in[1]
+ scanchain_115/module_data_in[2] scanchain_115/module_data_in[3] scanchain_115/module_data_in[4]
+ scanchain_115/module_data_in[5] scanchain_115/module_data_in[6] scanchain_115/module_data_in[7]
+ scanchain_115/module_data_out[0] scanchain_115/module_data_out[1] scanchain_115/module_data_out[2]
+ scanchain_115/module_data_out[3] scanchain_115/module_data_out[4] scanchain_115/module_data_out[5]
+ scanchain_115/module_data_out[6] scanchain_115/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_137 scanchain_137/module_data_in[0] scanchain_137/module_data_in[1]
+ scanchain_137/module_data_in[2] scanchain_137/module_data_in[3] scanchain_137/module_data_in[4]
+ scanchain_137/module_data_in[5] scanchain_137/module_data_in[6] scanchain_137/module_data_in[7]
+ scanchain_137/module_data_out[0] scanchain_137/module_data_out[1] scanchain_137/module_data_out[2]
+ scanchain_137/module_data_out[3] scanchain_137/module_data_out[4] scanchain_137/module_data_out[5]
+ scanchain_137/module_data_out[6] scanchain_137/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_126 scanchain_126/module_data_in[0] scanchain_126/module_data_in[1]
+ scanchain_126/module_data_in[2] scanchain_126/module_data_in[3] scanchain_126/module_data_in[4]
+ scanchain_126/module_data_in[5] scanchain_126/module_data_in[6] scanchain_126/module_data_in[7]
+ scanchain_126/module_data_out[0] scanchain_126/module_data_out[1] scanchain_126/module_data_out[2]
+ scanchain_126/module_data_out[3] scanchain_126/module_data_out[4] scanchain_126/module_data_out[5]
+ scanchain_126/module_data_out[6] scanchain_126/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_148 scanchain_148/module_data_in[0] scanchain_148/module_data_in[1]
+ scanchain_148/module_data_in[2] scanchain_148/module_data_in[3] scanchain_148/module_data_in[4]
+ scanchain_148/module_data_in[5] scanchain_148/module_data_in[6] scanchain_148/module_data_in[7]
+ scanchain_148/module_data_out[0] scanchain_148/module_data_out[1] scanchain_148/module_data_out[2]
+ scanchain_148/module_data_out[3] scanchain_148/module_data_out[4] scanchain_148/module_data_out[5]
+ scanchain_148/module_data_out[6] scanchain_148/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_159 scanchain_159/module_data_in[0] scanchain_159/module_data_in[1]
+ scanchain_159/module_data_in[2] scanchain_159/module_data_in[3] scanchain_159/module_data_in[4]
+ scanchain_159/module_data_in[5] scanchain_159/module_data_in[6] scanchain_159/module_data_in[7]
+ scanchain_159/module_data_out[0] scanchain_159/module_data_out[1] scanchain_159/module_data_out[2]
+ scanchain_159/module_data_out[3] scanchain_159/module_data_out[4] scanchain_159/module_data_out[5]
+ scanchain_159/module_data_out[6] scanchain_159/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341178154799333971_085 scanchain_085/module_data_in[0] scanchain_085/module_data_in[1]
+ scanchain_085/module_data_in[2] scanchain_085/module_data_in[3] scanchain_085/module_data_in[4]
+ scanchain_085/module_data_in[5] scanchain_085/module_data_in[6] scanchain_085/module_data_in[7]
+ scanchain_085/module_data_out[0] scanchain_085/module_data_out[1] scanchain_085/module_data_out[2]
+ scanchain_085/module_data_out[3] scanchain_085/module_data_out[4] scanchain_085/module_data_out[5]
+ scanchain_085/module_data_out[6] scanchain_085/module_data_out[7] vccd1 vssd1 user_module_341178154799333971
Xtt2_tholin_namebadge_055 scanchain_055/module_data_in[0] scanchain_055/module_data_in[1]
+ scanchain_055/module_data_in[2] scanchain_055/module_data_in[3] scanchain_055/module_data_in[4]
+ scanchain_055/module_data_in[5] scanchain_055/module_data_in[6] scanchain_055/module_data_in[7]
+ scanchain_055/module_data_out[0] scanchain_055/module_data_out[1] scanchain_055/module_data_out[2]
+ scanchain_055/module_data_out[3] scanchain_055/module_data_out[4] scanchain_055/module_data_out[5]
+ scanchain_055/module_data_out[6] scanchain_055/module_data_out[7] vccd1 vssd1 tt2_tholin_namebadge
Xscanchain_100 scanchain_100/clk_in scanchain_101/clk_in scanchain_100/data_in scanchain_101/data_in
+ scanchain_100/latch_enable_in scanchain_101/latch_enable_in scanchain_100/module_data_in[0]
+ scanchain_100/module_data_in[1] scanchain_100/module_data_in[2] scanchain_100/module_data_in[3]
+ scanchain_100/module_data_in[4] scanchain_100/module_data_in[5] scanchain_100/module_data_in[6]
+ scanchain_100/module_data_in[7] scanchain_100/module_data_out[0] scanchain_100/module_data_out[1]
+ scanchain_100/module_data_out[2] scanchain_100/module_data_out[3] scanchain_100/module_data_out[4]
+ scanchain_100/module_data_out[5] scanchain_100/module_data_out[6] scanchain_100/module_data_out[7]
+ scanchain_100/scan_select_in scanchain_101/scan_select_in vccd1 vssd1 scanchain
Xscanchain_111 scanchain_111/clk_in scanchain_112/clk_in scanchain_111/data_in scanchain_112/data_in
+ scanchain_111/latch_enable_in scanchain_112/latch_enable_in scanchain_111/module_data_in[0]
+ scanchain_111/module_data_in[1] scanchain_111/module_data_in[2] scanchain_111/module_data_in[3]
+ scanchain_111/module_data_in[4] scanchain_111/module_data_in[5] scanchain_111/module_data_in[6]
+ scanchain_111/module_data_in[7] scanchain_111/module_data_out[0] scanchain_111/module_data_out[1]
+ scanchain_111/module_data_out[2] scanchain_111/module_data_out[3] scanchain_111/module_data_out[4]
+ scanchain_111/module_data_out[5] scanchain_111/module_data_out[6] scanchain_111/module_data_out[7]
+ scanchain_111/scan_select_in scanchain_112/scan_select_in vccd1 vssd1 scanchain
Xscanchain_122 scanchain_122/clk_in scanchain_123/clk_in scanchain_122/data_in scanchain_123/data_in
+ scanchain_122/latch_enable_in scanchain_123/latch_enable_in scanchain_122/module_data_in[0]
+ scanchain_122/module_data_in[1] scanchain_122/module_data_in[2] scanchain_122/module_data_in[3]
+ scanchain_122/module_data_in[4] scanchain_122/module_data_in[5] scanchain_122/module_data_in[6]
+ scanchain_122/module_data_in[7] scanchain_122/module_data_out[0] scanchain_122/module_data_out[1]
+ scanchain_122/module_data_out[2] scanchain_122/module_data_out[3] scanchain_122/module_data_out[4]
+ scanchain_122/module_data_out[5] scanchain_122/module_data_out[6] scanchain_122/module_data_out[7]
+ scanchain_122/scan_select_in scanchain_123/scan_select_in vccd1 vssd1 scanchain
Xscanchain_133 scanchain_133/clk_in scanchain_134/clk_in scanchain_133/data_in scanchain_134/data_in
+ scanchain_133/latch_enable_in scanchain_134/latch_enable_in scanchain_133/module_data_in[0]
+ scanchain_133/module_data_in[1] scanchain_133/module_data_in[2] scanchain_133/module_data_in[3]
+ scanchain_133/module_data_in[4] scanchain_133/module_data_in[5] scanchain_133/module_data_in[6]
+ scanchain_133/module_data_in[7] scanchain_133/module_data_out[0] scanchain_133/module_data_out[1]
+ scanchain_133/module_data_out[2] scanchain_133/module_data_out[3] scanchain_133/module_data_out[4]
+ scanchain_133/module_data_out[5] scanchain_133/module_data_out[6] scanchain_133/module_data_out[7]
+ scanchain_133/scan_select_in scanchain_134/scan_select_in vccd1 vssd1 scanchain
Xscanchain_144 scanchain_144/clk_in scanchain_145/clk_in scanchain_144/data_in scanchain_145/data_in
+ scanchain_144/latch_enable_in scanchain_145/latch_enable_in scanchain_144/module_data_in[0]
+ scanchain_144/module_data_in[1] scanchain_144/module_data_in[2] scanchain_144/module_data_in[3]
+ scanchain_144/module_data_in[4] scanchain_144/module_data_in[5] scanchain_144/module_data_in[6]
+ scanchain_144/module_data_in[7] scanchain_144/module_data_out[0] scanchain_144/module_data_out[1]
+ scanchain_144/module_data_out[2] scanchain_144/module_data_out[3] scanchain_144/module_data_out[4]
+ scanchain_144/module_data_out[5] scanchain_144/module_data_out[6] scanchain_144/module_data_out[7]
+ scanchain_144/scan_select_in scanchain_145/scan_select_in vccd1 vssd1 scanchain
Xscanchain_155 scanchain_155/clk_in scanchain_156/clk_in scanchain_155/data_in scanchain_156/data_in
+ scanchain_155/latch_enable_in scanchain_156/latch_enable_in scanchain_155/module_data_in[0]
+ scanchain_155/module_data_in[1] scanchain_155/module_data_in[2] scanchain_155/module_data_in[3]
+ scanchain_155/module_data_in[4] scanchain_155/module_data_in[5] scanchain_155/module_data_in[6]
+ scanchain_155/module_data_in[7] scanchain_155/module_data_out[0] scanchain_155/module_data_out[1]
+ scanchain_155/module_data_out[2] scanchain_155/module_data_out[3] scanchain_155/module_data_out[4]
+ scanchain_155/module_data_out[5] scanchain_155/module_data_out[6] scanchain_155/module_data_out[7]
+ scanchain_155/scan_select_in scanchain_156/scan_select_in vccd1 vssd1 scanchain
Xscanchain_166 scanchain_166/clk_in scanchain_167/clk_in scanchain_166/data_in scanchain_167/data_in
+ scanchain_166/latch_enable_in scanchain_167/latch_enable_in scanchain_166/module_data_in[0]
+ scanchain_166/module_data_in[1] scanchain_166/module_data_in[2] scanchain_166/module_data_in[3]
+ scanchain_166/module_data_in[4] scanchain_166/module_data_in[5] scanchain_166/module_data_in[6]
+ scanchain_166/module_data_in[7] scanchain_166/module_data_out[0] scanchain_166/module_data_out[1]
+ scanchain_166/module_data_out[2] scanchain_166/module_data_out[3] scanchain_166/module_data_out[4]
+ scanchain_166/module_data_out[5] scanchain_166/module_data_out[6] scanchain_166/module_data_out[7]
+ scanchain_166/scan_select_in scanchain_167/scan_select_in vccd1 vssd1 scanchain
Xscanchain_199 scanchain_199/clk_in scanchain_200/clk_in scanchain_199/data_in scanchain_200/data_in
+ scanchain_199/latch_enable_in scanchain_200/latch_enable_in scanchain_199/module_data_in[0]
+ scanchain_199/module_data_in[1] scanchain_199/module_data_in[2] scanchain_199/module_data_in[3]
+ scanchain_199/module_data_in[4] scanchain_199/module_data_in[5] scanchain_199/module_data_in[6]
+ scanchain_199/module_data_in[7] scanchain_199/module_data_out[0] scanchain_199/module_data_out[1]
+ scanchain_199/module_data_out[2] scanchain_199/module_data_out[3] scanchain_199/module_data_out[4]
+ scanchain_199/module_data_out[5] scanchain_199/module_data_out[6] scanchain_199/module_data_out[7]
+ scanchain_199/scan_select_in scanchain_200/scan_select_in vccd1 vssd1 scanchain
Xscanchain_177 scanchain_177/clk_in scanchain_178/clk_in scanchain_177/data_in scanchain_178/data_in
+ scanchain_177/latch_enable_in scanchain_178/latch_enable_in scanchain_177/module_data_in[0]
+ scanchain_177/module_data_in[1] scanchain_177/module_data_in[2] scanchain_177/module_data_in[3]
+ scanchain_177/module_data_in[4] scanchain_177/module_data_in[5] scanchain_177/module_data_in[6]
+ scanchain_177/module_data_in[7] scanchain_177/module_data_out[0] scanchain_177/module_data_out[1]
+ scanchain_177/module_data_out[2] scanchain_177/module_data_out[3] scanchain_177/module_data_out[4]
+ scanchain_177/module_data_out[5] scanchain_177/module_data_out[6] scanchain_177/module_data_out[7]
+ scanchain_177/scan_select_in scanchain_178/scan_select_in vccd1 vssd1 scanchain
Xscanchain_188 scanchain_188/clk_in scanchain_189/clk_in scanchain_188/data_in scanchain_189/data_in
+ scanchain_188/latch_enable_in scanchain_189/latch_enable_in scanchain_188/module_data_in[0]
+ scanchain_188/module_data_in[1] scanchain_188/module_data_in[2] scanchain_188/module_data_in[3]
+ scanchain_188/module_data_in[4] scanchain_188/module_data_in[5] scanchain_188/module_data_in[6]
+ scanchain_188/module_data_in[7] scanchain_188/module_data_out[0] scanchain_188/module_data_out[1]
+ scanchain_188/module_data_out[2] scanchain_188/module_data_out[3] scanchain_188/module_data_out[4]
+ scanchain_188/module_data_out[5] scanchain_188/module_data_out[6] scanchain_188/module_data_out[7]
+ scanchain_188/scan_select_in scanchain_189/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341490465660469844_064 scanchain_064/module_data_in[0] scanchain_064/module_data_in[1]
+ scanchain_064/module_data_in[2] scanchain_064/module_data_in[3] scanchain_064/module_data_in[4]
+ scanchain_064/module_data_in[5] scanchain_064/module_data_in[6] scanchain_064/module_data_in[7]
+ scanchain_064/module_data_out[0] scanchain_064/module_data_out[1] scanchain_064/module_data_out[2]
+ scanchain_064/module_data_out[3] scanchain_064/module_data_out[4] scanchain_064/module_data_out[5]
+ scanchain_064/module_data_out[6] scanchain_064/module_data_out[7] vccd1 vssd1 user_module_341490465660469844
Xuser_module_341608574336631379_091 scanchain_091/module_data_in[0] scanchain_091/module_data_in[1]
+ scanchain_091/module_data_in[2] scanchain_091/module_data_in[3] scanchain_091/module_data_in[4]
+ scanchain_091/module_data_in[5] scanchain_091/module_data_in[6] scanchain_091/module_data_in[7]
+ scanchain_091/module_data_out[0] scanchain_091/module_data_out[1] scanchain_091/module_data_out[2]
+ scanchain_091/module_data_out[3] scanchain_091/module_data_out[4] scanchain_091/module_data_out[5]
+ scanchain_091/module_data_out[6] scanchain_091/module_data_out[7] vccd1 vssd1 user_module_341608574336631379
Xkrasin_3_bit_8_channel_pwm_driver_057 scanchain_057/module_data_in[0] scanchain_057/module_data_in[1]
+ scanchain_057/module_data_in[2] scanchain_057/module_data_in[3] scanchain_057/module_data_in[4]
+ scanchain_057/module_data_in[5] scanchain_057/module_data_in[6] scanchain_057/module_data_in[7]
+ scanchain_057/module_data_out[0] scanchain_057/module_data_out[1] scanchain_057/module_data_out[2]
+ scanchain_057/module_data_out[3] scanchain_057/module_data_out[4] scanchain_057/module_data_out[5]
+ scanchain_057/module_data_out[6] scanchain_057/module_data_out[7] vccd1 vssd1 krasin_3_bit_8_channel_pwm_driver
Xuser_module_341535056611770964_105 scanchain_105/module_data_in[0] scanchain_105/module_data_in[1]
+ scanchain_105/module_data_in[2] scanchain_105/module_data_in[3] scanchain_105/module_data_in[4]
+ scanchain_105/module_data_in[5] scanchain_105/module_data_in[6] scanchain_105/module_data_in[7]
+ scanchain_105/module_data_out[0] scanchain_105/module_data_out[1] scanchain_105/module_data_out[2]
+ scanchain_105/module_data_out[3] scanchain_105/module_data_out[4] scanchain_105/module_data_out[5]
+ scanchain_105/module_data_out[6] scanchain_105/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_116 scanchain_116/module_data_in[0] scanchain_116/module_data_in[1]
+ scanchain_116/module_data_in[2] scanchain_116/module_data_in[3] scanchain_116/module_data_in[4]
+ scanchain_116/module_data_in[5] scanchain_116/module_data_in[6] scanchain_116/module_data_in[7]
+ scanchain_116/module_data_out[0] scanchain_116/module_data_out[1] scanchain_116/module_data_out[2]
+ scanchain_116/module_data_out[3] scanchain_116/module_data_out[4] scanchain_116/module_data_out[5]
+ scanchain_116/module_data_out[6] scanchain_116/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_127 scanchain_127/module_data_in[0] scanchain_127/module_data_in[1]
+ scanchain_127/module_data_in[2] scanchain_127/module_data_in[3] scanchain_127/module_data_in[4]
+ scanchain_127/module_data_in[5] scanchain_127/module_data_in[6] scanchain_127/module_data_in[7]
+ scanchain_127/module_data_out[0] scanchain_127/module_data_out[1] scanchain_127/module_data_out[2]
+ scanchain_127/module_data_out[3] scanchain_127/module_data_out[4] scanchain_127/module_data_out[5]
+ scanchain_127/module_data_out[6] scanchain_127/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_138 scanchain_138/module_data_in[0] scanchain_138/module_data_in[1]
+ scanchain_138/module_data_in[2] scanchain_138/module_data_in[3] scanchain_138/module_data_in[4]
+ scanchain_138/module_data_in[5] scanchain_138/module_data_in[6] scanchain_138/module_data_in[7]
+ scanchain_138/module_data_out[0] scanchain_138/module_data_out[1] scanchain_138/module_data_out[2]
+ scanchain_138/module_data_out[3] scanchain_138/module_data_out[4] scanchain_138/module_data_out[5]
+ scanchain_138/module_data_out[6] scanchain_138/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_149 scanchain_149/module_data_in[0] scanchain_149/module_data_in[1]
+ scanchain_149/module_data_in[2] scanchain_149/module_data_in[3] scanchain_149/module_data_in[4]
+ scanchain_149/module_data_in[5] scanchain_149/module_data_in[6] scanchain_149/module_data_in[7]
+ scanchain_149/module_data_out[0] scanchain_149/module_data_out[1] scanchain_149/module_data_out[2]
+ scanchain_149/module_data_out[3] scanchain_149/module_data_out[4] scanchain_149/module_data_out[5]
+ scanchain_149/module_data_out[6] scanchain_149/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xthunderbird_taillight_ctrl_088 scanchain_088/module_data_in[0] scanchain_088/module_data_in[1]
+ scanchain_088/module_data_in[2] scanchain_088/module_data_in[3] scanchain_088/module_data_in[4]
+ scanchain_088/module_data_in[5] scanchain_088/module_data_in[6] scanchain_088/module_data_in[7]
+ scanchain_088/module_data_out[0] scanchain_088/module_data_out[1] scanchain_088/module_data_out[2]
+ scanchain_088/module_data_out[3] scanchain_088/module_data_out[4] scanchain_088/module_data_out[5]
+ scanchain_088/module_data_out[6] scanchain_088/module_data_out[7] vccd1 vssd1 thunderbird_taillight_ctrl
Xmbikovitsky_top_033 mbikovitsky_top_033/io_in[0] mbikovitsky_top_033/io_in[1] mbikovitsky_top_033/io_in[2]
+ mbikovitsky_top_033/io_in[3] mbikovitsky_top_033/io_in[4] mbikovitsky_top_033/io_in[5]
+ mbikovitsky_top_033/io_in[6] mbikovitsky_top_033/io_in[7] mbikovitsky_top_033/io_out[0]
+ mbikovitsky_top_033/io_out[1] mbikovitsky_top_033/io_out[2] mbikovitsky_top_033/io_out[3]
+ mbikovitsky_top_033/io_out[4] mbikovitsky_top_033/io_out[5] mbikovitsky_top_033/io_out[6]
+ mbikovitsky_top_033/io_out[7] vccd1 vssd1 mbikovitsky_top
Xscanchain_101 scanchain_101/clk_in scanchain_102/clk_in scanchain_101/data_in scanchain_102/data_in
+ scanchain_101/latch_enable_in scanchain_102/latch_enable_in scanchain_101/module_data_in[0]
+ scanchain_101/module_data_in[1] scanchain_101/module_data_in[2] scanchain_101/module_data_in[3]
+ scanchain_101/module_data_in[4] scanchain_101/module_data_in[5] scanchain_101/module_data_in[6]
+ scanchain_101/module_data_in[7] scanchain_101/module_data_out[0] scanchain_101/module_data_out[1]
+ scanchain_101/module_data_out[2] scanchain_101/module_data_out[3] scanchain_101/module_data_out[4]
+ scanchain_101/module_data_out[5] scanchain_101/module_data_out[6] scanchain_101/module_data_out[7]
+ scanchain_101/scan_select_in scanchain_102/scan_select_in vccd1 vssd1 scanchain
Xscanchain_112 scanchain_112/clk_in scanchain_113/clk_in scanchain_112/data_in scanchain_113/data_in
+ scanchain_112/latch_enable_in scanchain_113/latch_enable_in scanchain_112/module_data_in[0]
+ scanchain_112/module_data_in[1] scanchain_112/module_data_in[2] scanchain_112/module_data_in[3]
+ scanchain_112/module_data_in[4] scanchain_112/module_data_in[5] scanchain_112/module_data_in[6]
+ scanchain_112/module_data_in[7] scanchain_112/module_data_out[0] scanchain_112/module_data_out[1]
+ scanchain_112/module_data_out[2] scanchain_112/module_data_out[3] scanchain_112/module_data_out[4]
+ scanchain_112/module_data_out[5] scanchain_112/module_data_out[6] scanchain_112/module_data_out[7]
+ scanchain_112/scan_select_in scanchain_113/scan_select_in vccd1 vssd1 scanchain
Xscanchain_123 scanchain_123/clk_in scanchain_124/clk_in scanchain_123/data_in scanchain_124/data_in
+ scanchain_123/latch_enable_in scanchain_124/latch_enable_in scanchain_123/module_data_in[0]
+ scanchain_123/module_data_in[1] scanchain_123/module_data_in[2] scanchain_123/module_data_in[3]
+ scanchain_123/module_data_in[4] scanchain_123/module_data_in[5] scanchain_123/module_data_in[6]
+ scanchain_123/module_data_in[7] scanchain_123/module_data_out[0] scanchain_123/module_data_out[1]
+ scanchain_123/module_data_out[2] scanchain_123/module_data_out[3] scanchain_123/module_data_out[4]
+ scanchain_123/module_data_out[5] scanchain_123/module_data_out[6] scanchain_123/module_data_out[7]
+ scanchain_123/scan_select_in scanchain_124/scan_select_in vccd1 vssd1 scanchain
Xscanchain_134 scanchain_134/clk_in scanchain_135/clk_in scanchain_134/data_in scanchain_135/data_in
+ scanchain_134/latch_enable_in scanchain_135/latch_enable_in scanchain_134/module_data_in[0]
+ scanchain_134/module_data_in[1] scanchain_134/module_data_in[2] scanchain_134/module_data_in[3]
+ scanchain_134/module_data_in[4] scanchain_134/module_data_in[5] scanchain_134/module_data_in[6]
+ scanchain_134/module_data_in[7] scanchain_134/module_data_out[0] scanchain_134/module_data_out[1]
+ scanchain_134/module_data_out[2] scanchain_134/module_data_out[3] scanchain_134/module_data_out[4]
+ scanchain_134/module_data_out[5] scanchain_134/module_data_out[6] scanchain_134/module_data_out[7]
+ scanchain_134/scan_select_in scanchain_135/scan_select_in vccd1 vssd1 scanchain
Xscanchain_145 scanchain_145/clk_in scanchain_146/clk_in scanchain_145/data_in scanchain_146/data_in
+ scanchain_145/latch_enable_in scanchain_146/latch_enable_in scanchain_145/module_data_in[0]
+ scanchain_145/module_data_in[1] scanchain_145/module_data_in[2] scanchain_145/module_data_in[3]
+ scanchain_145/module_data_in[4] scanchain_145/module_data_in[5] scanchain_145/module_data_in[6]
+ scanchain_145/module_data_in[7] scanchain_145/module_data_out[0] scanchain_145/module_data_out[1]
+ scanchain_145/module_data_out[2] scanchain_145/module_data_out[3] scanchain_145/module_data_out[4]
+ scanchain_145/module_data_out[5] scanchain_145/module_data_out[6] scanchain_145/module_data_out[7]
+ scanchain_145/scan_select_in scanchain_146/scan_select_in vccd1 vssd1 scanchain
Xscanchain_156 scanchain_156/clk_in scanchain_157/clk_in scanchain_156/data_in scanchain_157/data_in
+ scanchain_156/latch_enable_in scanchain_157/latch_enable_in scanchain_156/module_data_in[0]
+ scanchain_156/module_data_in[1] scanchain_156/module_data_in[2] scanchain_156/module_data_in[3]
+ scanchain_156/module_data_in[4] scanchain_156/module_data_in[5] scanchain_156/module_data_in[6]
+ scanchain_156/module_data_in[7] scanchain_156/module_data_out[0] scanchain_156/module_data_out[1]
+ scanchain_156/module_data_out[2] scanchain_156/module_data_out[3] scanchain_156/module_data_out[4]
+ scanchain_156/module_data_out[5] scanchain_156/module_data_out[6] scanchain_156/module_data_out[7]
+ scanchain_156/scan_select_in scanchain_157/scan_select_in vccd1 vssd1 scanchain
Xscanchain_167 scanchain_167/clk_in scanchain_168/clk_in scanchain_167/data_in scanchain_168/data_in
+ scanchain_167/latch_enable_in scanchain_168/latch_enable_in scanchain_167/module_data_in[0]
+ scanchain_167/module_data_in[1] scanchain_167/module_data_in[2] scanchain_167/module_data_in[3]
+ scanchain_167/module_data_in[4] scanchain_167/module_data_in[5] scanchain_167/module_data_in[6]
+ scanchain_167/module_data_in[7] scanchain_167/module_data_out[0] scanchain_167/module_data_out[1]
+ scanchain_167/module_data_out[2] scanchain_167/module_data_out[3] scanchain_167/module_data_out[4]
+ scanchain_167/module_data_out[5] scanchain_167/module_data_out[6] scanchain_167/module_data_out[7]
+ scanchain_167/scan_select_in scanchain_168/scan_select_in vccd1 vssd1 scanchain
Xscanchain_178 scanchain_178/clk_in scanchain_179/clk_in scanchain_178/data_in scanchain_179/data_in
+ scanchain_178/latch_enable_in scanchain_179/latch_enable_in scanchain_178/module_data_in[0]
+ scanchain_178/module_data_in[1] scanchain_178/module_data_in[2] scanchain_178/module_data_in[3]
+ scanchain_178/module_data_in[4] scanchain_178/module_data_in[5] scanchain_178/module_data_in[6]
+ scanchain_178/module_data_in[7] scanchain_178/module_data_out[0] scanchain_178/module_data_out[1]
+ scanchain_178/module_data_out[2] scanchain_178/module_data_out[3] scanchain_178/module_data_out[4]
+ scanchain_178/module_data_out[5] scanchain_178/module_data_out[6] scanchain_178/module_data_out[7]
+ scanchain_178/scan_select_in scanchain_179/scan_select_in vccd1 vssd1 scanchain
Xscanchain_189 scanchain_189/clk_in scanchain_190/clk_in scanchain_189/data_in scanchain_190/data_in
+ scanchain_189/latch_enable_in scanchain_190/latch_enable_in scanchain_189/module_data_in[0]
+ scanchain_189/module_data_in[1] scanchain_189/module_data_in[2] scanchain_189/module_data_in[3]
+ scanchain_189/module_data_in[4] scanchain_189/module_data_in[5] scanchain_189/module_data_in[6]
+ scanchain_189/module_data_in[7] scanchain_189/module_data_out[0] scanchain_189/module_data_out[1]
+ scanchain_189/module_data_out[2] scanchain_189/module_data_out[3] scanchain_189/module_data_out[4]
+ scanchain_189/module_data_out[5] scanchain_189/module_data_out[6] scanchain_189/module_data_out[7]
+ scanchain_189/scan_select_in scanchain_190/scan_select_in vccd1 vssd1 scanchain
Xuser_module_347592305412145748_013 scanchain_013/module_data_in[0] scanchain_013/module_data_in[1]
+ scanchain_013/module_data_in[2] scanchain_013/module_data_in[3] scanchain_013/module_data_in[4]
+ scanchain_013/module_data_in[5] scanchain_013/module_data_in[6] scanchain_013/module_data_in[7]
+ scanchain_013/module_data_out[0] scanchain_013/module_data_out[1] scanchain_013/module_data_out[2]
+ scanchain_013/module_data_out[3] scanchain_013/module_data_out[4] scanchain_013/module_data_out[5]
+ scanchain_013/module_data_out[6] scanchain_013/module_data_out[7] vccd1 vssd1 user_module_347592305412145748
Xmoyes0_top_module_039 moyes0_top_module_039/io_in[0] moyes0_top_module_039/io_in[1]
+ moyes0_top_module_039/io_in[2] moyes0_top_module_039/io_in[3] moyes0_top_module_039/io_in[4]
+ moyes0_top_module_039/io_in[5] moyes0_top_module_039/io_in[6] moyes0_top_module_039/io_in[7]
+ moyes0_top_module_039/io_out[0] moyes0_top_module_039/io_out[1] moyes0_top_module_039/io_out[2]
+ moyes0_top_module_039/io_out[3] moyes0_top_module_039/io_out[4] moyes0_top_module_039/io_out[5]
+ moyes0_top_module_039/io_out[6] moyes0_top_module_039/io_out[7] vccd1 vssd1 moyes0_top_module
Xuser_module_341535056611770964_106 scanchain_106/module_data_in[0] scanchain_106/module_data_in[1]
+ scanchain_106/module_data_in[2] scanchain_106/module_data_in[3] scanchain_106/module_data_in[4]
+ scanchain_106/module_data_in[5] scanchain_106/module_data_in[6] scanchain_106/module_data_in[7]
+ scanchain_106/module_data_out[0] scanchain_106/module_data_out[1] scanchain_106/module_data_out[2]
+ scanchain_106/module_data_out[3] scanchain_106/module_data_out[4] scanchain_106/module_data_out[5]
+ scanchain_106/module_data_out[6] scanchain_106/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_117 scanchain_117/module_data_in[0] scanchain_117/module_data_in[1]
+ scanchain_117/module_data_in[2] scanchain_117/module_data_in[3] scanchain_117/module_data_in[4]
+ scanchain_117/module_data_in[5] scanchain_117/module_data_in[6] scanchain_117/module_data_in[7]
+ scanchain_117/module_data_out[0] scanchain_117/module_data_out[1] scanchain_117/module_data_out[2]
+ scanchain_117/module_data_out[3] scanchain_117/module_data_out[4] scanchain_117/module_data_out[5]
+ scanchain_117/module_data_out[6] scanchain_117/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_128 scanchain_128/module_data_in[0] scanchain_128/module_data_in[1]
+ scanchain_128/module_data_in[2] scanchain_128/module_data_in[3] scanchain_128/module_data_in[4]
+ scanchain_128/module_data_in[5] scanchain_128/module_data_in[6] scanchain_128/module_data_in[7]
+ scanchain_128/module_data_out[0] scanchain_128/module_data_out[1] scanchain_128/module_data_out[2]
+ scanchain_128/module_data_out[3] scanchain_128/module_data_out[4] scanchain_128/module_data_out[5]
+ scanchain_128/module_data_out[6] scanchain_128/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_139 scanchain_139/module_data_in[0] scanchain_139/module_data_in[1]
+ scanchain_139/module_data_in[2] scanchain_139/module_data_in[3] scanchain_139/module_data_in[4]
+ scanchain_139/module_data_in[5] scanchain_139/module_data_in[6] scanchain_139/module_data_in[7]
+ scanchain_139/module_data_out[0] scanchain_139/module_data_out[1] scanchain_139/module_data_out[2]
+ scanchain_139/module_data_out[3] scanchain_139/module_data_out[4] scanchain_139/module_data_out[5]
+ scanchain_139/module_data_out[6] scanchain_139/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xcpldcpu_MCPU5plus_077 cpldcpu_MCPU5plus_077/io_in[0] cpldcpu_MCPU5plus_077/io_in[1]
+ cpldcpu_MCPU5plus_077/io_in[2] cpldcpu_MCPU5plus_077/io_in[3] cpldcpu_MCPU5plus_077/io_in[4]
+ cpldcpu_MCPU5plus_077/io_in[5] cpldcpu_MCPU5plus_077/io_in[6] cpldcpu_MCPU5plus_077/io_in[7]
+ cpldcpu_MCPU5plus_077/io_out[0] cpldcpu_MCPU5plus_077/io_out[1] cpldcpu_MCPU5plus_077/io_out[2]
+ cpldcpu_MCPU5plus_077/io_out[3] cpldcpu_MCPU5plus_077/io_out[4] cpldcpu_MCPU5plus_077/io_out[5]
+ cpldcpu_MCPU5plus_077/io_out[6] cpldcpu_MCPU5plus_077/io_out[7] vccd1 vssd1 cpldcpu_MCPU5plus
Xscanchain_102 scanchain_102/clk_in scanchain_103/clk_in scanchain_102/data_in scanchain_103/data_in
+ scanchain_102/latch_enable_in scanchain_103/latch_enable_in scanchain_102/module_data_in[0]
+ scanchain_102/module_data_in[1] scanchain_102/module_data_in[2] scanchain_102/module_data_in[3]
+ scanchain_102/module_data_in[4] scanchain_102/module_data_in[5] scanchain_102/module_data_in[6]
+ scanchain_102/module_data_in[7] scanchain_102/module_data_out[0] scanchain_102/module_data_out[1]
+ scanchain_102/module_data_out[2] scanchain_102/module_data_out[3] scanchain_102/module_data_out[4]
+ scanchain_102/module_data_out[5] scanchain_102/module_data_out[6] scanchain_102/module_data_out[7]
+ scanchain_102/scan_select_in scanchain_103/scan_select_in vccd1 vssd1 scanchain
Xscanchain_113 scanchain_113/clk_in scanchain_114/clk_in scanchain_113/data_in scanchain_114/data_in
+ scanchain_113/latch_enable_in scanchain_114/latch_enable_in scanchain_113/module_data_in[0]
+ scanchain_113/module_data_in[1] scanchain_113/module_data_in[2] scanchain_113/module_data_in[3]
+ scanchain_113/module_data_in[4] scanchain_113/module_data_in[5] scanchain_113/module_data_in[6]
+ scanchain_113/module_data_in[7] scanchain_113/module_data_out[0] scanchain_113/module_data_out[1]
+ scanchain_113/module_data_out[2] scanchain_113/module_data_out[3] scanchain_113/module_data_out[4]
+ scanchain_113/module_data_out[5] scanchain_113/module_data_out[6] scanchain_113/module_data_out[7]
+ scanchain_113/scan_select_in scanchain_114/scan_select_in vccd1 vssd1 scanchain
Xscanchain_135 scanchain_135/clk_in scanchain_136/clk_in scanchain_135/data_in scanchain_136/data_in
+ scanchain_135/latch_enable_in scanchain_136/latch_enable_in scanchain_135/module_data_in[0]
+ scanchain_135/module_data_in[1] scanchain_135/module_data_in[2] scanchain_135/module_data_in[3]
+ scanchain_135/module_data_in[4] scanchain_135/module_data_in[5] scanchain_135/module_data_in[6]
+ scanchain_135/module_data_in[7] scanchain_135/module_data_out[0] scanchain_135/module_data_out[1]
+ scanchain_135/module_data_out[2] scanchain_135/module_data_out[3] scanchain_135/module_data_out[4]
+ scanchain_135/module_data_out[5] scanchain_135/module_data_out[6] scanchain_135/module_data_out[7]
+ scanchain_135/scan_select_in scanchain_136/scan_select_in vccd1 vssd1 scanchain
Xscanchain_124 scanchain_124/clk_in scanchain_125/clk_in scanchain_124/data_in scanchain_125/data_in
+ scanchain_124/latch_enable_in scanchain_125/latch_enable_in scanchain_124/module_data_in[0]
+ scanchain_124/module_data_in[1] scanchain_124/module_data_in[2] scanchain_124/module_data_in[3]
+ scanchain_124/module_data_in[4] scanchain_124/module_data_in[5] scanchain_124/module_data_in[6]
+ scanchain_124/module_data_in[7] scanchain_124/module_data_out[0] scanchain_124/module_data_out[1]
+ scanchain_124/module_data_out[2] scanchain_124/module_data_out[3] scanchain_124/module_data_out[4]
+ scanchain_124/module_data_out[5] scanchain_124/module_data_out[6] scanchain_124/module_data_out[7]
+ scanchain_124/scan_select_in scanchain_125/scan_select_in vccd1 vssd1 scanchain
Xscanchain_146 scanchain_146/clk_in scanchain_147/clk_in scanchain_146/data_in scanchain_147/data_in
+ scanchain_146/latch_enable_in scanchain_147/latch_enable_in scanchain_146/module_data_in[0]
+ scanchain_146/module_data_in[1] scanchain_146/module_data_in[2] scanchain_146/module_data_in[3]
+ scanchain_146/module_data_in[4] scanchain_146/module_data_in[5] scanchain_146/module_data_in[6]
+ scanchain_146/module_data_in[7] scanchain_146/module_data_out[0] scanchain_146/module_data_out[1]
+ scanchain_146/module_data_out[2] scanchain_146/module_data_out[3] scanchain_146/module_data_out[4]
+ scanchain_146/module_data_out[5] scanchain_146/module_data_out[6] scanchain_146/module_data_out[7]
+ scanchain_146/scan_select_in scanchain_147/scan_select_in vccd1 vssd1 scanchain
Xscanchain_157 scanchain_157/clk_in scanchain_158/clk_in scanchain_157/data_in scanchain_158/data_in
+ scanchain_157/latch_enable_in scanchain_158/latch_enable_in scanchain_157/module_data_in[0]
+ scanchain_157/module_data_in[1] scanchain_157/module_data_in[2] scanchain_157/module_data_in[3]
+ scanchain_157/module_data_in[4] scanchain_157/module_data_in[5] scanchain_157/module_data_in[6]
+ scanchain_157/module_data_in[7] scanchain_157/module_data_out[0] scanchain_157/module_data_out[1]
+ scanchain_157/module_data_out[2] scanchain_157/module_data_out[3] scanchain_157/module_data_out[4]
+ scanchain_157/module_data_out[5] scanchain_157/module_data_out[6] scanchain_157/module_data_out[7]
+ scanchain_157/scan_select_in scanchain_158/scan_select_in vccd1 vssd1 scanchain
Xscanchain_168 scanchain_168/clk_in scanchain_169/clk_in scanchain_168/data_in scanchain_169/data_in
+ scanchain_168/latch_enable_in scanchain_169/latch_enable_in scanchain_168/module_data_in[0]
+ scanchain_168/module_data_in[1] scanchain_168/module_data_in[2] scanchain_168/module_data_in[3]
+ scanchain_168/module_data_in[4] scanchain_168/module_data_in[5] scanchain_168/module_data_in[6]
+ scanchain_168/module_data_in[7] scanchain_168/module_data_out[0] scanchain_168/module_data_out[1]
+ scanchain_168/module_data_out[2] scanchain_168/module_data_out[3] scanchain_168/module_data_out[4]
+ scanchain_168/module_data_out[5] scanchain_168/module_data_out[6] scanchain_168/module_data_out[7]
+ scanchain_168/scan_select_in scanchain_169/scan_select_in vccd1 vssd1 scanchain
Xscanchain_179 scanchain_179/clk_in scanchain_180/clk_in scanchain_179/data_in scanchain_180/data_in
+ scanchain_179/latch_enable_in scanchain_180/latch_enable_in scanchain_179/module_data_in[0]
+ scanchain_179/module_data_in[1] scanchain_179/module_data_in[2] scanchain_179/module_data_in[3]
+ scanchain_179/module_data_in[4] scanchain_179/module_data_in[5] scanchain_179/module_data_in[6]
+ scanchain_179/module_data_in[7] scanchain_179/module_data_out[0] scanchain_179/module_data_out[1]
+ scanchain_179/module_data_out[2] scanchain_179/module_data_out[3] scanchain_179/module_data_out[4]
+ scanchain_179/module_data_out[5] scanchain_179/module_data_out[6] scanchain_179/module_data_out[7]
+ scanchain_179/scan_select_in scanchain_180/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_107 scanchain_107/module_data_in[0] scanchain_107/module_data_in[1]
+ scanchain_107/module_data_in[2] scanchain_107/module_data_in[3] scanchain_107/module_data_in[4]
+ scanchain_107/module_data_in[5] scanchain_107/module_data_in[6] scanchain_107/module_data_in[7]
+ scanchain_107/module_data_out[0] scanchain_107/module_data_out[1] scanchain_107/module_data_out[2]
+ scanchain_107/module_data_out[3] scanchain_107/module_data_out[4] scanchain_107/module_data_out[5]
+ scanchain_107/module_data_out[6] scanchain_107/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_118 scanchain_118/module_data_in[0] scanchain_118/module_data_in[1]
+ scanchain_118/module_data_in[2] scanchain_118/module_data_in[3] scanchain_118/module_data_in[4]
+ scanchain_118/module_data_in[5] scanchain_118/module_data_in[6] scanchain_118/module_data_in[7]
+ scanchain_118/module_data_out[0] scanchain_118/module_data_out[1] scanchain_118/module_data_out[2]
+ scanchain_118/module_data_out[3] scanchain_118/module_data_out[4] scanchain_118/module_data_out[5]
+ scanchain_118/module_data_out[6] scanchain_118/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_129 scanchain_129/module_data_in[0] scanchain_129/module_data_in[1]
+ scanchain_129/module_data_in[2] scanchain_129/module_data_in[3] scanchain_129/module_data_in[4]
+ scanchain_129/module_data_in[5] scanchain_129/module_data_in[6] scanchain_129/module_data_in[7]
+ scanchain_129/module_data_out[0] scanchain_129/module_data_out[1] scanchain_129/module_data_out[2]
+ scanchain_129/module_data_out[3] scanchain_129/module_data_out[4] scanchain_129/module_data_out[5]
+ scanchain_129/module_data_out[6] scanchain_129/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_342981109408072274_022 scanchain_022/module_data_in[0] scanchain_022/module_data_in[1]
+ scanchain_022/module_data_in[2] scanchain_022/module_data_in[3] scanchain_022/module_data_in[4]
+ scanchain_022/module_data_in[5] scanchain_022/module_data_in[6] scanchain_022/module_data_in[7]
+ scanchain_022/module_data_out[0] scanchain_022/module_data_out[1] scanchain_022/module_data_out[2]
+ scanchain_022/module_data_out[3] scanchain_022/module_data_out[4] scanchain_022/module_data_out[5]
+ scanchain_022/module_data_out[6] scanchain_022/module_data_out[7] vccd1 vssd1 user_module_342981109408072274
Xtt2_tholin_diceroll_060 scanchain_060/module_data_in[0] scanchain_060/module_data_in[1]
+ scanchain_060/module_data_in[2] scanchain_060/module_data_in[3] scanchain_060/module_data_in[4]
+ scanchain_060/module_data_in[5] scanchain_060/module_data_in[6] scanchain_060/module_data_in[7]
+ scanchain_060/module_data_out[0] scanchain_060/module_data_out[1] scanchain_060/module_data_out[2]
+ scanchain_060/module_data_out[3] scanchain_060/module_data_out[4] scanchain_060/module_data_out[5]
+ scanchain_060/module_data_out[6] scanchain_060/module_data_out[7] vccd1 vssd1 tt2_tholin_diceroll
Xuser_module_nickoe_058 user_module_nickoe_058/io_in[0] user_module_nickoe_058/io_in[1]
+ user_module_nickoe_058/io_in[2] user_module_nickoe_058/io_in[3] user_module_nickoe_058/io_in[4]
+ user_module_nickoe_058/io_in[5] user_module_nickoe_058/io_in[6] user_module_nickoe_058/io_in[7]
+ user_module_nickoe_058/io_out[0] user_module_nickoe_058/io_out[1] user_module_nickoe_058/io_out[2]
+ user_module_nickoe_058/io_out[3] user_module_nickoe_058/io_out[4] user_module_nickoe_058/io_out[5]
+ user_module_nickoe_058/io_out[6] user_module_nickoe_058/io_out[7] vccd1 vssd1 user_module_nickoe
Xscanchain_103 scanchain_103/clk_in scanchain_104/clk_in scanchain_103/data_in scanchain_104/data_in
+ scanchain_103/latch_enable_in scanchain_104/latch_enable_in scanchain_103/module_data_in[0]
+ scanchain_103/module_data_in[1] scanchain_103/module_data_in[2] scanchain_103/module_data_in[3]
+ scanchain_103/module_data_in[4] scanchain_103/module_data_in[5] scanchain_103/module_data_in[6]
+ scanchain_103/module_data_in[7] scanchain_103/module_data_out[0] scanchain_103/module_data_out[1]
+ scanchain_103/module_data_out[2] scanchain_103/module_data_out[3] scanchain_103/module_data_out[4]
+ scanchain_103/module_data_out[5] scanchain_103/module_data_out[6] scanchain_103/module_data_out[7]
+ scanchain_103/scan_select_in scanchain_104/scan_select_in vccd1 vssd1 scanchain
Xscanchain_114 scanchain_114/clk_in scanchain_115/clk_in scanchain_114/data_in scanchain_115/data_in
+ scanchain_114/latch_enable_in scanchain_115/latch_enable_in scanchain_114/module_data_in[0]
+ scanchain_114/module_data_in[1] scanchain_114/module_data_in[2] scanchain_114/module_data_in[3]
+ scanchain_114/module_data_in[4] scanchain_114/module_data_in[5] scanchain_114/module_data_in[6]
+ scanchain_114/module_data_in[7] scanchain_114/module_data_out[0] scanchain_114/module_data_out[1]
+ scanchain_114/module_data_out[2] scanchain_114/module_data_out[3] scanchain_114/module_data_out[4]
+ scanchain_114/module_data_out[5] scanchain_114/module_data_out[6] scanchain_114/module_data_out[7]
+ scanchain_114/scan_select_in scanchain_115/scan_select_in vccd1 vssd1 scanchain
Xscanchain_136 scanchain_136/clk_in scanchain_137/clk_in scanchain_136/data_in scanchain_137/data_in
+ scanchain_136/latch_enable_in scanchain_137/latch_enable_in scanchain_136/module_data_in[0]
+ scanchain_136/module_data_in[1] scanchain_136/module_data_in[2] scanchain_136/module_data_in[3]
+ scanchain_136/module_data_in[4] scanchain_136/module_data_in[5] scanchain_136/module_data_in[6]
+ scanchain_136/module_data_in[7] scanchain_136/module_data_out[0] scanchain_136/module_data_out[1]
+ scanchain_136/module_data_out[2] scanchain_136/module_data_out[3] scanchain_136/module_data_out[4]
+ scanchain_136/module_data_out[5] scanchain_136/module_data_out[6] scanchain_136/module_data_out[7]
+ scanchain_136/scan_select_in scanchain_137/scan_select_in vccd1 vssd1 scanchain
Xscanchain_125 scanchain_125/clk_in scanchain_126/clk_in scanchain_125/data_in scanchain_126/data_in
+ scanchain_125/latch_enable_in scanchain_126/latch_enable_in scanchain_125/module_data_in[0]
+ scanchain_125/module_data_in[1] scanchain_125/module_data_in[2] scanchain_125/module_data_in[3]
+ scanchain_125/module_data_in[4] scanchain_125/module_data_in[5] scanchain_125/module_data_in[6]
+ scanchain_125/module_data_in[7] scanchain_125/module_data_out[0] scanchain_125/module_data_out[1]
+ scanchain_125/module_data_out[2] scanchain_125/module_data_out[3] scanchain_125/module_data_out[4]
+ scanchain_125/module_data_out[5] scanchain_125/module_data_out[6] scanchain_125/module_data_out[7]
+ scanchain_125/scan_select_in scanchain_126/scan_select_in vccd1 vssd1 scanchain
Xscanchain_147 scanchain_147/clk_in scanchain_148/clk_in scanchain_147/data_in scanchain_148/data_in
+ scanchain_147/latch_enable_in scanchain_148/latch_enable_in scanchain_147/module_data_in[0]
+ scanchain_147/module_data_in[1] scanchain_147/module_data_in[2] scanchain_147/module_data_in[3]
+ scanchain_147/module_data_in[4] scanchain_147/module_data_in[5] scanchain_147/module_data_in[6]
+ scanchain_147/module_data_in[7] scanchain_147/module_data_out[0] scanchain_147/module_data_out[1]
+ scanchain_147/module_data_out[2] scanchain_147/module_data_out[3] scanchain_147/module_data_out[4]
+ scanchain_147/module_data_out[5] scanchain_147/module_data_out[6] scanchain_147/module_data_out[7]
+ scanchain_147/scan_select_in scanchain_148/scan_select_in vccd1 vssd1 scanchain
Xscanchain_158 scanchain_158/clk_in scanchain_159/clk_in scanchain_158/data_in scanchain_159/data_in
+ scanchain_158/latch_enable_in scanchain_159/latch_enable_in scanchain_158/module_data_in[0]
+ scanchain_158/module_data_in[1] scanchain_158/module_data_in[2] scanchain_158/module_data_in[3]
+ scanchain_158/module_data_in[4] scanchain_158/module_data_in[5] scanchain_158/module_data_in[6]
+ scanchain_158/module_data_in[7] scanchain_158/module_data_out[0] scanchain_158/module_data_out[1]
+ scanchain_158/module_data_out[2] scanchain_158/module_data_out[3] scanchain_158/module_data_out[4]
+ scanchain_158/module_data_out[5] scanchain_158/module_data_out[6] scanchain_158/module_data_out[7]
+ scanchain_158/scan_select_in scanchain_159/scan_select_in vccd1 vssd1 scanchain
Xscanchain_169 scanchain_169/clk_in scanchain_170/clk_in scanchain_169/data_in scanchain_170/data_in
+ scanchain_169/latch_enable_in scanchain_170/latch_enable_in scanchain_169/module_data_in[0]
+ scanchain_169/module_data_in[1] scanchain_169/module_data_in[2] scanchain_169/module_data_in[3]
+ scanchain_169/module_data_in[4] scanchain_169/module_data_in[5] scanchain_169/module_data_in[6]
+ scanchain_169/module_data_in[7] scanchain_169/module_data_out[0] scanchain_169/module_data_out[1]
+ scanchain_169/module_data_out[2] scanchain_169/module_data_out[3] scanchain_169/module_data_out[4]
+ scanchain_169/module_data_out[5] scanchain_169/module_data_out[6] scanchain_169/module_data_out[7]
+ scanchain_169/scan_select_in scanchain_170/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_108 scanchain_108/module_data_in[0] scanchain_108/module_data_in[1]
+ scanchain_108/module_data_in[2] scanchain_108/module_data_in[3] scanchain_108/module_data_in[4]
+ scanchain_108/module_data_in[5] scanchain_108/module_data_in[6] scanchain_108/module_data_in[7]
+ scanchain_108/module_data_out[0] scanchain_108/module_data_out[1] scanchain_108/module_data_out[2]
+ scanchain_108/module_data_out[3] scanchain_108/module_data_out[4] scanchain_108/module_data_out[5]
+ scanchain_108/module_data_out[6] scanchain_108/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_119 scanchain_119/module_data_in[0] scanchain_119/module_data_in[1]
+ scanchain_119/module_data_in[2] scanchain_119/module_data_in[3] scanchain_119/module_data_in[4]
+ scanchain_119/module_data_in[5] scanchain_119/module_data_in[6] scanchain_119/module_data_in[7]
+ scanchain_119/module_data_out[0] scanchain_119/module_data_out[1] scanchain_119/module_data_out[2]
+ scanchain_119/module_data_out[3] scanchain_119/module_data_out[4] scanchain_119/module_data_out[5]
+ scanchain_119/module_data_out[6] scanchain_119/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341541108650607187_047 scanchain_047/module_data_in[0] scanchain_047/module_data_in[1]
+ scanchain_047/module_data_in[2] scanchain_047/module_data_in[3] scanchain_047/module_data_in[4]
+ scanchain_047/module_data_in[5] scanchain_047/module_data_in[6] scanchain_047/module_data_in[7]
+ scanchain_047/module_data_out[0] scanchain_047/module_data_out[1] scanchain_047/module_data_out[2]
+ scanchain_047/module_data_out[3] scanchain_047/module_data_out[4] scanchain_047/module_data_out[5]
+ scanchain_047/module_data_out[6] scanchain_047/module_data_out[7] vccd1 vssd1 user_module_341541108650607187
Xuser_module_349546262775726676_086 scanchain_086/module_data_in[0] scanchain_086/module_data_in[1]
+ scanchain_086/module_data_in[2] scanchain_086/module_data_in[3] scanchain_086/module_data_in[4]
+ scanchain_086/module_data_in[5] scanchain_086/module_data_in[6] scanchain_086/module_data_in[7]
+ scanchain_086/module_data_out[0] scanchain_086/module_data_out[1] scanchain_086/module_data_out[2]
+ scanchain_086/module_data_out[3] scanchain_086/module_data_out[4] scanchain_086/module_data_out[5]
+ scanchain_086/module_data_out[6] scanchain_086/module_data_out[7] vccd1 vssd1 user_module_349546262775726676
Xscanchain_104 scanchain_104/clk_in scanchain_105/clk_in scanchain_104/data_in scanchain_105/data_in
+ scanchain_104/latch_enable_in scanchain_105/latch_enable_in scanchain_104/module_data_in[0]
+ scanchain_104/module_data_in[1] scanchain_104/module_data_in[2] scanchain_104/module_data_in[3]
+ scanchain_104/module_data_in[4] scanchain_104/module_data_in[5] scanchain_104/module_data_in[6]
+ scanchain_104/module_data_in[7] scanchain_104/module_data_out[0] scanchain_104/module_data_out[1]
+ scanchain_104/module_data_out[2] scanchain_104/module_data_out[3] scanchain_104/module_data_out[4]
+ scanchain_104/module_data_out[5] scanchain_104/module_data_out[6] scanchain_104/module_data_out[7]
+ scanchain_104/scan_select_in scanchain_105/scan_select_in vccd1 vssd1 scanchain
Xscanchain_115 scanchain_115/clk_in scanchain_116/clk_in scanchain_115/data_in scanchain_116/data_in
+ scanchain_115/latch_enable_in scanchain_116/latch_enable_in scanchain_115/module_data_in[0]
+ scanchain_115/module_data_in[1] scanchain_115/module_data_in[2] scanchain_115/module_data_in[3]
+ scanchain_115/module_data_in[4] scanchain_115/module_data_in[5] scanchain_115/module_data_in[6]
+ scanchain_115/module_data_in[7] scanchain_115/module_data_out[0] scanchain_115/module_data_out[1]
+ scanchain_115/module_data_out[2] scanchain_115/module_data_out[3] scanchain_115/module_data_out[4]
+ scanchain_115/module_data_out[5] scanchain_115/module_data_out[6] scanchain_115/module_data_out[7]
+ scanchain_115/scan_select_in scanchain_116/scan_select_in vccd1 vssd1 scanchain
Xscanchain_137 scanchain_137/clk_in scanchain_138/clk_in scanchain_137/data_in scanchain_138/data_in
+ scanchain_137/latch_enable_in scanchain_138/latch_enable_in scanchain_137/module_data_in[0]
+ scanchain_137/module_data_in[1] scanchain_137/module_data_in[2] scanchain_137/module_data_in[3]
+ scanchain_137/module_data_in[4] scanchain_137/module_data_in[5] scanchain_137/module_data_in[6]
+ scanchain_137/module_data_in[7] scanchain_137/module_data_out[0] scanchain_137/module_data_out[1]
+ scanchain_137/module_data_out[2] scanchain_137/module_data_out[3] scanchain_137/module_data_out[4]
+ scanchain_137/module_data_out[5] scanchain_137/module_data_out[6] scanchain_137/module_data_out[7]
+ scanchain_137/scan_select_in scanchain_138/scan_select_in vccd1 vssd1 scanchain
Xscanchain_126 scanchain_126/clk_in scanchain_127/clk_in scanchain_126/data_in scanchain_127/data_in
+ scanchain_126/latch_enable_in scanchain_127/latch_enable_in scanchain_126/module_data_in[0]
+ scanchain_126/module_data_in[1] scanchain_126/module_data_in[2] scanchain_126/module_data_in[3]
+ scanchain_126/module_data_in[4] scanchain_126/module_data_in[5] scanchain_126/module_data_in[6]
+ scanchain_126/module_data_in[7] scanchain_126/module_data_out[0] scanchain_126/module_data_out[1]
+ scanchain_126/module_data_out[2] scanchain_126/module_data_out[3] scanchain_126/module_data_out[4]
+ scanchain_126/module_data_out[5] scanchain_126/module_data_out[6] scanchain_126/module_data_out[7]
+ scanchain_126/scan_select_in scanchain_127/scan_select_in vccd1 vssd1 scanchain
Xscanchain_148 scanchain_148/clk_in scanchain_149/clk_in scanchain_148/data_in scanchain_149/data_in
+ scanchain_148/latch_enable_in scanchain_149/latch_enable_in scanchain_148/module_data_in[0]
+ scanchain_148/module_data_in[1] scanchain_148/module_data_in[2] scanchain_148/module_data_in[3]
+ scanchain_148/module_data_in[4] scanchain_148/module_data_in[5] scanchain_148/module_data_in[6]
+ scanchain_148/module_data_in[7] scanchain_148/module_data_out[0] scanchain_148/module_data_out[1]
+ scanchain_148/module_data_out[2] scanchain_148/module_data_out[3] scanchain_148/module_data_out[4]
+ scanchain_148/module_data_out[5] scanchain_148/module_data_out[6] scanchain_148/module_data_out[7]
+ scanchain_148/scan_select_in scanchain_149/scan_select_in vccd1 vssd1 scanchain
Xscanchain_159 scanchain_159/clk_in scanchain_160/clk_in scanchain_159/data_in scanchain_160/data_in
+ scanchain_159/latch_enable_in scanchain_160/latch_enable_in scanchain_159/module_data_in[0]
+ scanchain_159/module_data_in[1] scanchain_159/module_data_in[2] scanchain_159/module_data_in[3]
+ scanchain_159/module_data_in[4] scanchain_159/module_data_in[5] scanchain_159/module_data_in[6]
+ scanchain_159/module_data_in[7] scanchain_159/module_data_out[0] scanchain_159/module_data_out[1]
+ scanchain_159/module_data_out[2] scanchain_159/module_data_out[3] scanchain_159/module_data_out[4]
+ scanchain_159/module_data_out[5] scanchain_159/module_data_out[6] scanchain_159/module_data_out[7]
+ scanchain_159/scan_select_in scanchain_160/scan_select_in vccd1 vssd1 scanchain
Xgithub_com_proppy_tt02_xls_popcount_042 scanchain_042/module_data_in[0] scanchain_042/module_data_in[1]
+ scanchain_042/module_data_in[2] scanchain_042/module_data_in[3] scanchain_042/module_data_in[4]
+ scanchain_042/module_data_in[5] scanchain_042/module_data_in[6] scanchain_042/module_data_in[7]
+ scanchain_042/module_data_out[0] scanchain_042/module_data_out[1] scanchain_042/module_data_out[2]
+ scanchain_042/module_data_out[3] scanchain_042/module_data_out[4] scanchain_042/module_data_out[5]
+ scanchain_042/module_data_out[6] scanchain_042/module_data_out[7] vccd1 vssd1 github_com_proppy_tt02_xls_popcount
Xuser_module_341614374571475540_044 scanchain_044/module_data_in[0] scanchain_044/module_data_in[1]
+ scanchain_044/module_data_in[2] scanchain_044/module_data_in[3] scanchain_044/module_data_in[4]
+ scanchain_044/module_data_in[5] scanchain_044/module_data_in[6] scanchain_044/module_data_in[7]
+ scanchain_044/module_data_out[0] scanchain_044/module_data_out[1] scanchain_044/module_data_out[2]
+ scanchain_044/module_data_out[3] scanchain_044/module_data_out[4] scanchain_044/module_data_out[5]
+ scanchain_044/module_data_out[6] scanchain_044/module_data_out[7] vccd1 vssd1 user_module_341614374571475540
Xkrasin_tt02_verilog_spi_7_channel_pwm_driver_072 scanchain_072/module_data_in[0]
+ scanchain_072/module_data_in[1] scanchain_072/module_data_in[2] scanchain_072/module_data_in[3]
+ scanchain_072/module_data_in[4] scanchain_072/module_data_in[5] scanchain_072/module_data_in[6]
+ scanchain_072/module_data_in[7] scanchain_072/module_data_out[0] scanchain_072/module_data_out[1]
+ scanchain_072/module_data_out[2] scanchain_072/module_data_out[3] scanchain_072/module_data_out[4]
+ scanchain_072/module_data_out[5] scanchain_072/module_data_out[6] scanchain_072/module_data_out[7]
+ vccd1 vssd1 krasin_tt02_verilog_spi_7_channel_pwm_driver
Xuser_module_341535056611770964_109 scanchain_109/module_data_in[0] scanchain_109/module_data_in[1]
+ scanchain_109/module_data_in[2] scanchain_109/module_data_in[3] scanchain_109/module_data_in[4]
+ scanchain_109/module_data_in[5] scanchain_109/module_data_in[6] scanchain_109/module_data_in[7]
+ scanchain_109/module_data_out[0] scanchain_109/module_data_out[1] scanchain_109/module_data_out[2]
+ scanchain_109/module_data_out[3] scanchain_109/module_data_out[4] scanchain_109/module_data_out[5]
+ scanchain_109/module_data_out[6] scanchain_109/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_105 scanchain_105/clk_in scanchain_106/clk_in scanchain_105/data_in scanchain_106/data_in
+ scanchain_105/latch_enable_in scanchain_106/latch_enable_in scanchain_105/module_data_in[0]
+ scanchain_105/module_data_in[1] scanchain_105/module_data_in[2] scanchain_105/module_data_in[3]
+ scanchain_105/module_data_in[4] scanchain_105/module_data_in[5] scanchain_105/module_data_in[6]
+ scanchain_105/module_data_in[7] scanchain_105/module_data_out[0] scanchain_105/module_data_out[1]
+ scanchain_105/module_data_out[2] scanchain_105/module_data_out[3] scanchain_105/module_data_out[4]
+ scanchain_105/module_data_out[5] scanchain_105/module_data_out[6] scanchain_105/module_data_out[7]
+ scanchain_105/scan_select_in scanchain_106/scan_select_in vccd1 vssd1 scanchain
Xscanchain_116 scanchain_116/clk_in scanchain_117/clk_in scanchain_116/data_in scanchain_117/data_in
+ scanchain_116/latch_enable_in scanchain_117/latch_enable_in scanchain_116/module_data_in[0]
+ scanchain_116/module_data_in[1] scanchain_116/module_data_in[2] scanchain_116/module_data_in[3]
+ scanchain_116/module_data_in[4] scanchain_116/module_data_in[5] scanchain_116/module_data_in[6]
+ scanchain_116/module_data_in[7] scanchain_116/module_data_out[0] scanchain_116/module_data_out[1]
+ scanchain_116/module_data_out[2] scanchain_116/module_data_out[3] scanchain_116/module_data_out[4]
+ scanchain_116/module_data_out[5] scanchain_116/module_data_out[6] scanchain_116/module_data_out[7]
+ scanchain_116/scan_select_in scanchain_117/scan_select_in vccd1 vssd1 scanchain
Xscanchain_127 scanchain_127/clk_in scanchain_128/clk_in scanchain_127/data_in scanchain_128/data_in
+ scanchain_127/latch_enable_in scanchain_128/latch_enable_in scanchain_127/module_data_in[0]
+ scanchain_127/module_data_in[1] scanchain_127/module_data_in[2] scanchain_127/module_data_in[3]
+ scanchain_127/module_data_in[4] scanchain_127/module_data_in[5] scanchain_127/module_data_in[6]
+ scanchain_127/module_data_in[7] scanchain_127/module_data_out[0] scanchain_127/module_data_out[1]
+ scanchain_127/module_data_out[2] scanchain_127/module_data_out[3] scanchain_127/module_data_out[4]
+ scanchain_127/module_data_out[5] scanchain_127/module_data_out[6] scanchain_127/module_data_out[7]
+ scanchain_127/scan_select_in scanchain_128/scan_select_in vccd1 vssd1 scanchain
Xscanchain_138 scanchain_138/clk_in scanchain_139/clk_in scanchain_138/data_in scanchain_139/data_in
+ scanchain_138/latch_enable_in scanchain_139/latch_enable_in scanchain_138/module_data_in[0]
+ scanchain_138/module_data_in[1] scanchain_138/module_data_in[2] scanchain_138/module_data_in[3]
+ scanchain_138/module_data_in[4] scanchain_138/module_data_in[5] scanchain_138/module_data_in[6]
+ scanchain_138/module_data_in[7] scanchain_138/module_data_out[0] scanchain_138/module_data_out[1]
+ scanchain_138/module_data_out[2] scanchain_138/module_data_out[3] scanchain_138/module_data_out[4]
+ scanchain_138/module_data_out[5] scanchain_138/module_data_out[6] scanchain_138/module_data_out[7]
+ scanchain_138/scan_select_in scanchain_139/scan_select_in vccd1 vssd1 scanchain
Xscanchain_149 scanchain_149/clk_in scanchain_150/clk_in scanchain_149/data_in scanchain_150/data_in
+ scanchain_149/latch_enable_in scanchain_150/latch_enable_in scanchain_149/module_data_in[0]
+ scanchain_149/module_data_in[1] scanchain_149/module_data_in[2] scanchain_149/module_data_in[3]
+ scanchain_149/module_data_in[4] scanchain_149/module_data_in[5] scanchain_149/module_data_in[6]
+ scanchain_149/module_data_in[7] scanchain_149/module_data_out[0] scanchain_149/module_data_out[1]
+ scanchain_149/module_data_out[2] scanchain_149/module_data_out[3] scanchain_149/module_data_out[4]
+ scanchain_149/module_data_out[5] scanchain_149/module_data_out[6] scanchain_149/module_data_out[7]
+ scanchain_149/scan_select_in scanchain_150/scan_select_in vccd1 vssd1 scanchain
Xudxs_sqrt_top_066 udxs_sqrt_top_066/io_in[0] udxs_sqrt_top_066/io_in[1] udxs_sqrt_top_066/io_in[2]
+ udxs_sqrt_top_066/io_in[3] udxs_sqrt_top_066/io_in[4] udxs_sqrt_top_066/io_in[5]
+ udxs_sqrt_top_066/io_in[6] udxs_sqrt_top_066/io_in[7] udxs_sqrt_top_066/io_out[0]
+ udxs_sqrt_top_066/io_out[1] udxs_sqrt_top_066/io_out[2] udxs_sqrt_top_066/io_out[3]
+ udxs_sqrt_top_066/io_out[4] udxs_sqrt_top_066/io_out[5] udxs_sqrt_top_066/io_out[6]
+ udxs_sqrt_top_066/io_out[7] vccd1 vssd1 udxs_sqrt_top
Xmoonbase_cpu_8bit_084 moonbase_cpu_8bit_084/io_in[0] moonbase_cpu_8bit_084/io_in[1]
+ moonbase_cpu_8bit_084/io_in[2] moonbase_cpu_8bit_084/io_in[3] moonbase_cpu_8bit_084/io_in[4]
+ moonbase_cpu_8bit_084/io_in[5] moonbase_cpu_8bit_084/io_in[6] moonbase_cpu_8bit_084/io_in[7]
+ moonbase_cpu_8bit_084/io_out[0] moonbase_cpu_8bit_084/io_out[1] moonbase_cpu_8bit_084/io_out[2]
+ moonbase_cpu_8bit_084/io_out[3] moonbase_cpu_8bit_084/io_out[4] moonbase_cpu_8bit_084/io_out[5]
+ moonbase_cpu_8bit_084/io_out[6] moonbase_cpu_8bit_084/io_out[7] vccd1 vssd1 moonbase_cpu_8bit
Xloxodes_sequencer_004 loxodes_sequencer_004/io_in[0] loxodes_sequencer_004/io_in[1]
+ loxodes_sequencer_004/io_in[2] loxodes_sequencer_004/io_in[3] loxodes_sequencer_004/io_in[4]
+ loxodes_sequencer_004/io_in[5] loxodes_sequencer_004/io_in[6] loxodes_sequencer_004/io_in[7]
+ loxodes_sequencer_004/io_out[0] loxodes_sequencer_004/io_out[1] loxodes_sequencer_004/io_out[2]
+ loxodes_sequencer_004/io_out[3] loxodes_sequencer_004/io_out[4] loxodes_sequencer_004/io_out[5]
+ loxodes_sequencer_004/io_out[6] loxodes_sequencer_004/io_out[7] vccd1 vssd1 loxodes_sequencer
Xscanchain_106 scanchain_106/clk_in scanchain_107/clk_in scanchain_106/data_in scanchain_107/data_in
+ scanchain_106/latch_enable_in scanchain_107/latch_enable_in scanchain_106/module_data_in[0]
+ scanchain_106/module_data_in[1] scanchain_106/module_data_in[2] scanchain_106/module_data_in[3]
+ scanchain_106/module_data_in[4] scanchain_106/module_data_in[5] scanchain_106/module_data_in[6]
+ scanchain_106/module_data_in[7] scanchain_106/module_data_out[0] scanchain_106/module_data_out[1]
+ scanchain_106/module_data_out[2] scanchain_106/module_data_out[3] scanchain_106/module_data_out[4]
+ scanchain_106/module_data_out[5] scanchain_106/module_data_out[6] scanchain_106/module_data_out[7]
+ scanchain_106/scan_select_in scanchain_107/scan_select_in vccd1 vssd1 scanchain
Xscanchain_117 scanchain_117/clk_in scanchain_118/clk_in scanchain_117/data_in scanchain_118/data_in
+ scanchain_117/latch_enable_in scanchain_118/latch_enable_in scanchain_117/module_data_in[0]
+ scanchain_117/module_data_in[1] scanchain_117/module_data_in[2] scanchain_117/module_data_in[3]
+ scanchain_117/module_data_in[4] scanchain_117/module_data_in[5] scanchain_117/module_data_in[6]
+ scanchain_117/module_data_in[7] scanchain_117/module_data_out[0] scanchain_117/module_data_out[1]
+ scanchain_117/module_data_out[2] scanchain_117/module_data_out[3] scanchain_117/module_data_out[4]
+ scanchain_117/module_data_out[5] scanchain_117/module_data_out[6] scanchain_117/module_data_out[7]
+ scanchain_117/scan_select_in scanchain_118/scan_select_in vccd1 vssd1 scanchain
Xscanchain_128 scanchain_128/clk_in scanchain_129/clk_in scanchain_128/data_in scanchain_129/data_in
+ scanchain_128/latch_enable_in scanchain_129/latch_enable_in scanchain_128/module_data_in[0]
+ scanchain_128/module_data_in[1] scanchain_128/module_data_in[2] scanchain_128/module_data_in[3]
+ scanchain_128/module_data_in[4] scanchain_128/module_data_in[5] scanchain_128/module_data_in[6]
+ scanchain_128/module_data_in[7] scanchain_128/module_data_out[0] scanchain_128/module_data_out[1]
+ scanchain_128/module_data_out[2] scanchain_128/module_data_out[3] scanchain_128/module_data_out[4]
+ scanchain_128/module_data_out[5] scanchain_128/module_data_out[6] scanchain_128/module_data_out[7]
+ scanchain_128/scan_select_in scanchain_129/scan_select_in vccd1 vssd1 scanchain
Xscanchain_139 scanchain_139/clk_in scanchain_140/clk_in scanchain_139/data_in scanchain_140/data_in
+ scanchain_139/latch_enable_in scanchain_140/latch_enable_in scanchain_139/module_data_in[0]
+ scanchain_139/module_data_in[1] scanchain_139/module_data_in[2] scanchain_139/module_data_in[3]
+ scanchain_139/module_data_in[4] scanchain_139/module_data_in[5] scanchain_139/module_data_in[6]
+ scanchain_139/module_data_in[7] scanchain_139/module_data_out[0] scanchain_139/module_data_out[1]
+ scanchain_139/module_data_out[2] scanchain_139/module_data_out[3] scanchain_139/module_data_out[4]
+ scanchain_139/module_data_out[5] scanchain_139/module_data_out[6] scanchain_139/module_data_out[7]
+ scanchain_139/scan_select_in scanchain_140/scan_select_in vccd1 vssd1 scanchain
Xuser_module_347594509754827347_019 scanchain_019/module_data_in[0] scanchain_019/module_data_in[1]
+ scanchain_019/module_data_in[2] scanchain_019/module_data_in[3] scanchain_019/module_data_in[4]
+ scanchain_019/module_data_in[5] scanchain_019/module_data_in[6] scanchain_019/module_data_in[7]
+ scanchain_019/module_data_out[0] scanchain_019/module_data_out[1] scanchain_019/module_data_out[2]
+ scanchain_019/module_data_out[3] scanchain_019/module_data_out[4] scanchain_019/module_data_out[5]
+ scanchain_019/module_data_out[6] scanchain_019/module_data_out[7] vccd1 vssd1 user_module_347594509754827347
Xyupferris_bitslam_040 yupferris_bitslam_040/io_in[0] yupferris_bitslam_040/io_in[1]
+ yupferris_bitslam_040/io_in[2] yupferris_bitslam_040/io_in[3] yupferris_bitslam_040/io_in[4]
+ yupferris_bitslam_040/io_in[5] yupferris_bitslam_040/io_in[6] yupferris_bitslam_040/io_in[7]
+ yupferris_bitslam_040/io_out[0] yupferris_bitslam_040/io_out[1] yupferris_bitslam_040/io_out[2]
+ yupferris_bitslam_040/io_out[3] yupferris_bitslam_040/io_out[4] yupferris_bitslam_040/io_out[5]
+ yupferris_bitslam_040/io_out[6] yupferris_bitslam_040/io_out[7] vccd1 vssd1 yupferris_bitslam
Xphasenoisepon_seven_segment_seconds_046 scanchain_046/module_data_in[0] scanchain_046/module_data_in[1]
+ scanchain_046/module_data_in[2] scanchain_046/module_data_in[3] scanchain_046/module_data_in[4]
+ scanchain_046/module_data_in[5] scanchain_046/module_data_in[6] scanchain_046/module_data_in[7]
+ scanchain_046/module_data_out[0] scanchain_046/module_data_out[1] scanchain_046/module_data_out[2]
+ scanchain_046/module_data_out[3] scanchain_046/module_data_out[4] scanchain_046/module_data_out[5]
+ scanchain_046/module_data_out[6] scanchain_046/module_data_out[7] vccd1 vssd1 phasenoisepon_seven_segment_seconds
Xuser_module_348961139276644947_062 scanchain_062/module_data_in[0] scanchain_062/module_data_in[1]
+ scanchain_062/module_data_in[2] scanchain_062/module_data_in[3] scanchain_062/module_data_in[4]
+ scanchain_062/module_data_in[5] scanchain_062/module_data_in[6] scanchain_062/module_data_in[7]
+ scanchain_062/module_data_out[0] scanchain_062/module_data_out[1] scanchain_062/module_data_out[2]
+ scanchain_062/module_data_out[3] scanchain_062/module_data_out[4] scanchain_062/module_data_out[5]
+ scanchain_062/module_data_out[6] scanchain_062/module_data_out[7] vccd1 vssd1 user_module_348961139276644947
Xmigcorre_pwm_005 migcorre_pwm_005/io_in[0] migcorre_pwm_005/io_in[1] migcorre_pwm_005/io_in[2]
+ migcorre_pwm_005/io_in[3] migcorre_pwm_005/io_in[4] migcorre_pwm_005/io_in[5] migcorre_pwm_005/io_in[6]
+ migcorre_pwm_005/io_in[7] migcorre_pwm_005/io_out[0] migcorre_pwm_005/io_out[1]
+ migcorre_pwm_005/io_out[2] migcorre_pwm_005/io_out[3] migcorre_pwm_005/io_out[4]
+ migcorre_pwm_005/io_out[5] migcorre_pwm_005/io_out[6] migcorre_pwm_005/io_out[7]
+ vccd1 vssd1 migcorre_pwm
Xscanchain_107 scanchain_107/clk_in scanchain_108/clk_in scanchain_107/data_in scanchain_108/data_in
+ scanchain_107/latch_enable_in scanchain_108/latch_enable_in scanchain_107/module_data_in[0]
+ scanchain_107/module_data_in[1] scanchain_107/module_data_in[2] scanchain_107/module_data_in[3]
+ scanchain_107/module_data_in[4] scanchain_107/module_data_in[5] scanchain_107/module_data_in[6]
+ scanchain_107/module_data_in[7] scanchain_107/module_data_out[0] scanchain_107/module_data_out[1]
+ scanchain_107/module_data_out[2] scanchain_107/module_data_out[3] scanchain_107/module_data_out[4]
+ scanchain_107/module_data_out[5] scanchain_107/module_data_out[6] scanchain_107/module_data_out[7]
+ scanchain_107/scan_select_in scanchain_108/scan_select_in vccd1 vssd1 scanchain
Xscanchain_118 scanchain_118/clk_in scanchain_119/clk_in scanchain_118/data_in scanchain_119/data_in
+ scanchain_118/latch_enable_in scanchain_119/latch_enable_in scanchain_118/module_data_in[0]
+ scanchain_118/module_data_in[1] scanchain_118/module_data_in[2] scanchain_118/module_data_in[3]
+ scanchain_118/module_data_in[4] scanchain_118/module_data_in[5] scanchain_118/module_data_in[6]
+ scanchain_118/module_data_in[7] scanchain_118/module_data_out[0] scanchain_118/module_data_out[1]
+ scanchain_118/module_data_out[2] scanchain_118/module_data_out[3] scanchain_118/module_data_out[4]
+ scanchain_118/module_data_out[5] scanchain_118/module_data_out[6] scanchain_118/module_data_out[7]
+ scanchain_118/scan_select_in scanchain_119/scan_select_in vccd1 vssd1 scanchain
Xscanchain_129 scanchain_129/clk_in scanchain_130/clk_in scanchain_129/data_in scanchain_130/data_in
+ scanchain_129/latch_enable_in scanchain_130/latch_enable_in scanchain_129/module_data_in[0]
+ scanchain_129/module_data_in[1] scanchain_129/module_data_in[2] scanchain_129/module_data_in[3]
+ scanchain_129/module_data_in[4] scanchain_129/module_data_in[5] scanchain_129/module_data_in[6]
+ scanchain_129/module_data_in[7] scanchain_129/module_data_out[0] scanchain_129/module_data_out[1]
+ scanchain_129/module_data_out[2] scanchain_129/module_data_out[3] scanchain_129/module_data_out[4]
+ scanchain_129/module_data_out[5] scanchain_129/module_data_out[6] scanchain_129/module_data_out[7]
+ scanchain_129/scan_select_in scanchain_130/scan_select_in vccd1 vssd1 scanchain
Xuser_module_346553315158393428_016 scanchain_016/module_data_in[0] scanchain_016/module_data_in[1]
+ scanchain_016/module_data_in[2] scanchain_016/module_data_in[3] scanchain_016/module_data_in[4]
+ scanchain_016/module_data_in[5] scanchain_016/module_data_in[6] scanchain_016/module_data_in[7]
+ scanchain_016/module_data_out[0] scanchain_016/module_data_out[1] scanchain_016/module_data_out[2]
+ scanchain_016/module_data_out[3] scanchain_016/module_data_out[4] scanchain_016/module_data_out[5]
+ scanchain_016/module_data_out[6] scanchain_016/module_data_out[7] vccd1 vssd1 user_module_346553315158393428
Xjar_sram_top_011 jar_sram_top_011/io_in[0] jar_sram_top_011/io_in[1] jar_sram_top_011/io_in[2]
+ jar_sram_top_011/io_in[3] jar_sram_top_011/io_in[4] jar_sram_top_011/io_in[5] jar_sram_top_011/io_in[6]
+ jar_sram_top_011/io_in[7] jar_sram_top_011/io_out[0] jar_sram_top_011/io_out[1]
+ jar_sram_top_011/io_out[2] jar_sram_top_011/io_out[3] jar_sram_top_011/io_out[4]
+ jar_sram_top_011/io_out[5] jar_sram_top_011/io_out[6] jar_sram_top_011/io_out[7]
+ vccd1 vssd1 jar_sram_top
Xuser_module_341535056611770964_240 scanchain_240/module_data_in[0] scanchain_240/module_data_in[1]
+ scanchain_240/module_data_in[2] scanchain_240/module_data_in[3] scanchain_240/module_data_in[4]
+ scanchain_240/module_data_in[5] scanchain_240/module_data_in[6] scanchain_240/module_data_in[7]
+ scanchain_240/module_data_out[0] scanchain_240/module_data_out[1] scanchain_240/module_data_out[2]
+ scanchain_240/module_data_out[3] scanchain_240/module_data_out[4] scanchain_240/module_data_out[5]
+ scanchain_240/module_data_out[6] scanchain_240/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_108 scanchain_108/clk_in scanchain_109/clk_in scanchain_108/data_in scanchain_109/data_in
+ scanchain_108/latch_enable_in scanchain_109/latch_enable_in scanchain_108/module_data_in[0]
+ scanchain_108/module_data_in[1] scanchain_108/module_data_in[2] scanchain_108/module_data_in[3]
+ scanchain_108/module_data_in[4] scanchain_108/module_data_in[5] scanchain_108/module_data_in[6]
+ scanchain_108/module_data_in[7] scanchain_108/module_data_out[0] scanchain_108/module_data_out[1]
+ scanchain_108/module_data_out[2] scanchain_108/module_data_out[3] scanchain_108/module_data_out[4]
+ scanchain_108/module_data_out[5] scanchain_108/module_data_out[6] scanchain_108/module_data_out[7]
+ scanchain_108/scan_select_in scanchain_109/scan_select_in vccd1 vssd1 scanchain
Xscanchain_119 scanchain_119/clk_in scanchain_120/clk_in scanchain_119/data_in scanchain_120/data_in
+ scanchain_119/latch_enable_in scanchain_120/latch_enable_in scanchain_119/module_data_in[0]
+ scanchain_119/module_data_in[1] scanchain_119/module_data_in[2] scanchain_119/module_data_in[3]
+ scanchain_119/module_data_in[4] scanchain_119/module_data_in[5] scanchain_119/module_data_in[6]
+ scanchain_119/module_data_in[7] scanchain_119/module_data_out[0] scanchain_119/module_data_out[1]
+ scanchain_119/module_data_out[2] scanchain_119/module_data_out[3] scanchain_119/module_data_out[4]
+ scanchain_119/module_data_out[5] scanchain_119/module_data_out[6] scanchain_119/module_data_out[7]
+ scanchain_119/scan_select_in scanchain_120/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_241 scanchain_241/module_data_in[0] scanchain_241/module_data_in[1]
+ scanchain_241/module_data_in[2] scanchain_241/module_data_in[3] scanchain_241/module_data_in[4]
+ scanchain_241/module_data_in[5] scanchain_241/module_data_in[6] scanchain_241/module_data_in[7]
+ scanchain_241/module_data_out[0] scanchain_241/module_data_out[1] scanchain_241/module_data_out[2]
+ scanchain_241/module_data_out[3] scanchain_241/module_data_out[4] scanchain_241/module_data_out[5]
+ scanchain_241/module_data_out[6] scanchain_241/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_230 scanchain_230/module_data_in[0] scanchain_230/module_data_in[1]
+ scanchain_230/module_data_in[2] scanchain_230/module_data_in[3] scanchain_230/module_data_in[4]
+ scanchain_230/module_data_in[5] scanchain_230/module_data_in[6] scanchain_230/module_data_in[7]
+ scanchain_230/module_data_out[0] scanchain_230/module_data_out[1] scanchain_230/module_data_out[2]
+ scanchain_230/module_data_out[3] scanchain_230/module_data_out[4] scanchain_230/module_data_out[5]
+ scanchain_230/module_data_out[6] scanchain_230/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_109 scanchain_109/clk_in scanchain_110/clk_in scanchain_109/data_in scanchain_110/data_in
+ scanchain_109/latch_enable_in scanchain_110/latch_enable_in scanchain_109/module_data_in[0]
+ scanchain_109/module_data_in[1] scanchain_109/module_data_in[2] scanchain_109/module_data_in[3]
+ scanchain_109/module_data_in[4] scanchain_109/module_data_in[5] scanchain_109/module_data_in[6]
+ scanchain_109/module_data_in[7] scanchain_109/module_data_out[0] scanchain_109/module_data_out[1]
+ scanchain_109/module_data_out[2] scanchain_109/module_data_out[3] scanchain_109/module_data_out[4]
+ scanchain_109/module_data_out[5] scanchain_109/module_data_out[6] scanchain_109/module_data_out[7]
+ scanchain_109/scan_select_in scanchain_110/scan_select_in vccd1 vssd1 scanchain
Xyubex_egg_timer_029 yubex_egg_timer_029/io_in[0] yubex_egg_timer_029/io_in[1] yubex_egg_timer_029/io_in[2]
+ yubex_egg_timer_029/io_in[3] yubex_egg_timer_029/io_in[4] yubex_egg_timer_029/io_in[5]
+ yubex_egg_timer_029/io_in[6] yubex_egg_timer_029/io_in[7] yubex_egg_timer_029/io_out[0]
+ yubex_egg_timer_029/io_out[1] yubex_egg_timer_029/io_out[2] yubex_egg_timer_029/io_out[3]
+ yubex_egg_timer_029/io_out[4] yubex_egg_timer_029/io_out[5] yubex_egg_timer_029/io_out[6]
+ yubex_egg_timer_029/io_out[7] vccd1 vssd1 yubex_egg_timer
Xflygoat_tt02_play_tune_054 scanchain_054/module_data_in[0] scanchain_054/module_data_in[1]
+ scanchain_054/module_data_in[2] scanchain_054/module_data_in[3] scanchain_054/module_data_in[4]
+ scanchain_054/module_data_in[5] scanchain_054/module_data_in[6] scanchain_054/module_data_in[7]
+ scanchain_054/module_data_out[0] scanchain_054/module_data_out[1] scanchain_054/module_data_out[2]
+ scanchain_054/module_data_out[3] scanchain_054/module_data_out[4] scanchain_054/module_data_out[5]
+ scanchain_054/module_data_out[6] scanchain_054/module_data_out[7] vccd1 vssd1 flygoat_tt02_play_tune
Xs4ga_006 s4ga_006/io_in[0] s4ga_006/io_in[1] s4ga_006/io_in[2] s4ga_006/io_in[3]
+ s4ga_006/io_in[4] s4ga_006/io_in[5] s4ga_006/io_in[6] s4ga_006/io_in[7] s4ga_006/io_out[0]
+ s4ga_006/io_out[1] s4ga_006/io_out[2] s4ga_006/io_out[3] s4ga_006/io_out[4] s4ga_006/io_out[5]
+ s4ga_006/io_out[6] s4ga_006/io_out[7] vccd1 vssd1 s4ga
Xuser_module_341535056611770964_242 scanchain_242/module_data_in[0] scanchain_242/module_data_in[1]
+ scanchain_242/module_data_in[2] scanchain_242/module_data_in[3] scanchain_242/module_data_in[4]
+ scanchain_242/module_data_in[5] scanchain_242/module_data_in[6] scanchain_242/module_data_in[7]
+ scanchain_242/module_data_out[0] scanchain_242/module_data_out[1] scanchain_242/module_data_out[2]
+ scanchain_242/module_data_out[3] scanchain_242/module_data_out[4] scanchain_242/module_data_out[5]
+ scanchain_242/module_data_out[6] scanchain_242/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_231 scanchain_231/module_data_in[0] scanchain_231/module_data_in[1]
+ scanchain_231/module_data_in[2] scanchain_231/module_data_in[3] scanchain_231/module_data_in[4]
+ scanchain_231/module_data_in[5] scanchain_231/module_data_in[6] scanchain_231/module_data_in[7]
+ scanchain_231/module_data_out[0] scanchain_231/module_data_out[1] scanchain_231/module_data_out[2]
+ scanchain_231/module_data_out[3] scanchain_231/module_data_out[4] scanchain_231/module_data_out[5]
+ scanchain_231/module_data_out[6] scanchain_231/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_220 scanchain_220/module_data_in[0] scanchain_220/module_data_in[1]
+ scanchain_220/module_data_in[2] scanchain_220/module_data_in[3] scanchain_220/module_data_in[4]
+ scanchain_220/module_data_in[5] scanchain_220/module_data_in[6] scanchain_220/module_data_in[7]
+ scanchain_220/module_data_out[0] scanchain_220/module_data_out[1] scanchain_220/module_data_out[2]
+ scanchain_220/module_data_out[3] scanchain_220/module_data_out[4] scanchain_220/module_data_out[5]
+ scanchain_220/module_data_out[6] scanchain_220/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xrc5_top_043 rc5_top_043/io_in[0] rc5_top_043/io_in[1] rc5_top_043/io_in[2] rc5_top_043/io_in[3]
+ rc5_top_043/io_in[4] rc5_top_043/io_in[5] rc5_top_043/io_in[6] rc5_top_043/io_in[7]
+ rc5_top_043/io_out[0] rc5_top_043/io_out[1] rc5_top_043/io_out[2] rc5_top_043/io_out[3]
+ rc5_top_043/io_out[4] rc5_top_043/io_out[5] rc5_top_043/io_out[6] rc5_top_043/io_out[7]
+ vccd1 vssd1 rc5_top
Xscanchain_090 scanchain_090/clk_in scanchain_091/clk_in scanchain_090/data_in scanchain_091/data_in
+ scanchain_090/latch_enable_in scanchain_091/latch_enable_in scanchain_090/module_data_in[0]
+ scanchain_090/module_data_in[1] scanchain_090/module_data_in[2] scanchain_090/module_data_in[3]
+ scanchain_090/module_data_in[4] scanchain_090/module_data_in[5] scanchain_090/module_data_in[6]
+ scanchain_090/module_data_in[7] scanchain_090/module_data_out[0] scanchain_090/module_data_out[1]
+ scanchain_090/module_data_out[2] scanchain_090/module_data_out[3] scanchain_090/module_data_out[4]
+ scanchain_090/module_data_out[5] scanchain_090/module_data_out[6] scanchain_090/module_data_out[7]
+ scanchain_090/scan_select_in scanchain_091/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_243 scanchain_243/module_data_in[0] scanchain_243/module_data_in[1]
+ scanchain_243/module_data_in[2] scanchain_243/module_data_in[3] scanchain_243/module_data_in[4]
+ scanchain_243/module_data_in[5] scanchain_243/module_data_in[6] scanchain_243/module_data_in[7]
+ scanchain_243/module_data_out[0] scanchain_243/module_data_out[1] scanchain_243/module_data_out[2]
+ scanchain_243/module_data_out[3] scanchain_243/module_data_out[4] scanchain_243/module_data_out[5]
+ scanchain_243/module_data_out[6] scanchain_243/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_232 scanchain_232/module_data_in[0] scanchain_232/module_data_in[1]
+ scanchain_232/module_data_in[2] scanchain_232/module_data_in[3] scanchain_232/module_data_in[4]
+ scanchain_232/module_data_in[5] scanchain_232/module_data_in[6] scanchain_232/module_data_in[7]
+ scanchain_232/module_data_out[0] scanchain_232/module_data_out[1] scanchain_232/module_data_out[2]
+ scanchain_232/module_data_out[3] scanchain_232/module_data_out[4] scanchain_232/module_data_out[5]
+ scanchain_232/module_data_out[6] scanchain_232/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_210 scanchain_210/module_data_in[0] scanchain_210/module_data_in[1]
+ scanchain_210/module_data_in[2] scanchain_210/module_data_in[3] scanchain_210/module_data_in[4]
+ scanchain_210/module_data_in[5] scanchain_210/module_data_in[6] scanchain_210/module_data_in[7]
+ scanchain_210/module_data_out[0] scanchain_210/module_data_out[1] scanchain_210/module_data_out[2]
+ scanchain_210/module_data_out[3] scanchain_210/module_data_out[4] scanchain_210/module_data_out[5]
+ scanchain_210/module_data_out[6] scanchain_210/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_221 scanchain_221/module_data_in[0] scanchain_221/module_data_in[1]
+ scanchain_221/module_data_in[2] scanchain_221/module_data_in[3] scanchain_221/module_data_in[4]
+ scanchain_221/module_data_in[5] scanchain_221/module_data_in[6] scanchain_221/module_data_in[7]
+ scanchain_221/module_data_out[0] scanchain_221/module_data_out[1] scanchain_221/module_data_out[2]
+ scanchain_221/module_data_out[3] scanchain_221/module_data_out[4] scanchain_221/module_data_out[5]
+ scanchain_221/module_data_out[6] scanchain_221/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_349228308755382868_081 scanchain_081/module_data_in[0] scanchain_081/module_data_in[1]
+ scanchain_081/module_data_in[2] scanchain_081/module_data_in[3] scanchain_081/module_data_in[4]
+ scanchain_081/module_data_in[5] scanchain_081/module_data_in[6] scanchain_081/module_data_in[7]
+ scanchain_081/module_data_out[0] scanchain_081/module_data_out[1] scanchain_081/module_data_out[2]
+ scanchain_081/module_data_out[3] scanchain_081/module_data_out[4] scanchain_081/module_data_out[5]
+ scanchain_081/module_data_out[6] scanchain_081/module_data_out[7] vccd1 vssd1 user_module_349228308755382868
Xscanchain_080 scanchain_080/clk_in scanchain_081/clk_in scanchain_080/data_in scanchain_081/data_in
+ scanchain_080/latch_enable_in scanchain_081/latch_enable_in scanchain_080/module_data_in[0]
+ scanchain_080/module_data_in[1] scanchain_080/module_data_in[2] scanchain_080/module_data_in[3]
+ scanchain_080/module_data_in[4] scanchain_080/module_data_in[5] scanchain_080/module_data_in[6]
+ scanchain_080/module_data_in[7] scanchain_080/module_data_out[0] scanchain_080/module_data_out[1]
+ scanchain_080/module_data_out[2] scanchain_080/module_data_out[3] scanchain_080/module_data_out[4]
+ scanchain_080/module_data_out[5] scanchain_080/module_data_out[6] scanchain_080/module_data_out[7]
+ scanchain_080/scan_select_in scanchain_081/scan_select_in vccd1 vssd1 scanchain
Xscanchain_091 scanchain_091/clk_in scanchain_092/clk_in scanchain_091/data_in scanchain_092/data_in
+ scanchain_091/latch_enable_in scanchain_092/latch_enable_in scanchain_091/module_data_in[0]
+ scanchain_091/module_data_in[1] scanchain_091/module_data_in[2] scanchain_091/module_data_in[3]
+ scanchain_091/module_data_in[4] scanchain_091/module_data_in[5] scanchain_091/module_data_in[6]
+ scanchain_091/module_data_in[7] scanchain_091/module_data_out[0] scanchain_091/module_data_out[1]
+ scanchain_091/module_data_out[2] scanchain_091/module_data_out[3] scanchain_091/module_data_out[4]
+ scanchain_091/module_data_out[5] scanchain_091/module_data_out[6] scanchain_091/module_data_out[7]
+ scanchain_091/scan_select_in scanchain_092/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_244 scanchain_244/module_data_in[0] scanchain_244/module_data_in[1]
+ scanchain_244/module_data_in[2] scanchain_244/module_data_in[3] scanchain_244/module_data_in[4]
+ scanchain_244/module_data_in[5] scanchain_244/module_data_in[6] scanchain_244/module_data_in[7]
+ scanchain_244/module_data_out[0] scanchain_244/module_data_out[1] scanchain_244/module_data_out[2]
+ scanchain_244/module_data_out[3] scanchain_244/module_data_out[4] scanchain_244/module_data_out[5]
+ scanchain_244/module_data_out[6] scanchain_244/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_233 scanchain_233/module_data_in[0] scanchain_233/module_data_in[1]
+ scanchain_233/module_data_in[2] scanchain_233/module_data_in[3] scanchain_233/module_data_in[4]
+ scanchain_233/module_data_in[5] scanchain_233/module_data_in[6] scanchain_233/module_data_in[7]
+ scanchain_233/module_data_out[0] scanchain_233/module_data_out[1] scanchain_233/module_data_out[2]
+ scanchain_233/module_data_out[3] scanchain_233/module_data_out[4] scanchain_233/module_data_out[5]
+ scanchain_233/module_data_out[6] scanchain_233/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_222 scanchain_222/module_data_in[0] scanchain_222/module_data_in[1]
+ scanchain_222/module_data_in[2] scanchain_222/module_data_in[3] scanchain_222/module_data_in[4]
+ scanchain_222/module_data_in[5] scanchain_222/module_data_in[6] scanchain_222/module_data_in[7]
+ scanchain_222/module_data_out[0] scanchain_222/module_data_out[1] scanchain_222/module_data_out[2]
+ scanchain_222/module_data_out[3] scanchain_222/module_data_out[4] scanchain_222/module_data_out[5]
+ scanchain_222/module_data_out[6] scanchain_222/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_211 scanchain_211/module_data_in[0] scanchain_211/module_data_in[1]
+ scanchain_211/module_data_in[2] scanchain_211/module_data_in[3] scanchain_211/module_data_in[4]
+ scanchain_211/module_data_in[5] scanchain_211/module_data_in[6] scanchain_211/module_data_in[7]
+ scanchain_211/module_data_out[0] scanchain_211/module_data_out[1] scanchain_211/module_data_out[2]
+ scanchain_211/module_data_out[3] scanchain_211/module_data_out[4] scanchain_211/module_data_out[5]
+ scanchain_211/module_data_out[6] scanchain_211/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_200 scanchain_200/module_data_in[0] scanchain_200/module_data_in[1]
+ scanchain_200/module_data_in[2] scanchain_200/module_data_in[3] scanchain_200/module_data_in[4]
+ scanchain_200/module_data_in[5] scanchain_200/module_data_in[6] scanchain_200/module_data_in[7]
+ scanchain_200/module_data_out[0] scanchain_200/module_data_out[1] scanchain_200/module_data_out[2]
+ scanchain_200/module_data_out[3] scanchain_200/module_data_out[4] scanchain_200/module_data_out[5]
+ scanchain_200/module_data_out[6] scanchain_200/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xmm21_LEDMatrixTop_026 mm21_LEDMatrixTop_026/io_in[0] mm21_LEDMatrixTop_026/io_in[1]
+ mm21_LEDMatrixTop_026/io_in[2] mm21_LEDMatrixTop_026/io_in[3] mm21_LEDMatrixTop_026/io_in[4]
+ mm21_LEDMatrixTop_026/io_in[5] mm21_LEDMatrixTop_026/io_in[6] mm21_LEDMatrixTop_026/io_in[7]
+ mm21_LEDMatrixTop_026/io_out[0] mm21_LEDMatrixTop_026/io_out[1] mm21_LEDMatrixTop_026/io_out[2]
+ mm21_LEDMatrixTop_026/io_out[3] mm21_LEDMatrixTop_026/io_out[4] mm21_LEDMatrixTop_026/io_out[5]
+ mm21_LEDMatrixTop_026/io_out[6] mm21_LEDMatrixTop_026/io_out[7] vccd1 vssd1 mm21_LEDMatrixTop
Xcchan_fp8_multiplier_059 scanchain_059/module_data_in[0] scanchain_059/module_data_in[1]
+ scanchain_059/module_data_in[2] scanchain_059/module_data_in[3] scanchain_059/module_data_in[4]
+ scanchain_059/module_data_in[5] scanchain_059/module_data_in[6] scanchain_059/module_data_in[7]
+ scanchain_059/module_data_out[0] scanchain_059/module_data_out[1] scanchain_059/module_data_out[2]
+ scanchain_059/module_data_out[3] scanchain_059/module_data_out[4] scanchain_059/module_data_out[5]
+ scanchain_059/module_data_out[6] scanchain_059/module_data_out[7] vccd1 vssd1 cchan_fp8_multiplier
Xuser_module_341516949939814994_048 scanchain_048/module_data_in[0] scanchain_048/module_data_in[1]
+ scanchain_048/module_data_in[2] scanchain_048/module_data_in[3] scanchain_048/module_data_in[4]
+ scanchain_048/module_data_in[5] scanchain_048/module_data_in[6] scanchain_048/module_data_in[7]
+ scanchain_048/module_data_out[0] scanchain_048/module_data_out[1] scanchain_048/module_data_out[2]
+ scanchain_048/module_data_out[3] scanchain_048/module_data_out[4] scanchain_048/module_data_out[5]
+ scanchain_048/module_data_out[6] scanchain_048/module_data_out[7] vccd1 vssd1 user_module_341516949939814994
Xuser_module_341535056611770964_096 scanchain_096/module_data_in[0] scanchain_096/module_data_in[1]
+ scanchain_096/module_data_in[2] scanchain_096/module_data_in[3] scanchain_096/module_data_in[4]
+ scanchain_096/module_data_in[5] scanchain_096/module_data_in[6] scanchain_096/module_data_in[7]
+ scanchain_096/module_data_out[0] scanchain_096/module_data_out[1] scanchain_096/module_data_out[2]
+ scanchain_096/module_data_out[3] scanchain_096/module_data_out[4] scanchain_096/module_data_out[5]
+ scanchain_096/module_data_out[6] scanchain_096/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xtholin_avalonsemi_tbb1143_024 scanchain_024/module_data_in[0] scanchain_024/module_data_in[1]
+ scanchain_024/module_data_in[2] scanchain_024/module_data_in[3] scanchain_024/module_data_in[4]
+ scanchain_024/module_data_in[5] scanchain_024/module_data_in[6] scanchain_024/module_data_in[7]
+ scanchain_024/module_data_out[0] scanchain_024/module_data_out[1] scanchain_024/module_data_out[2]
+ scanchain_024/module_data_out[3] scanchain_024/module_data_out[4] scanchain_024/module_data_out[5]
+ scanchain_024/module_data_out[6] scanchain_024/module_data_out[7] vccd1 vssd1 tholin_avalonsemi_tbb1143
Xscanchain_240 scanchain_240/clk_in scanchain_241/clk_in scanchain_240/data_in scanchain_241/data_in
+ scanchain_240/latch_enable_in scanchain_241/latch_enable_in scanchain_240/module_data_in[0]
+ scanchain_240/module_data_in[1] scanchain_240/module_data_in[2] scanchain_240/module_data_in[3]
+ scanchain_240/module_data_in[4] scanchain_240/module_data_in[5] scanchain_240/module_data_in[6]
+ scanchain_240/module_data_in[7] scanchain_240/module_data_out[0] scanchain_240/module_data_out[1]
+ scanchain_240/module_data_out[2] scanchain_240/module_data_out[3] scanchain_240/module_data_out[4]
+ scanchain_240/module_data_out[5] scanchain_240/module_data_out[6] scanchain_240/module_data_out[7]
+ scanchain_240/scan_select_in scanchain_241/scan_select_in vccd1 vssd1 scanchain
Xwren6991_whisk_tt2_io_wrapper_092 scanchain_092/module_data_in[0] scanchain_092/module_data_in[1]
+ scanchain_092/module_data_in[2] scanchain_092/module_data_in[3] scanchain_092/module_data_in[4]
+ scanchain_092/module_data_in[5] scanchain_092/module_data_in[6] scanchain_092/module_data_in[7]
+ scanchain_092/module_data_out[0] scanchain_092/module_data_out[1] scanchain_092/module_data_out[2]
+ scanchain_092/module_data_out[3] scanchain_092/module_data_out[4] scanchain_092/module_data_out[5]
+ scanchain_092/module_data_out[6] scanchain_092/module_data_out[7] vccd1 vssd1 wren6991_whisk_tt2_io_wrapper
Xazdle_binary_clock_009 scanchain_009/module_data_in[0] scanchain_009/module_data_in[1]
+ scanchain_009/module_data_in[2] scanchain_009/module_data_in[3] scanchain_009/module_data_in[4]
+ scanchain_009/module_data_in[5] scanchain_009/module_data_in[6] scanchain_009/module_data_in[7]
+ scanchain_009/module_data_out[0] scanchain_009/module_data_out[1] scanchain_009/module_data_out[2]
+ scanchain_009/module_data_out[3] scanchain_009/module_data_out[4] scanchain_009/module_data_out[5]
+ scanchain_009/module_data_out[6] scanchain_009/module_data_out[7] vccd1 vssd1 azdle_binary_clock
Xscanchain_081 scanchain_081/clk_in scanchain_082/clk_in scanchain_081/data_in scanchain_082/data_in
+ scanchain_081/latch_enable_in scanchain_082/latch_enable_in scanchain_081/module_data_in[0]
+ scanchain_081/module_data_in[1] scanchain_081/module_data_in[2] scanchain_081/module_data_in[3]
+ scanchain_081/module_data_in[4] scanchain_081/module_data_in[5] scanchain_081/module_data_in[6]
+ scanchain_081/module_data_in[7] scanchain_081/module_data_out[0] scanchain_081/module_data_out[1]
+ scanchain_081/module_data_out[2] scanchain_081/module_data_out[3] scanchain_081/module_data_out[4]
+ scanchain_081/module_data_out[5] scanchain_081/module_data_out[6] scanchain_081/module_data_out[7]
+ scanchain_081/scan_select_in scanchain_082/scan_select_in vccd1 vssd1 scanchain
Xscanchain_070 scanchain_070/clk_in scanchain_071/clk_in scanchain_070/data_in scanchain_071/data_in
+ scanchain_070/latch_enable_in scanchain_071/latch_enable_in navray_top_070/io_in[0]
+ navray_top_070/io_in[1] navray_top_070/io_in[2] navray_top_070/io_in[3] navray_top_070/io_in[4]
+ navray_top_070/io_in[5] navray_top_070/io_in[6] navray_top_070/io_in[7] navray_top_070/io_out[0]
+ navray_top_070/io_out[1] navray_top_070/io_out[2] navray_top_070/io_out[3] navray_top_070/io_out[4]
+ navray_top_070/io_out[5] navray_top_070/io_out[6] navray_top_070/io_out[7] scanchain_070/scan_select_in
+ scanchain_071/scan_select_in vccd1 vssd1 scanchain
Xscanchain_092 scanchain_092/clk_in scanchain_093/clk_in scanchain_092/data_in scanchain_093/data_in
+ scanchain_092/latch_enable_in scanchain_093/latch_enable_in scanchain_092/module_data_in[0]
+ scanchain_092/module_data_in[1] scanchain_092/module_data_in[2] scanchain_092/module_data_in[3]
+ scanchain_092/module_data_in[4] scanchain_092/module_data_in[5] scanchain_092/module_data_in[6]
+ scanchain_092/module_data_in[7] scanchain_092/module_data_out[0] scanchain_092/module_data_out[1]
+ scanchain_092/module_data_out[2] scanchain_092/module_data_out[3] scanchain_092/module_data_out[4]
+ scanchain_092/module_data_out[5] scanchain_092/module_data_out[6] scanchain_092/module_data_out[7]
+ scanchain_092/scan_select_in scanchain_093/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_245 scanchain_245/module_data_in[0] scanchain_245/module_data_in[1]
+ scanchain_245/module_data_in[2] scanchain_245/module_data_in[3] scanchain_245/module_data_in[4]
+ scanchain_245/module_data_in[5] scanchain_245/module_data_in[6] scanchain_245/module_data_in[7]
+ scanchain_245/module_data_out[0] scanchain_245/module_data_out[1] scanchain_245/module_data_out[2]
+ scanchain_245/module_data_out[3] scanchain_245/module_data_out[4] scanchain_245/module_data_out[5]
+ scanchain_245/module_data_out[6] scanchain_245/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_234 scanchain_234/module_data_in[0] scanchain_234/module_data_in[1]
+ scanchain_234/module_data_in[2] scanchain_234/module_data_in[3] scanchain_234/module_data_in[4]
+ scanchain_234/module_data_in[5] scanchain_234/module_data_in[6] scanchain_234/module_data_in[7]
+ scanchain_234/module_data_out[0] scanchain_234/module_data_out[1] scanchain_234/module_data_out[2]
+ scanchain_234/module_data_out[3] scanchain_234/module_data_out[4] scanchain_234/module_data_out[5]
+ scanchain_234/module_data_out[6] scanchain_234/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_223 scanchain_223/module_data_in[0] scanchain_223/module_data_in[1]
+ scanchain_223/module_data_in[2] scanchain_223/module_data_in[3] scanchain_223/module_data_in[4]
+ scanchain_223/module_data_in[5] scanchain_223/module_data_in[6] scanchain_223/module_data_in[7]
+ scanchain_223/module_data_out[0] scanchain_223/module_data_out[1] scanchain_223/module_data_out[2]
+ scanchain_223/module_data_out[3] scanchain_223/module_data_out[4] scanchain_223/module_data_out[5]
+ scanchain_223/module_data_out[6] scanchain_223/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_212 scanchain_212/module_data_in[0] scanchain_212/module_data_in[1]
+ scanchain_212/module_data_in[2] scanchain_212/module_data_in[3] scanchain_212/module_data_in[4]
+ scanchain_212/module_data_in[5] scanchain_212/module_data_in[6] scanchain_212/module_data_in[7]
+ scanchain_212/module_data_out[0] scanchain_212/module_data_out[1] scanchain_212/module_data_out[2]
+ scanchain_212/module_data_out[3] scanchain_212/module_data_out[4] scanchain_212/module_data_out[5]
+ scanchain_212/module_data_out[6] scanchain_212/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_201 scanchain_201/module_data_in[0] scanchain_201/module_data_in[1]
+ scanchain_201/module_data_in[2] scanchain_201/module_data_in[3] scanchain_201/module_data_in[4]
+ scanchain_201/module_data_in[5] scanchain_201/module_data_in[6] scanchain_201/module_data_in[7]
+ scanchain_201/module_data_out[0] scanchain_201/module_data_out[1] scanchain_201/module_data_out[2]
+ scanchain_201/module_data_out[3] scanchain_201/module_data_out[4] scanchain_201/module_data_out[5]
+ scanchain_201/module_data_out[6] scanchain_201/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_097 scanchain_097/module_data_in[0] scanchain_097/module_data_in[1]
+ scanchain_097/module_data_in[2] scanchain_097/module_data_in[3] scanchain_097/module_data_in[4]
+ scanchain_097/module_data_in[5] scanchain_097/module_data_in[6] scanchain_097/module_data_in[7]
+ scanchain_097/module_data_out[0] scanchain_097/module_data_out[1] scanchain_097/module_data_out[2]
+ scanchain_097/module_data_out[3] scanchain_097/module_data_out[4] scanchain_097/module_data_out[5]
+ scanchain_097/module_data_out[6] scanchain_097/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_346916357828248146_018 scanchain_018/module_data_in[0] scanchain_018/module_data_in[1]
+ scanchain_018/module_data_in[2] scanchain_018/module_data_in[3] scanchain_018/module_data_in[4]
+ scanchain_018/module_data_in[5] scanchain_018/module_data_in[6] scanchain_018/module_data_in[7]
+ scanchain_018/module_data_out[0] scanchain_018/module_data_out[1] scanchain_018/module_data_out[2]
+ scanchain_018/module_data_out[3] scanchain_018/module_data_out[4] scanchain_018/module_data_out[5]
+ scanchain_018/module_data_out[6] scanchain_018/module_data_out[7] vccd1 vssd1 user_module_346916357828248146
Xscanchain_241 scanchain_241/clk_in scanchain_242/clk_in scanchain_241/data_in scanchain_242/data_in
+ scanchain_241/latch_enable_in scanchain_242/latch_enable_in scanchain_241/module_data_in[0]
+ scanchain_241/module_data_in[1] scanchain_241/module_data_in[2] scanchain_241/module_data_in[3]
+ scanchain_241/module_data_in[4] scanchain_241/module_data_in[5] scanchain_241/module_data_in[6]
+ scanchain_241/module_data_in[7] scanchain_241/module_data_out[0] scanchain_241/module_data_out[1]
+ scanchain_241/module_data_out[2] scanchain_241/module_data_out[3] scanchain_241/module_data_out[4]
+ scanchain_241/module_data_out[5] scanchain_241/module_data_out[6] scanchain_241/module_data_out[7]
+ scanchain_241/scan_select_in scanchain_242/scan_select_in vccd1 vssd1 scanchain
Xscanchain_230 scanchain_230/clk_in scanchain_231/clk_in scanchain_230/data_in scanchain_231/data_in
+ scanchain_230/latch_enable_in scanchain_231/latch_enable_in scanchain_230/module_data_in[0]
+ scanchain_230/module_data_in[1] scanchain_230/module_data_in[2] scanchain_230/module_data_in[3]
+ scanchain_230/module_data_in[4] scanchain_230/module_data_in[5] scanchain_230/module_data_in[6]
+ scanchain_230/module_data_in[7] scanchain_230/module_data_out[0] scanchain_230/module_data_out[1]
+ scanchain_230/module_data_out[2] scanchain_230/module_data_out[3] scanchain_230/module_data_out[4]
+ scanchain_230/module_data_out[5] scanchain_230/module_data_out[6] scanchain_230/module_data_out[7]
+ scanchain_230/scan_select_in scanchain_231/scan_select_in vccd1 vssd1 scanchain
Xscanchain_060 scanchain_060/clk_in scanchain_061/clk_in scanchain_060/data_in scanchain_061/data_in
+ scanchain_060/latch_enable_in scanchain_061/latch_enable_in scanchain_060/module_data_in[0]
+ scanchain_060/module_data_in[1] scanchain_060/module_data_in[2] scanchain_060/module_data_in[3]
+ scanchain_060/module_data_in[4] scanchain_060/module_data_in[5] scanchain_060/module_data_in[6]
+ scanchain_060/module_data_in[7] scanchain_060/module_data_out[0] scanchain_060/module_data_out[1]
+ scanchain_060/module_data_out[2] scanchain_060/module_data_out[3] scanchain_060/module_data_out[4]
+ scanchain_060/module_data_out[5] scanchain_060/module_data_out[6] scanchain_060/module_data_out[7]
+ scanchain_060/scan_select_in scanchain_061/scan_select_in vccd1 vssd1 scanchain
Xscanchain_071 scanchain_071/clk_in scanchain_072/clk_in scanchain_071/data_in scanchain_072/data_in
+ scanchain_071/latch_enable_in scanchain_072/latch_enable_in scanchain_071/module_data_in[0]
+ scanchain_071/module_data_in[1] scanchain_071/module_data_in[2] scanchain_071/module_data_in[3]
+ scanchain_071/module_data_in[4] scanchain_071/module_data_in[5] scanchain_071/module_data_in[6]
+ scanchain_071/module_data_in[7] scanchain_071/module_data_out[0] scanchain_071/module_data_out[1]
+ scanchain_071/module_data_out[2] scanchain_071/module_data_out[3] scanchain_071/module_data_out[4]
+ scanchain_071/module_data_out[5] scanchain_071/module_data_out[6] scanchain_071/module_data_out[7]
+ scanchain_071/scan_select_in scanchain_072/scan_select_in vccd1 vssd1 scanchain
Xscanchain_082 scanchain_082/clk_in scanchain_083/clk_in scanchain_082/data_in scanchain_083/data_in
+ scanchain_082/latch_enable_in scanchain_083/latch_enable_in scanchain_082/module_data_in[0]
+ scanchain_082/module_data_in[1] scanchain_082/module_data_in[2] scanchain_082/module_data_in[3]
+ scanchain_082/module_data_in[4] scanchain_082/module_data_in[5] scanchain_082/module_data_in[6]
+ scanchain_082/module_data_in[7] scanchain_082/module_data_out[0] scanchain_082/module_data_out[1]
+ scanchain_082/module_data_out[2] scanchain_082/module_data_out[3] scanchain_082/module_data_out[4]
+ scanchain_082/module_data_out[5] scanchain_082/module_data_out[6] scanchain_082/module_data_out[7]
+ scanchain_082/scan_select_in scanchain_083/scan_select_in vccd1 vssd1 scanchain
Xscanchain_093 scanchain_093/clk_in scanchain_094/clk_in scanchain_093/data_in scanchain_094/data_in
+ scanchain_093/latch_enable_in scanchain_094/latch_enable_in scanchain_093/module_data_in[0]
+ scanchain_093/module_data_in[1] scanchain_093/module_data_in[2] scanchain_093/module_data_in[3]
+ scanchain_093/module_data_in[4] scanchain_093/module_data_in[5] scanchain_093/module_data_in[6]
+ scanchain_093/module_data_in[7] scanchain_093/module_data_out[0] scanchain_093/module_data_out[1]
+ scanchain_093/module_data_out[2] scanchain_093/module_data_out[3] scanchain_093/module_data_out[4]
+ scanchain_093/module_data_out[5] scanchain_093/module_data_out[6] scanchain_093/module_data_out[7]
+ scanchain_093/scan_select_in scanchain_094/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_246 scanchain_246/module_data_in[0] scanchain_246/module_data_in[1]
+ scanchain_246/module_data_in[2] scanchain_246/module_data_in[3] scanchain_246/module_data_in[4]
+ scanchain_246/module_data_in[5] scanchain_246/module_data_in[6] scanchain_246/module_data_in[7]
+ scanchain_246/module_data_out[0] scanchain_246/module_data_out[1] scanchain_246/module_data_out[2]
+ scanchain_246/module_data_out[3] scanchain_246/module_data_out[4] scanchain_246/module_data_out[5]
+ scanchain_246/module_data_out[6] scanchain_246/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_235 scanchain_235/module_data_in[0] scanchain_235/module_data_in[1]
+ scanchain_235/module_data_in[2] scanchain_235/module_data_in[3] scanchain_235/module_data_in[4]
+ scanchain_235/module_data_in[5] scanchain_235/module_data_in[6] scanchain_235/module_data_in[7]
+ scanchain_235/module_data_out[0] scanchain_235/module_data_out[1] scanchain_235/module_data_out[2]
+ scanchain_235/module_data_out[3] scanchain_235/module_data_out[4] scanchain_235/module_data_out[5]
+ scanchain_235/module_data_out[6] scanchain_235/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_224 scanchain_224/module_data_in[0] scanchain_224/module_data_in[1]
+ scanchain_224/module_data_in[2] scanchain_224/module_data_in[3] scanchain_224/module_data_in[4]
+ scanchain_224/module_data_in[5] scanchain_224/module_data_in[6] scanchain_224/module_data_in[7]
+ scanchain_224/module_data_out[0] scanchain_224/module_data_out[1] scanchain_224/module_data_out[2]
+ scanchain_224/module_data_out[3] scanchain_224/module_data_out[4] scanchain_224/module_data_out[5]
+ scanchain_224/module_data_out[6] scanchain_224/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_213 scanchain_213/module_data_in[0] scanchain_213/module_data_in[1]
+ scanchain_213/module_data_in[2] scanchain_213/module_data_in[3] scanchain_213/module_data_in[4]
+ scanchain_213/module_data_in[5] scanchain_213/module_data_in[6] scanchain_213/module_data_in[7]
+ scanchain_213/module_data_out[0] scanchain_213/module_data_out[1] scanchain_213/module_data_out[2]
+ scanchain_213/module_data_out[3] scanchain_213/module_data_out[4] scanchain_213/module_data_out[5]
+ scanchain_213/module_data_out[6] scanchain_213/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_202 scanchain_202/module_data_in[0] scanchain_202/module_data_in[1]
+ scanchain_202/module_data_in[2] scanchain_202/module_data_in[3] scanchain_202/module_data_in[4]
+ scanchain_202/module_data_in[5] scanchain_202/module_data_in[6] scanchain_202/module_data_in[7]
+ scanchain_202/module_data_out[0] scanchain_202/module_data_out[1] scanchain_202/module_data_out[2]
+ scanchain_202/module_data_out[3] scanchain_202/module_data_out[4] scanchain_202/module_data_out[5]
+ scanchain_202/module_data_out[6] scanchain_202/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_098 scanchain_098/module_data_in[0] scanchain_098/module_data_in[1]
+ scanchain_098/module_data_in[2] scanchain_098/module_data_in[3] scanchain_098/module_data_in[4]
+ scanchain_098/module_data_in[5] scanchain_098/module_data_in[6] scanchain_098/module_data_in[7]
+ scanchain_098/module_data_out[0] scanchain_098/module_data_out[1] scanchain_098/module_data_out[2]
+ scanchain_098/module_data_out[3] scanchain_098/module_data_out[4] scanchain_098/module_data_out[5]
+ scanchain_098/module_data_out[6] scanchain_098/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_242 scanchain_242/clk_in scanchain_243/clk_in scanchain_242/data_in scanchain_243/data_in
+ scanchain_242/latch_enable_in scanchain_243/latch_enable_in scanchain_242/module_data_in[0]
+ scanchain_242/module_data_in[1] scanchain_242/module_data_in[2] scanchain_242/module_data_in[3]
+ scanchain_242/module_data_in[4] scanchain_242/module_data_in[5] scanchain_242/module_data_in[6]
+ scanchain_242/module_data_in[7] scanchain_242/module_data_out[0] scanchain_242/module_data_out[1]
+ scanchain_242/module_data_out[2] scanchain_242/module_data_out[3] scanchain_242/module_data_out[4]
+ scanchain_242/module_data_out[5] scanchain_242/module_data_out[6] scanchain_242/module_data_out[7]
+ scanchain_242/scan_select_in scanchain_243/scan_select_in vccd1 vssd1 scanchain
Xscanchain_231 scanchain_231/clk_in scanchain_232/clk_in scanchain_231/data_in scanchain_232/data_in
+ scanchain_231/latch_enable_in scanchain_232/latch_enable_in scanchain_231/module_data_in[0]
+ scanchain_231/module_data_in[1] scanchain_231/module_data_in[2] scanchain_231/module_data_in[3]
+ scanchain_231/module_data_in[4] scanchain_231/module_data_in[5] scanchain_231/module_data_in[6]
+ scanchain_231/module_data_in[7] scanchain_231/module_data_out[0] scanchain_231/module_data_out[1]
+ scanchain_231/module_data_out[2] scanchain_231/module_data_out[3] scanchain_231/module_data_out[4]
+ scanchain_231/module_data_out[5] scanchain_231/module_data_out[6] scanchain_231/module_data_out[7]
+ scanchain_231/scan_select_in scanchain_232/scan_select_in vccd1 vssd1 scanchain
Xscanchain_220 scanchain_220/clk_in scanchain_221/clk_in scanchain_220/data_in scanchain_221/data_in
+ scanchain_220/latch_enable_in scanchain_221/latch_enable_in scanchain_220/module_data_in[0]
+ scanchain_220/module_data_in[1] scanchain_220/module_data_in[2] scanchain_220/module_data_in[3]
+ scanchain_220/module_data_in[4] scanchain_220/module_data_in[5] scanchain_220/module_data_in[6]
+ scanchain_220/module_data_in[7] scanchain_220/module_data_out[0] scanchain_220/module_data_out[1]
+ scanchain_220/module_data_out[2] scanchain_220/module_data_out[3] scanchain_220/module_data_out[4]
+ scanchain_220/module_data_out[5] scanchain_220/module_data_out[6] scanchain_220/module_data_out[7]
+ scanchain_220/scan_select_in scanchain_221/scan_select_in vccd1 vssd1 scanchain
Xscanchain_050 scanchain_050/clk_in scanchain_051/clk_in scanchain_050/data_in scanchain_051/data_in
+ scanchain_050/latch_enable_in scanchain_051/latch_enable_in scanchain_050/module_data_in[0]
+ scanchain_050/module_data_in[1] scanchain_050/module_data_in[2] scanchain_050/module_data_in[3]
+ scanchain_050/module_data_in[4] scanchain_050/module_data_in[5] scanchain_050/module_data_in[6]
+ scanchain_050/module_data_in[7] scanchain_050/module_data_out[0] scanchain_050/module_data_out[1]
+ scanchain_050/module_data_out[2] scanchain_050/module_data_out[3] scanchain_050/module_data_out[4]
+ scanchain_050/module_data_out[5] scanchain_050/module_data_out[6] scanchain_050/module_data_out[7]
+ scanchain_050/scan_select_in scanchain_051/scan_select_in vccd1 vssd1 scanchain
Xscanchain_061 scanchain_061/clk_in scanchain_062/clk_in scanchain_061/data_in scanchain_062/data_in
+ scanchain_061/latch_enable_in scanchain_062/latch_enable_in scanchain_061/module_data_in[0]
+ scanchain_061/module_data_in[1] scanchain_061/module_data_in[2] scanchain_061/module_data_in[3]
+ scanchain_061/module_data_in[4] scanchain_061/module_data_in[5] scanchain_061/module_data_in[6]
+ scanchain_061/module_data_in[7] scanchain_061/module_data_out[0] scanchain_061/module_data_out[1]
+ scanchain_061/module_data_out[2] scanchain_061/module_data_out[3] scanchain_061/module_data_out[4]
+ scanchain_061/module_data_out[5] scanchain_061/module_data_out[6] scanchain_061/module_data_out[7]
+ scanchain_061/scan_select_in scanchain_062/scan_select_in vccd1 vssd1 scanchain
Xscanchain_072 scanchain_072/clk_in scanchain_073/clk_in scanchain_072/data_in scanchain_073/data_in
+ scanchain_072/latch_enable_in scanchain_073/latch_enable_in scanchain_072/module_data_in[0]
+ scanchain_072/module_data_in[1] scanchain_072/module_data_in[2] scanchain_072/module_data_in[3]
+ scanchain_072/module_data_in[4] scanchain_072/module_data_in[5] scanchain_072/module_data_in[6]
+ scanchain_072/module_data_in[7] scanchain_072/module_data_out[0] scanchain_072/module_data_out[1]
+ scanchain_072/module_data_out[2] scanchain_072/module_data_out[3] scanchain_072/module_data_out[4]
+ scanchain_072/module_data_out[5] scanchain_072/module_data_out[6] scanchain_072/module_data_out[7]
+ scanchain_072/scan_select_in scanchain_073/scan_select_in vccd1 vssd1 scanchain
Xscanchain_083 scanchain_083/clk_in scanchain_084/clk_in scanchain_083/data_in scanchain_084/data_in
+ scanchain_083/latch_enable_in scanchain_084/latch_enable_in scanchain_083/module_data_in[0]
+ scanchain_083/module_data_in[1] scanchain_083/module_data_in[2] scanchain_083/module_data_in[3]
+ scanchain_083/module_data_in[4] scanchain_083/module_data_in[5] scanchain_083/module_data_in[6]
+ scanchain_083/module_data_in[7] scanchain_083/module_data_out[0] scanchain_083/module_data_out[1]
+ scanchain_083/module_data_out[2] scanchain_083/module_data_out[3] scanchain_083/module_data_out[4]
+ scanchain_083/module_data_out[5] scanchain_083/module_data_out[6] scanchain_083/module_data_out[7]
+ scanchain_083/scan_select_in scanchain_084/scan_select_in vccd1 vssd1 scanchain
Xscanchain_094 scanchain_094/clk_in scanchain_095/clk_in scanchain_094/data_in scanchain_095/data_in
+ scanchain_094/latch_enable_in scanchain_095/latch_enable_in scanchain_094/module_data_in[0]
+ scanchain_094/module_data_in[1] scanchain_094/module_data_in[2] scanchain_094/module_data_in[3]
+ scanchain_094/module_data_in[4] scanchain_094/module_data_in[5] scanchain_094/module_data_in[6]
+ scanchain_094/module_data_in[7] scanchain_094/module_data_out[0] scanchain_094/module_data_out[1]
+ scanchain_094/module_data_out[2] scanchain_094/module_data_out[3] scanchain_094/module_data_out[4]
+ scanchain_094/module_data_out[5] scanchain_094/module_data_out[6] scanchain_094/module_data_out[7]
+ scanchain_094/scan_select_in scanchain_095/scan_select_in vccd1 vssd1 scanchain
Xtomkeddie_top_tto_a_025 scanchain_025/module_data_in[0] scanchain_025/module_data_in[1]
+ scanchain_025/module_data_in[2] scanchain_025/module_data_in[3] scanchain_025/module_data_in[4]
+ scanchain_025/module_data_in[5] scanchain_025/module_data_in[6] scanchain_025/module_data_in[7]
+ scanchain_025/module_data_out[0] scanchain_025/module_data_out[1] scanchain_025/module_data_out[2]
+ scanchain_025/module_data_out[3] scanchain_025/module_data_out[4] scanchain_025/module_data_out[5]
+ scanchain_025/module_data_out[6] scanchain_025/module_data_out[7] vccd1 vssd1 tomkeddie_top_tto_a
Xuser_module_341535056611770964_236 scanchain_236/module_data_in[0] scanchain_236/module_data_in[1]
+ scanchain_236/module_data_in[2] scanchain_236/module_data_in[3] scanchain_236/module_data_in[4]
+ scanchain_236/module_data_in[5] scanchain_236/module_data_in[6] scanchain_236/module_data_in[7]
+ scanchain_236/module_data_out[0] scanchain_236/module_data_out[1] scanchain_236/module_data_out[2]
+ scanchain_236/module_data_out[3] scanchain_236/module_data_out[4] scanchain_236/module_data_out[5]
+ scanchain_236/module_data_out[6] scanchain_236/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_247 scanchain_247/module_data_in[0] scanchain_247/module_data_in[1]
+ scanchain_247/module_data_in[2] scanchain_247/module_data_in[3] scanchain_247/module_data_in[4]
+ scanchain_247/module_data_in[5] scanchain_247/module_data_in[6] scanchain_247/module_data_in[7]
+ scanchain_247/module_data_out[0] scanchain_247/module_data_out[1] scanchain_247/module_data_out[2]
+ scanchain_247/module_data_out[3] scanchain_247/module_data_out[4] scanchain_247/module_data_out[5]
+ scanchain_247/module_data_out[6] scanchain_247/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_225 scanchain_225/module_data_in[0] scanchain_225/module_data_in[1]
+ scanchain_225/module_data_in[2] scanchain_225/module_data_in[3] scanchain_225/module_data_in[4]
+ scanchain_225/module_data_in[5] scanchain_225/module_data_in[6] scanchain_225/module_data_in[7]
+ scanchain_225/module_data_out[0] scanchain_225/module_data_out[1] scanchain_225/module_data_out[2]
+ scanchain_225/module_data_out[3] scanchain_225/module_data_out[4] scanchain_225/module_data_out[5]
+ scanchain_225/module_data_out[6] scanchain_225/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_214 scanchain_214/module_data_in[0] scanchain_214/module_data_in[1]
+ scanchain_214/module_data_in[2] scanchain_214/module_data_in[3] scanchain_214/module_data_in[4]
+ scanchain_214/module_data_in[5] scanchain_214/module_data_in[6] scanchain_214/module_data_in[7]
+ scanchain_214/module_data_out[0] scanchain_214/module_data_out[1] scanchain_214/module_data_out[2]
+ scanchain_214/module_data_out[3] scanchain_214/module_data_out[4] scanchain_214/module_data_out[5]
+ scanchain_214/module_data_out[6] scanchain_214/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_203 scanchain_203/module_data_in[0] scanchain_203/module_data_in[1]
+ scanchain_203/module_data_in[2] scanchain_203/module_data_in[3] scanchain_203/module_data_in[4]
+ scanchain_203/module_data_in[5] scanchain_203/module_data_in[6] scanchain_203/module_data_in[7]
+ scanchain_203/module_data_out[0] scanchain_203/module_data_out[1] scanchain_203/module_data_out[2]
+ scanchain_203/module_data_out[3] scanchain_203/module_data_out[4] scanchain_203/module_data_out[5]
+ scanchain_203/module_data_out[6] scanchain_203/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xtiny_fft_015 tiny_fft_015/io_in[0] tiny_fft_015/io_in[1] tiny_fft_015/io_in[2] tiny_fft_015/io_in[3]
+ tiny_fft_015/io_in[4] tiny_fft_015/io_in[5] tiny_fft_015/io_in[6] tiny_fft_015/io_in[7]
+ tiny_fft_015/io_out[0] tiny_fft_015/io_out[1] tiny_fft_015/io_out[2] tiny_fft_015/io_out[3]
+ tiny_fft_015/io_out[4] tiny_fft_015/io_out[5] tiny_fft_015/io_out[6] tiny_fft_015/io_out[7]
+ vccd1 vssd1 tiny_fft
Xrolfmobile99_alu_fsm_top_035 scanchain_035/module_data_in[0] scanchain_035/module_data_in[1]
+ scanchain_035/module_data_in[2] scanchain_035/module_data_in[3] scanchain_035/module_data_in[4]
+ scanchain_035/module_data_in[5] scanchain_035/module_data_in[6] scanchain_035/module_data_in[7]
+ scanchain_035/module_data_out[0] scanchain_035/module_data_out[1] scanchain_035/module_data_out[2]
+ scanchain_035/module_data_out[3] scanchain_035/module_data_out[4] scanchain_035/module_data_out[5]
+ scanchain_035/module_data_out[6] scanchain_035/module_data_out[7] vccd1 vssd1 rolfmobile99_alu_fsm_top
Xuser_module_341535056611770964_000 scanchain_000/module_data_in[0] scanchain_000/module_data_in[1]
+ scanchain_000/module_data_in[2] scanchain_000/module_data_in[3] scanchain_000/module_data_in[4]
+ scanchain_000/module_data_in[5] scanchain_000/module_data_in[6] scanchain_000/module_data_in[7]
+ scanchain_000/module_data_out[0] scanchain_000/module_data_out[1] scanchain_000/module_data_out[2]
+ scanchain_000/module_data_out[3] scanchain_000/module_data_out[4] scanchain_000/module_data_out[5]
+ scanchain_000/module_data_out[6] scanchain_000/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_348260124451668562_034 scanchain_034/module_data_in[0] scanchain_034/module_data_in[1]
+ scanchain_034/module_data_in[2] scanchain_034/module_data_in[3] scanchain_034/module_data_in[4]
+ scanchain_034/module_data_in[5] scanchain_034/module_data_in[6] scanchain_034/module_data_in[7]
+ scanchain_034/module_data_out[0] scanchain_034/module_data_out[1] scanchain_034/module_data_out[2]
+ scanchain_034/module_data_out[3] scanchain_034/module_data_out[4] scanchain_034/module_data_out[5]
+ scanchain_034/module_data_out[6] scanchain_034/module_data_out[7] vccd1 vssd1 user_module_348260124451668562
Xuser_module_341535056611770964_099 scanchain_099/module_data_in[0] scanchain_099/module_data_in[1]
+ scanchain_099/module_data_in[2] scanchain_099/module_data_in[3] scanchain_099/module_data_in[4]
+ scanchain_099/module_data_in[5] scanchain_099/module_data_in[6] scanchain_099/module_data_in[7]
+ scanchain_099/module_data_out[0] scanchain_099/module_data_out[1] scanchain_099/module_data_out[2]
+ scanchain_099/module_data_out[3] scanchain_099/module_data_out[4] scanchain_099/module_data_out[5]
+ scanchain_099/module_data_out[6] scanchain_099/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_243 scanchain_243/clk_in scanchain_244/clk_in scanchain_243/data_in scanchain_244/data_in
+ scanchain_243/latch_enable_in scanchain_244/latch_enable_in scanchain_243/module_data_in[0]
+ scanchain_243/module_data_in[1] scanchain_243/module_data_in[2] scanchain_243/module_data_in[3]
+ scanchain_243/module_data_in[4] scanchain_243/module_data_in[5] scanchain_243/module_data_in[6]
+ scanchain_243/module_data_in[7] scanchain_243/module_data_out[0] scanchain_243/module_data_out[1]
+ scanchain_243/module_data_out[2] scanchain_243/module_data_out[3] scanchain_243/module_data_out[4]
+ scanchain_243/module_data_out[5] scanchain_243/module_data_out[6] scanchain_243/module_data_out[7]
+ scanchain_243/scan_select_in scanchain_244/scan_select_in vccd1 vssd1 scanchain
Xscanchain_232 scanchain_232/clk_in scanchain_233/clk_in scanchain_232/data_in scanchain_233/data_in
+ scanchain_232/latch_enable_in scanchain_233/latch_enable_in scanchain_232/module_data_in[0]
+ scanchain_232/module_data_in[1] scanchain_232/module_data_in[2] scanchain_232/module_data_in[3]
+ scanchain_232/module_data_in[4] scanchain_232/module_data_in[5] scanchain_232/module_data_in[6]
+ scanchain_232/module_data_in[7] scanchain_232/module_data_out[0] scanchain_232/module_data_out[1]
+ scanchain_232/module_data_out[2] scanchain_232/module_data_out[3] scanchain_232/module_data_out[4]
+ scanchain_232/module_data_out[5] scanchain_232/module_data_out[6] scanchain_232/module_data_out[7]
+ scanchain_232/scan_select_in scanchain_233/scan_select_in vccd1 vssd1 scanchain
Xscanchain_210 scanchain_210/clk_in scanchain_211/clk_in scanchain_210/data_in scanchain_211/data_in
+ scanchain_210/latch_enable_in scanchain_211/latch_enable_in scanchain_210/module_data_in[0]
+ scanchain_210/module_data_in[1] scanchain_210/module_data_in[2] scanchain_210/module_data_in[3]
+ scanchain_210/module_data_in[4] scanchain_210/module_data_in[5] scanchain_210/module_data_in[6]
+ scanchain_210/module_data_in[7] scanchain_210/module_data_out[0] scanchain_210/module_data_out[1]
+ scanchain_210/module_data_out[2] scanchain_210/module_data_out[3] scanchain_210/module_data_out[4]
+ scanchain_210/module_data_out[5] scanchain_210/module_data_out[6] scanchain_210/module_data_out[7]
+ scanchain_210/scan_select_in scanchain_211/scan_select_in vccd1 vssd1 scanchain
Xscanchain_221 scanchain_221/clk_in scanchain_222/clk_in scanchain_221/data_in scanchain_222/data_in
+ scanchain_221/latch_enable_in scanchain_222/latch_enable_in scanchain_221/module_data_in[0]
+ scanchain_221/module_data_in[1] scanchain_221/module_data_in[2] scanchain_221/module_data_in[3]
+ scanchain_221/module_data_in[4] scanchain_221/module_data_in[5] scanchain_221/module_data_in[6]
+ scanchain_221/module_data_in[7] scanchain_221/module_data_out[0] scanchain_221/module_data_out[1]
+ scanchain_221/module_data_out[2] scanchain_221/module_data_out[3] scanchain_221/module_data_out[4]
+ scanchain_221/module_data_out[5] scanchain_221/module_data_out[6] scanchain_221/module_data_out[7]
+ scanchain_221/scan_select_in scanchain_222/scan_select_in vccd1 vssd1 scanchain
Xscanchain_051 scanchain_051/clk_in scanchain_052/clk_in scanchain_051/data_in scanchain_052/data_in
+ scanchain_051/latch_enable_in scanchain_052/latch_enable_in scanchain_051/module_data_in[0]
+ scanchain_051/module_data_in[1] scanchain_051/module_data_in[2] scanchain_051/module_data_in[3]
+ scanchain_051/module_data_in[4] scanchain_051/module_data_in[5] scanchain_051/module_data_in[6]
+ scanchain_051/module_data_in[7] scanchain_051/module_data_out[0] scanchain_051/module_data_out[1]
+ scanchain_051/module_data_out[2] scanchain_051/module_data_out[3] scanchain_051/module_data_out[4]
+ scanchain_051/module_data_out[5] scanchain_051/module_data_out[6] scanchain_051/module_data_out[7]
+ scanchain_051/scan_select_in scanchain_052/scan_select_in vccd1 vssd1 scanchain
Xzoechip_031 zoechip_031/io_in[0] zoechip_031/io_in[1] zoechip_031/io_in[2] zoechip_031/io_in[3]
+ zoechip_031/io_in[4] zoechip_031/io_in[5] zoechip_031/io_in[6] zoechip_031/io_in[7]
+ zoechip_031/io_out[0] zoechip_031/io_out[1] zoechip_031/io_out[2] zoechip_031/io_out[3]
+ zoechip_031/io_out[4] zoechip_031/io_out[5] zoechip_031/io_out[6] zoechip_031/io_out[7]
+ vccd1 vssd1 zoechip
Xscanchain_040 scanchain_040/clk_in scanchain_041/clk_in scanchain_040/data_in scanchain_041/data_in
+ scanchain_040/latch_enable_in scanchain_041/latch_enable_in yupferris_bitslam_040/io_in[0]
+ yupferris_bitslam_040/io_in[1] yupferris_bitslam_040/io_in[2] yupferris_bitslam_040/io_in[3]
+ yupferris_bitslam_040/io_in[4] yupferris_bitslam_040/io_in[5] yupferris_bitslam_040/io_in[6]
+ yupferris_bitslam_040/io_in[7] yupferris_bitslam_040/io_out[0] yupferris_bitslam_040/io_out[1]
+ yupferris_bitslam_040/io_out[2] yupferris_bitslam_040/io_out[3] yupferris_bitslam_040/io_out[4]
+ yupferris_bitslam_040/io_out[5] yupferris_bitslam_040/io_out[6] yupferris_bitslam_040/io_out[7]
+ scanchain_040/scan_select_in scanchain_041/scan_select_in vccd1 vssd1 scanchain
Xscanchain_062 scanchain_062/clk_in scanchain_063/clk_in scanchain_062/data_in scanchain_063/data_in
+ scanchain_062/latch_enable_in scanchain_063/latch_enable_in scanchain_062/module_data_in[0]
+ scanchain_062/module_data_in[1] scanchain_062/module_data_in[2] scanchain_062/module_data_in[3]
+ scanchain_062/module_data_in[4] scanchain_062/module_data_in[5] scanchain_062/module_data_in[6]
+ scanchain_062/module_data_in[7] scanchain_062/module_data_out[0] scanchain_062/module_data_out[1]
+ scanchain_062/module_data_out[2] scanchain_062/module_data_out[3] scanchain_062/module_data_out[4]
+ scanchain_062/module_data_out[5] scanchain_062/module_data_out[6] scanchain_062/module_data_out[7]
+ scanchain_062/scan_select_in scanchain_063/scan_select_in vccd1 vssd1 scanchain
Xscanchain_073 scanchain_073/clk_in scanchain_074/clk_in scanchain_073/data_in scanchain_074/data_in
+ scanchain_073/latch_enable_in scanchain_074/latch_enable_in hex_sr_073/io_in[0]
+ hex_sr_073/io_in[1] hex_sr_073/io_in[2] hex_sr_073/io_in[3] hex_sr_073/io_in[4]
+ hex_sr_073/io_in[5] hex_sr_073/io_in[6] hex_sr_073/io_in[7] hex_sr_073/io_out[0]
+ hex_sr_073/io_out[1] hex_sr_073/io_out[2] hex_sr_073/io_out[3] hex_sr_073/io_out[4]
+ hex_sr_073/io_out[5] hex_sr_073/io_out[6] hex_sr_073/io_out[7] scanchain_073/scan_select_in
+ scanchain_074/scan_select_in vccd1 vssd1 scanchain
Xscanchain_084 scanchain_084/clk_in scanchain_085/clk_in scanchain_084/data_in scanchain_085/data_in
+ scanchain_084/latch_enable_in scanchain_085/latch_enable_in moonbase_cpu_8bit_084/io_in[0]
+ moonbase_cpu_8bit_084/io_in[1] moonbase_cpu_8bit_084/io_in[2] moonbase_cpu_8bit_084/io_in[3]
+ moonbase_cpu_8bit_084/io_in[4] moonbase_cpu_8bit_084/io_in[5] moonbase_cpu_8bit_084/io_in[6]
+ moonbase_cpu_8bit_084/io_in[7] moonbase_cpu_8bit_084/io_out[0] moonbase_cpu_8bit_084/io_out[1]
+ moonbase_cpu_8bit_084/io_out[2] moonbase_cpu_8bit_084/io_out[3] moonbase_cpu_8bit_084/io_out[4]
+ moonbase_cpu_8bit_084/io_out[5] moonbase_cpu_8bit_084/io_out[6] moonbase_cpu_8bit_084/io_out[7]
+ scanchain_084/scan_select_in scanchain_085/scan_select_in vccd1 vssd1 scanchain
Xscanchain_095 scanchain_095/clk_in scanchain_096/clk_in scanchain_095/data_in scanchain_096/data_in
+ scanchain_095/latch_enable_in scanchain_096/latch_enable_in scanchain_095/module_data_in[0]
+ scanchain_095/module_data_in[1] scanchain_095/module_data_in[2] scanchain_095/module_data_in[3]
+ scanchain_095/module_data_in[4] scanchain_095/module_data_in[5] scanchain_095/module_data_in[6]
+ scanchain_095/module_data_in[7] scanchain_095/module_data_out[0] scanchain_095/module_data_out[1]
+ scanchain_095/module_data_out[2] scanchain_095/module_data_out[3] scanchain_095/module_data_out[4]
+ scanchain_095/module_data_out[5] scanchain_095/module_data_out[6] scanchain_095/module_data_out[7]
+ scanchain_095/scan_select_in scanchain_096/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_237 scanchain_237/module_data_in[0] scanchain_237/module_data_in[1]
+ scanchain_237/module_data_in[2] scanchain_237/module_data_in[3] scanchain_237/module_data_in[4]
+ scanchain_237/module_data_in[5] scanchain_237/module_data_in[6] scanchain_237/module_data_in[7]
+ scanchain_237/module_data_out[0] scanchain_237/module_data_out[1] scanchain_237/module_data_out[2]
+ scanchain_237/module_data_out[3] scanchain_237/module_data_out[4] scanchain_237/module_data_out[5]
+ scanchain_237/module_data_out[6] scanchain_237/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_248 scanchain_248/module_data_in[0] scanchain_248/module_data_in[1]
+ scanchain_248/module_data_in[2] scanchain_248/module_data_in[3] scanchain_248/module_data_in[4]
+ scanchain_248/module_data_in[5] scanchain_248/module_data_in[6] scanchain_248/module_data_in[7]
+ scanchain_248/module_data_out[0] scanchain_248/module_data_out[1] scanchain_248/module_data_out[2]
+ scanchain_248/module_data_out[3] scanchain_248/module_data_out[4] scanchain_248/module_data_out[5]
+ scanchain_248/module_data_out[6] scanchain_248/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_226 scanchain_226/module_data_in[0] scanchain_226/module_data_in[1]
+ scanchain_226/module_data_in[2] scanchain_226/module_data_in[3] scanchain_226/module_data_in[4]
+ scanchain_226/module_data_in[5] scanchain_226/module_data_in[6] scanchain_226/module_data_in[7]
+ scanchain_226/module_data_out[0] scanchain_226/module_data_out[1] scanchain_226/module_data_out[2]
+ scanchain_226/module_data_out[3] scanchain_226/module_data_out[4] scanchain_226/module_data_out[5]
+ scanchain_226/module_data_out[6] scanchain_226/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_215 scanchain_215/module_data_in[0] scanchain_215/module_data_in[1]
+ scanchain_215/module_data_in[2] scanchain_215/module_data_in[3] scanchain_215/module_data_in[4]
+ scanchain_215/module_data_in[5] scanchain_215/module_data_in[6] scanchain_215/module_data_in[7]
+ scanchain_215/module_data_out[0] scanchain_215/module_data_out[1] scanchain_215/module_data_out[2]
+ scanchain_215/module_data_out[3] scanchain_215/module_data_out[4] scanchain_215/module_data_out[5]
+ scanchain_215/module_data_out[6] scanchain_215/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_204 scanchain_204/module_data_in[0] scanchain_204/module_data_in[1]
+ scanchain_204/module_data_in[2] scanchain_204/module_data_in[3] scanchain_204/module_data_in[4]
+ scanchain_204/module_data_in[5] scanchain_204/module_data_in[6] scanchain_204/module_data_in[7]
+ scanchain_204/module_data_out[0] scanchain_204/module_data_out[1] scanchain_204/module_data_out[2]
+ scanchain_204/module_data_out[3] scanchain_204/module_data_out[4] scanchain_204/module_data_out[5]
+ scanchain_204/module_data_out[6] scanchain_204/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_244 scanchain_244/clk_in scanchain_245/clk_in scanchain_244/data_in scanchain_245/data_in
+ scanchain_244/latch_enable_in scanchain_245/latch_enable_in scanchain_244/module_data_in[0]
+ scanchain_244/module_data_in[1] scanchain_244/module_data_in[2] scanchain_244/module_data_in[3]
+ scanchain_244/module_data_in[4] scanchain_244/module_data_in[5] scanchain_244/module_data_in[6]
+ scanchain_244/module_data_in[7] scanchain_244/module_data_out[0] scanchain_244/module_data_out[1]
+ scanchain_244/module_data_out[2] scanchain_244/module_data_out[3] scanchain_244/module_data_out[4]
+ scanchain_244/module_data_out[5] scanchain_244/module_data_out[6] scanchain_244/module_data_out[7]
+ scanchain_244/scan_select_in scanchain_245/scan_select_in vccd1 vssd1 scanchain
Xscanchain_233 scanchain_233/clk_in scanchain_234/clk_in scanchain_233/data_in scanchain_234/data_in
+ scanchain_233/latch_enable_in scanchain_234/latch_enable_in scanchain_233/module_data_in[0]
+ scanchain_233/module_data_in[1] scanchain_233/module_data_in[2] scanchain_233/module_data_in[3]
+ scanchain_233/module_data_in[4] scanchain_233/module_data_in[5] scanchain_233/module_data_in[6]
+ scanchain_233/module_data_in[7] scanchain_233/module_data_out[0] scanchain_233/module_data_out[1]
+ scanchain_233/module_data_out[2] scanchain_233/module_data_out[3] scanchain_233/module_data_out[4]
+ scanchain_233/module_data_out[5] scanchain_233/module_data_out[6] scanchain_233/module_data_out[7]
+ scanchain_233/scan_select_in scanchain_234/scan_select_in vccd1 vssd1 scanchain
Xscanchain_222 scanchain_222/clk_in scanchain_223/clk_in scanchain_222/data_in scanchain_223/data_in
+ scanchain_222/latch_enable_in scanchain_223/latch_enable_in scanchain_222/module_data_in[0]
+ scanchain_222/module_data_in[1] scanchain_222/module_data_in[2] scanchain_222/module_data_in[3]
+ scanchain_222/module_data_in[4] scanchain_222/module_data_in[5] scanchain_222/module_data_in[6]
+ scanchain_222/module_data_in[7] scanchain_222/module_data_out[0] scanchain_222/module_data_out[1]
+ scanchain_222/module_data_out[2] scanchain_222/module_data_out[3] scanchain_222/module_data_out[4]
+ scanchain_222/module_data_out[5] scanchain_222/module_data_out[6] scanchain_222/module_data_out[7]
+ scanchain_222/scan_select_in scanchain_223/scan_select_in vccd1 vssd1 scanchain
Xscanchain_211 scanchain_211/clk_in scanchain_212/clk_in scanchain_211/data_in scanchain_212/data_in
+ scanchain_211/latch_enable_in scanchain_212/latch_enable_in scanchain_211/module_data_in[0]
+ scanchain_211/module_data_in[1] scanchain_211/module_data_in[2] scanchain_211/module_data_in[3]
+ scanchain_211/module_data_in[4] scanchain_211/module_data_in[5] scanchain_211/module_data_in[6]
+ scanchain_211/module_data_in[7] scanchain_211/module_data_out[0] scanchain_211/module_data_out[1]
+ scanchain_211/module_data_out[2] scanchain_211/module_data_out[3] scanchain_211/module_data_out[4]
+ scanchain_211/module_data_out[5] scanchain_211/module_data_out[6] scanchain_211/module_data_out[7]
+ scanchain_211/scan_select_in scanchain_212/scan_select_in vccd1 vssd1 scanchain
Xscanchain_200 scanchain_200/clk_in scanchain_201/clk_in scanchain_200/data_in scanchain_201/data_in
+ scanchain_200/latch_enable_in scanchain_201/latch_enable_in scanchain_200/module_data_in[0]
+ scanchain_200/module_data_in[1] scanchain_200/module_data_in[2] scanchain_200/module_data_in[3]
+ scanchain_200/module_data_in[4] scanchain_200/module_data_in[5] scanchain_200/module_data_in[6]
+ scanchain_200/module_data_in[7] scanchain_200/module_data_out[0] scanchain_200/module_data_out[1]
+ scanchain_200/module_data_out[2] scanchain_200/module_data_out[3] scanchain_200/module_data_out[4]
+ scanchain_200/module_data_out[5] scanchain_200/module_data_out[6] scanchain_200/module_data_out[7]
+ scanchain_200/scan_select_in scanchain_201/scan_select_in vccd1 vssd1 scanchain
Xxyz_peppergray_Potato1_top_030 scanchain_030/module_data_in[0] scanchain_030/module_data_in[1]
+ scanchain_030/module_data_in[2] scanchain_030/module_data_in[3] scanchain_030/module_data_in[4]
+ scanchain_030/module_data_in[5] scanchain_030/module_data_in[6] scanchain_030/module_data_in[7]
+ scanchain_030/module_data_out[0] scanchain_030/module_data_out[1] scanchain_030/module_data_out[2]
+ scanchain_030/module_data_out[3] scanchain_030/module_data_out[4] scanchain_030/module_data_out[5]
+ scanchain_030/module_data_out[6] scanchain_030/module_data_out[7] vccd1 vssd1 xyz_peppergray_Potato1_top
Xscanchain_030 scanchain_030/clk_in scanchain_031/clk_in scanchain_030/data_in scanchain_031/data_in
+ scanchain_030/latch_enable_in scanchain_031/latch_enable_in scanchain_030/module_data_in[0]
+ scanchain_030/module_data_in[1] scanchain_030/module_data_in[2] scanchain_030/module_data_in[3]
+ scanchain_030/module_data_in[4] scanchain_030/module_data_in[5] scanchain_030/module_data_in[6]
+ scanchain_030/module_data_in[7] scanchain_030/module_data_out[0] scanchain_030/module_data_out[1]
+ scanchain_030/module_data_out[2] scanchain_030/module_data_out[3] scanchain_030/module_data_out[4]
+ scanchain_030/module_data_out[5] scanchain_030/module_data_out[6] scanchain_030/module_data_out[7]
+ scanchain_030/scan_select_in scanchain_031/scan_select_in vccd1 vssd1 scanchain
Xscanchain_041 scanchain_041/clk_in scanchain_042/clk_in scanchain_041/data_in scanchain_042/data_in
+ scanchain_041/latch_enable_in scanchain_042/latch_enable_in scanchain_041/module_data_in[0]
+ scanchain_041/module_data_in[1] scanchain_041/module_data_in[2] scanchain_041/module_data_in[3]
+ scanchain_041/module_data_in[4] scanchain_041/module_data_in[5] scanchain_041/module_data_in[6]
+ scanchain_041/module_data_in[7] scanchain_041/module_data_out[0] scanchain_041/module_data_out[1]
+ scanchain_041/module_data_out[2] scanchain_041/module_data_out[3] scanchain_041/module_data_out[4]
+ scanchain_041/module_data_out[5] scanchain_041/module_data_out[6] scanchain_041/module_data_out[7]
+ scanchain_041/scan_select_in scanchain_042/scan_select_in vccd1 vssd1 scanchain
Xscanchain_052 scanchain_052/clk_in scanchain_053/clk_in scanchain_052/data_in scanchain_053/data_in
+ scanchain_052/latch_enable_in scanchain_053/latch_enable_in scanchain_052/module_data_in[0]
+ scanchain_052/module_data_in[1] scanchain_052/module_data_in[2] scanchain_052/module_data_in[3]
+ scanchain_052/module_data_in[4] scanchain_052/module_data_in[5] scanchain_052/module_data_in[6]
+ scanchain_052/module_data_in[7] scanchain_052/module_data_out[0] scanchain_052/module_data_out[1]
+ scanchain_052/module_data_out[2] scanchain_052/module_data_out[3] scanchain_052/module_data_out[4]
+ scanchain_052/module_data_out[5] scanchain_052/module_data_out[6] scanchain_052/module_data_out[7]
+ scanchain_052/scan_select_in scanchain_053/scan_select_in vccd1 vssd1 scanchain
Xscanchain_063 scanchain_063/clk_in scanchain_064/clk_in scanchain_063/data_in scanchain_064/data_in
+ scanchain_063/latch_enable_in scanchain_064/latch_enable_in scanchain_063/module_data_in[0]
+ scanchain_063/module_data_in[1] scanchain_063/module_data_in[2] scanchain_063/module_data_in[3]
+ scanchain_063/module_data_in[4] scanchain_063/module_data_in[5] scanchain_063/module_data_in[6]
+ scanchain_063/module_data_in[7] scanchain_063/module_data_out[0] scanchain_063/module_data_out[1]
+ scanchain_063/module_data_out[2] scanchain_063/module_data_out[3] scanchain_063/module_data_out[4]
+ scanchain_063/module_data_out[5] scanchain_063/module_data_out[6] scanchain_063/module_data_out[7]
+ scanchain_063/scan_select_in scanchain_064/scan_select_in vccd1 vssd1 scanchain
Xscanchain_074 scanchain_074/clk_in scanchain_075/clk_in scanchain_074/data_in scanchain_075/data_in
+ scanchain_074/latch_enable_in scanchain_075/latch_enable_in scanchain_074/module_data_in[0]
+ scanchain_074/module_data_in[1] scanchain_074/module_data_in[2] scanchain_074/module_data_in[3]
+ scanchain_074/module_data_in[4] scanchain_074/module_data_in[5] scanchain_074/module_data_in[6]
+ scanchain_074/module_data_in[7] scanchain_074/module_data_out[0] scanchain_074/module_data_out[1]
+ scanchain_074/module_data_out[2] scanchain_074/module_data_out[3] scanchain_074/module_data_out[4]
+ scanchain_074/module_data_out[5] scanchain_074/module_data_out[6] scanchain_074/module_data_out[7]
+ scanchain_074/scan_select_in scanchain_075/scan_select_in vccd1 vssd1 scanchain
Xscanchain_085 scanchain_085/clk_in scanchain_086/clk_in scanchain_085/data_in scanchain_086/data_in
+ scanchain_085/latch_enable_in scanchain_086/latch_enable_in scanchain_085/module_data_in[0]
+ scanchain_085/module_data_in[1] scanchain_085/module_data_in[2] scanchain_085/module_data_in[3]
+ scanchain_085/module_data_in[4] scanchain_085/module_data_in[5] scanchain_085/module_data_in[6]
+ scanchain_085/module_data_in[7] scanchain_085/module_data_out[0] scanchain_085/module_data_out[1]
+ scanchain_085/module_data_out[2] scanchain_085/module_data_out[3] scanchain_085/module_data_out[4]
+ scanchain_085/module_data_out[5] scanchain_085/module_data_out[6] scanchain_085/module_data_out[7]
+ scanchain_085/scan_select_in scanchain_086/scan_select_in vccd1 vssd1 scanchain
Xscanchain_096 scanchain_096/clk_in scanchain_097/clk_in scanchain_096/data_in scanchain_097/data_in
+ scanchain_096/latch_enable_in scanchain_097/latch_enable_in scanchain_096/module_data_in[0]
+ scanchain_096/module_data_in[1] scanchain_096/module_data_in[2] scanchain_096/module_data_in[3]
+ scanchain_096/module_data_in[4] scanchain_096/module_data_in[5] scanchain_096/module_data_in[6]
+ scanchain_096/module_data_in[7] scanchain_096/module_data_out[0] scanchain_096/module_data_out[1]
+ scanchain_096/module_data_out[2] scanchain_096/module_data_out[3] scanchain_096/module_data_out[4]
+ scanchain_096/module_data_out[5] scanchain_096/module_data_out[6] scanchain_096/module_data_out[7]
+ scanchain_096/scan_select_in scanchain_097/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_238 scanchain_238/module_data_in[0] scanchain_238/module_data_in[1]
+ scanchain_238/module_data_in[2] scanchain_238/module_data_in[3] scanchain_238/module_data_in[4]
+ scanchain_238/module_data_in[5] scanchain_238/module_data_in[6] scanchain_238/module_data_in[7]
+ scanchain_238/module_data_out[0] scanchain_238/module_data_out[1] scanchain_238/module_data_out[2]
+ scanchain_238/module_data_out[3] scanchain_238/module_data_out[4] scanchain_238/module_data_out[5]
+ scanchain_238/module_data_out[6] scanchain_238/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_249 scanchain_249/module_data_in[0] scanchain_249/module_data_in[1]
+ scanchain_249/module_data_in[2] scanchain_249/module_data_in[3] scanchain_249/module_data_in[4]
+ scanchain_249/module_data_in[5] scanchain_249/module_data_in[6] scanchain_249/module_data_in[7]
+ scanchain_249/module_data_out[0] scanchain_249/module_data_out[1] scanchain_249/module_data_out[2]
+ scanchain_249/module_data_out[3] scanchain_249/module_data_out[4] scanchain_249/module_data_out[5]
+ scanchain_249/module_data_out[6] scanchain_249/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_227 scanchain_227/module_data_in[0] scanchain_227/module_data_in[1]
+ scanchain_227/module_data_in[2] scanchain_227/module_data_in[3] scanchain_227/module_data_in[4]
+ scanchain_227/module_data_in[5] scanchain_227/module_data_in[6] scanchain_227/module_data_in[7]
+ scanchain_227/module_data_out[0] scanchain_227/module_data_out[1] scanchain_227/module_data_out[2]
+ scanchain_227/module_data_out[3] scanchain_227/module_data_out[4] scanchain_227/module_data_out[5]
+ scanchain_227/module_data_out[6] scanchain_227/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_216 scanchain_216/module_data_in[0] scanchain_216/module_data_in[1]
+ scanchain_216/module_data_in[2] scanchain_216/module_data_in[3] scanchain_216/module_data_in[4]
+ scanchain_216/module_data_in[5] scanchain_216/module_data_in[6] scanchain_216/module_data_in[7]
+ scanchain_216/module_data_out[0] scanchain_216/module_data_out[1] scanchain_216/module_data_out[2]
+ scanchain_216/module_data_out[3] scanchain_216/module_data_out[4] scanchain_216/module_data_out[5]
+ scanchain_216/module_data_out[6] scanchain_216/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_205 scanchain_205/module_data_in[0] scanchain_205/module_data_in[1]
+ scanchain_205/module_data_in[2] scanchain_205/module_data_in[3] scanchain_205/module_data_in[4]
+ scanchain_205/module_data_in[5] scanchain_205/module_data_in[6] scanchain_205/module_data_in[7]
+ scanchain_205/module_data_out[0] scanchain_205/module_data_out[1] scanchain_205/module_data_out[2]
+ scanchain_205/module_data_out[3] scanchain_205/module_data_out[4] scanchain_205/module_data_out[5]
+ scanchain_205/module_data_out[6] scanchain_205/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_245 scanchain_245/clk_in scanchain_246/clk_in scanchain_245/data_in scanchain_246/data_in
+ scanchain_245/latch_enable_in scanchain_246/latch_enable_in scanchain_245/module_data_in[0]
+ scanchain_245/module_data_in[1] scanchain_245/module_data_in[2] scanchain_245/module_data_in[3]
+ scanchain_245/module_data_in[4] scanchain_245/module_data_in[5] scanchain_245/module_data_in[6]
+ scanchain_245/module_data_in[7] scanchain_245/module_data_out[0] scanchain_245/module_data_out[1]
+ scanchain_245/module_data_out[2] scanchain_245/module_data_out[3] scanchain_245/module_data_out[4]
+ scanchain_245/module_data_out[5] scanchain_245/module_data_out[6] scanchain_245/module_data_out[7]
+ scanchain_245/scan_select_in scanchain_246/scan_select_in vccd1 vssd1 scanchain
Xscanchain_234 scanchain_234/clk_in scanchain_235/clk_in scanchain_234/data_in scanchain_235/data_in
+ scanchain_234/latch_enable_in scanchain_235/latch_enable_in scanchain_234/module_data_in[0]
+ scanchain_234/module_data_in[1] scanchain_234/module_data_in[2] scanchain_234/module_data_in[3]
+ scanchain_234/module_data_in[4] scanchain_234/module_data_in[5] scanchain_234/module_data_in[6]
+ scanchain_234/module_data_in[7] scanchain_234/module_data_out[0] scanchain_234/module_data_out[1]
+ scanchain_234/module_data_out[2] scanchain_234/module_data_out[3] scanchain_234/module_data_out[4]
+ scanchain_234/module_data_out[5] scanchain_234/module_data_out[6] scanchain_234/module_data_out[7]
+ scanchain_234/scan_select_in scanchain_235/scan_select_in vccd1 vssd1 scanchain
Xscanchain_223 scanchain_223/clk_in scanchain_224/clk_in scanchain_223/data_in scanchain_224/data_in
+ scanchain_223/latch_enable_in scanchain_224/latch_enable_in scanchain_223/module_data_in[0]
+ scanchain_223/module_data_in[1] scanchain_223/module_data_in[2] scanchain_223/module_data_in[3]
+ scanchain_223/module_data_in[4] scanchain_223/module_data_in[5] scanchain_223/module_data_in[6]
+ scanchain_223/module_data_in[7] scanchain_223/module_data_out[0] scanchain_223/module_data_out[1]
+ scanchain_223/module_data_out[2] scanchain_223/module_data_out[3] scanchain_223/module_data_out[4]
+ scanchain_223/module_data_out[5] scanchain_223/module_data_out[6] scanchain_223/module_data_out[7]
+ scanchain_223/scan_select_in scanchain_224/scan_select_in vccd1 vssd1 scanchain
Xscanchain_212 scanchain_212/clk_in scanchain_213/clk_in scanchain_212/data_in scanchain_213/data_in
+ scanchain_212/latch_enable_in scanchain_213/latch_enable_in scanchain_212/module_data_in[0]
+ scanchain_212/module_data_in[1] scanchain_212/module_data_in[2] scanchain_212/module_data_in[3]
+ scanchain_212/module_data_in[4] scanchain_212/module_data_in[5] scanchain_212/module_data_in[6]
+ scanchain_212/module_data_in[7] scanchain_212/module_data_out[0] scanchain_212/module_data_out[1]
+ scanchain_212/module_data_out[2] scanchain_212/module_data_out[3] scanchain_212/module_data_out[4]
+ scanchain_212/module_data_out[5] scanchain_212/module_data_out[6] scanchain_212/module_data_out[7]
+ scanchain_212/scan_select_in scanchain_213/scan_select_in vccd1 vssd1 scanchain
Xscanchain_201 scanchain_201/clk_in scanchain_202/clk_in scanchain_201/data_in scanchain_202/data_in
+ scanchain_201/latch_enable_in scanchain_202/latch_enable_in scanchain_201/module_data_in[0]
+ scanchain_201/module_data_in[1] scanchain_201/module_data_in[2] scanchain_201/module_data_in[3]
+ scanchain_201/module_data_in[4] scanchain_201/module_data_in[5] scanchain_201/module_data_in[6]
+ scanchain_201/module_data_in[7] scanchain_201/module_data_out[0] scanchain_201/module_data_out[1]
+ scanchain_201/module_data_out[2] scanchain_201/module_data_out[3] scanchain_201/module_data_out[4]
+ scanchain_201/module_data_out[5] scanchain_201/module_data_out[6] scanchain_201/module_data_out[7]
+ scanchain_201/scan_select_in scanchain_202/scan_select_in vccd1 vssd1 scanchain
Xhex_sr_073 hex_sr_073/io_in[0] hex_sr_073/io_in[1] hex_sr_073/io_in[2] hex_sr_073/io_in[3]
+ hex_sr_073/io_in[4] hex_sr_073/io_in[5] hex_sr_073/io_in[6] hex_sr_073/io_in[7]
+ hex_sr_073/io_out[0] hex_sr_073/io_out[1] hex_sr_073/io_out[2] hex_sr_073/io_out[3]
+ hex_sr_073/io_out[4] hex_sr_073/io_out[5] hex_sr_073/io_out[6] hex_sr_073/io_out[7]
+ vccd1 vssd1 hex_sr
Xuser_module_341277789473735250_094 scanchain_094/module_data_in[0] scanchain_094/module_data_in[1]
+ scanchain_094/module_data_in[2] scanchain_094/module_data_in[3] scanchain_094/module_data_in[4]
+ scanchain_094/module_data_in[5] scanchain_094/module_data_in[6] scanchain_094/module_data_in[7]
+ scanchain_094/module_data_out[0] scanchain_094/module_data_out[1] scanchain_094/module_data_out[2]
+ scanchain_094/module_data_out[3] scanchain_094/module_data_out[4] scanchain_094/module_data_out[5]
+ scanchain_094/module_data_out[6] scanchain_094/module_data_out[7] vccd1 vssd1 user_module_341277789473735250
Xscanchain_053 scanchain_053/clk_in scanchain_054/clk_in scanchain_053/data_in scanchain_054/data_in
+ scanchain_053/latch_enable_in scanchain_054/latch_enable_in xor_shift32_evango_053/io_in[0]
+ xor_shift32_evango_053/io_in[1] xor_shift32_evango_053/io_in[2] xor_shift32_evango_053/io_in[3]
+ xor_shift32_evango_053/io_in[4] xor_shift32_evango_053/io_in[5] xor_shift32_evango_053/io_in[6]
+ xor_shift32_evango_053/io_in[7] xor_shift32_evango_053/io_out[0] xor_shift32_evango_053/io_out[1]
+ xor_shift32_evango_053/io_out[2] xor_shift32_evango_053/io_out[3] xor_shift32_evango_053/io_out[4]
+ xor_shift32_evango_053/io_out[5] xor_shift32_evango_053/io_out[6] xor_shift32_evango_053/io_out[7]
+ scanchain_053/scan_select_in scanchain_054/scan_select_in vccd1 vssd1 scanchain
Xscanchain_031 scanchain_031/clk_in scanchain_032/clk_in scanchain_031/data_in scanchain_032/data_in
+ scanchain_031/latch_enable_in scanchain_032/latch_enable_in zoechip_031/io_in[0]
+ zoechip_031/io_in[1] zoechip_031/io_in[2] zoechip_031/io_in[3] zoechip_031/io_in[4]
+ zoechip_031/io_in[5] zoechip_031/io_in[6] zoechip_031/io_in[7] zoechip_031/io_out[0]
+ zoechip_031/io_out[1] zoechip_031/io_out[2] zoechip_031/io_out[3] zoechip_031/io_out[4]
+ zoechip_031/io_out[5] zoechip_031/io_out[6] zoechip_031/io_out[7] scanchain_031/scan_select_in
+ scanchain_032/scan_select_in vccd1 vssd1 scanchain
Xscanchain_020 scanchain_020/clk_in scanchain_021/clk_in scanchain_020/data_in scanchain_021/data_in
+ scanchain_020/latch_enable_in scanchain_021/latch_enable_in chase_the_beat_020/io_in[0]
+ chase_the_beat_020/io_in[1] chase_the_beat_020/io_in[2] chase_the_beat_020/io_in[3]
+ chase_the_beat_020/io_in[4] chase_the_beat_020/io_in[5] chase_the_beat_020/io_in[6]
+ chase_the_beat_020/io_in[7] chase_the_beat_020/io_out[0] chase_the_beat_020/io_out[1]
+ chase_the_beat_020/io_out[2] chase_the_beat_020/io_out[3] chase_the_beat_020/io_out[4]
+ chase_the_beat_020/io_out[5] chase_the_beat_020/io_out[6] chase_the_beat_020/io_out[7]
+ scanchain_020/scan_select_in scanchain_021/scan_select_in vccd1 vssd1 scanchain
Xscanchain_042 scanchain_042/clk_in scanchain_043/clk_in scanchain_042/data_in scanchain_043/data_in
+ scanchain_042/latch_enable_in scanchain_043/latch_enable_in scanchain_042/module_data_in[0]
+ scanchain_042/module_data_in[1] scanchain_042/module_data_in[2] scanchain_042/module_data_in[3]
+ scanchain_042/module_data_in[4] scanchain_042/module_data_in[5] scanchain_042/module_data_in[6]
+ scanchain_042/module_data_in[7] scanchain_042/module_data_out[0] scanchain_042/module_data_out[1]
+ scanchain_042/module_data_out[2] scanchain_042/module_data_out[3] scanchain_042/module_data_out[4]
+ scanchain_042/module_data_out[5] scanchain_042/module_data_out[6] scanchain_042/module_data_out[7]
+ scanchain_042/scan_select_in scanchain_043/scan_select_in vccd1 vssd1 scanchain
Xscanchain_064 scanchain_064/clk_in scanchain_065/clk_in scanchain_064/data_in scanchain_065/data_in
+ scanchain_064/latch_enable_in scanchain_065/latch_enable_in scanchain_064/module_data_in[0]
+ scanchain_064/module_data_in[1] scanchain_064/module_data_in[2] scanchain_064/module_data_in[3]
+ scanchain_064/module_data_in[4] scanchain_064/module_data_in[5] scanchain_064/module_data_in[6]
+ scanchain_064/module_data_in[7] scanchain_064/module_data_out[0] scanchain_064/module_data_out[1]
+ scanchain_064/module_data_out[2] scanchain_064/module_data_out[3] scanchain_064/module_data_out[4]
+ scanchain_064/module_data_out[5] scanchain_064/module_data_out[6] scanchain_064/module_data_out[7]
+ scanchain_064/scan_select_in scanchain_065/scan_select_in vccd1 vssd1 scanchain
Xscanchain_075 scanchain_075/clk_in scanchain_076/clk_in scanchain_075/data_in scanchain_076/data_in
+ scanchain_075/latch_enable_in scanchain_076/latch_enable_in scanchain_075/module_data_in[0]
+ scanchain_075/module_data_in[1] scanchain_075/module_data_in[2] scanchain_075/module_data_in[3]
+ scanchain_075/module_data_in[4] scanchain_075/module_data_in[5] scanchain_075/module_data_in[6]
+ scanchain_075/module_data_in[7] scanchain_075/module_data_out[0] scanchain_075/module_data_out[1]
+ scanchain_075/module_data_out[2] scanchain_075/module_data_out[3] scanchain_075/module_data_out[4]
+ scanchain_075/module_data_out[5] scanchain_075/module_data_out[6] scanchain_075/module_data_out[7]
+ scanchain_075/scan_select_in scanchain_076/scan_select_in vccd1 vssd1 scanchain
Xscanchain_086 scanchain_086/clk_in scanchain_087/clk_in scanchain_086/data_in scanchain_087/data_in
+ scanchain_086/latch_enable_in scanchain_087/latch_enable_in scanchain_086/module_data_in[0]
+ scanchain_086/module_data_in[1] scanchain_086/module_data_in[2] scanchain_086/module_data_in[3]
+ scanchain_086/module_data_in[4] scanchain_086/module_data_in[5] scanchain_086/module_data_in[6]
+ scanchain_086/module_data_in[7] scanchain_086/module_data_out[0] scanchain_086/module_data_out[1]
+ scanchain_086/module_data_out[2] scanchain_086/module_data_out[3] scanchain_086/module_data_out[4]
+ scanchain_086/module_data_out[5] scanchain_086/module_data_out[6] scanchain_086/module_data_out[7]
+ scanchain_086/scan_select_in scanchain_087/scan_select_in vccd1 vssd1 scanchain
Xscanchain_097 scanchain_097/clk_in scanchain_098/clk_in scanchain_097/data_in scanchain_098/data_in
+ scanchain_097/latch_enable_in scanchain_098/latch_enable_in scanchain_097/module_data_in[0]
+ scanchain_097/module_data_in[1] scanchain_097/module_data_in[2] scanchain_097/module_data_in[3]
+ scanchain_097/module_data_in[4] scanchain_097/module_data_in[5] scanchain_097/module_data_in[6]
+ scanchain_097/module_data_in[7] scanchain_097/module_data_out[0] scanchain_097/module_data_out[1]
+ scanchain_097/module_data_out[2] scanchain_097/module_data_out[3] scanchain_097/module_data_out[4]
+ scanchain_097/module_data_out[5] scanchain_097/module_data_out[6] scanchain_097/module_data_out[7]
+ scanchain_097/scan_select_in scanchain_098/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_239 scanchain_239/module_data_in[0] scanchain_239/module_data_in[1]
+ scanchain_239/module_data_in[2] scanchain_239/module_data_in[3] scanchain_239/module_data_in[4]
+ scanchain_239/module_data_in[5] scanchain_239/module_data_in[6] scanchain_239/module_data_in[7]
+ scanchain_239/module_data_out[0] scanchain_239/module_data_out[1] scanchain_239/module_data_out[2]
+ scanchain_239/module_data_out[3] scanchain_239/module_data_out[4] scanchain_239/module_data_out[5]
+ scanchain_239/module_data_out[6] scanchain_239/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_228 scanchain_228/module_data_in[0] scanchain_228/module_data_in[1]
+ scanchain_228/module_data_in[2] scanchain_228/module_data_in[3] scanchain_228/module_data_in[4]
+ scanchain_228/module_data_in[5] scanchain_228/module_data_in[6] scanchain_228/module_data_in[7]
+ scanchain_228/module_data_out[0] scanchain_228/module_data_out[1] scanchain_228/module_data_out[2]
+ scanchain_228/module_data_out[3] scanchain_228/module_data_out[4] scanchain_228/module_data_out[5]
+ scanchain_228/module_data_out[6] scanchain_228/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_217 scanchain_217/module_data_in[0] scanchain_217/module_data_in[1]
+ scanchain_217/module_data_in[2] scanchain_217/module_data_in[3] scanchain_217/module_data_in[4]
+ scanchain_217/module_data_in[5] scanchain_217/module_data_in[6] scanchain_217/module_data_in[7]
+ scanchain_217/module_data_out[0] scanchain_217/module_data_out[1] scanchain_217/module_data_out[2]
+ scanchain_217/module_data_out[3] scanchain_217/module_data_out[4] scanchain_217/module_data_out[5]
+ scanchain_217/module_data_out[6] scanchain_217/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_206 scanchain_206/module_data_in[0] scanchain_206/module_data_in[1]
+ scanchain_206/module_data_in[2] scanchain_206/module_data_in[3] scanchain_206/module_data_in[4]
+ scanchain_206/module_data_in[5] scanchain_206/module_data_in[6] scanchain_206/module_data_in[7]
+ scanchain_206/module_data_out[0] scanchain_206/module_data_out[1] scanchain_206/module_data_out[2]
+ scanchain_206/module_data_out[3] scanchain_206/module_data_out[4] scanchain_206/module_data_out[5]
+ scanchain_206/module_data_out[6] scanchain_206/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_246 scanchain_246/clk_in scanchain_247/clk_in scanchain_246/data_in scanchain_247/data_in
+ scanchain_246/latch_enable_in scanchain_247/latch_enable_in scanchain_246/module_data_in[0]
+ scanchain_246/module_data_in[1] scanchain_246/module_data_in[2] scanchain_246/module_data_in[3]
+ scanchain_246/module_data_in[4] scanchain_246/module_data_in[5] scanchain_246/module_data_in[6]
+ scanchain_246/module_data_in[7] scanchain_246/module_data_out[0] scanchain_246/module_data_out[1]
+ scanchain_246/module_data_out[2] scanchain_246/module_data_out[3] scanchain_246/module_data_out[4]
+ scanchain_246/module_data_out[5] scanchain_246/module_data_out[6] scanchain_246/module_data_out[7]
+ scanchain_246/scan_select_in scanchain_247/scan_select_in vccd1 vssd1 scanchain
Xscanchain_235 scanchain_235/clk_in scanchain_236/clk_in scanchain_235/data_in scanchain_236/data_in
+ scanchain_235/latch_enable_in scanchain_236/latch_enable_in scanchain_235/module_data_in[0]
+ scanchain_235/module_data_in[1] scanchain_235/module_data_in[2] scanchain_235/module_data_in[3]
+ scanchain_235/module_data_in[4] scanchain_235/module_data_in[5] scanchain_235/module_data_in[6]
+ scanchain_235/module_data_in[7] scanchain_235/module_data_out[0] scanchain_235/module_data_out[1]
+ scanchain_235/module_data_out[2] scanchain_235/module_data_out[3] scanchain_235/module_data_out[4]
+ scanchain_235/module_data_out[5] scanchain_235/module_data_out[6] scanchain_235/module_data_out[7]
+ scanchain_235/scan_select_in scanchain_236/scan_select_in vccd1 vssd1 scanchain
Xscanchain_224 scanchain_224/clk_in scanchain_225/clk_in scanchain_224/data_in scanchain_225/data_in
+ scanchain_224/latch_enable_in scanchain_225/latch_enable_in scanchain_224/module_data_in[0]
+ scanchain_224/module_data_in[1] scanchain_224/module_data_in[2] scanchain_224/module_data_in[3]
+ scanchain_224/module_data_in[4] scanchain_224/module_data_in[5] scanchain_224/module_data_in[6]
+ scanchain_224/module_data_in[7] scanchain_224/module_data_out[0] scanchain_224/module_data_out[1]
+ scanchain_224/module_data_out[2] scanchain_224/module_data_out[3] scanchain_224/module_data_out[4]
+ scanchain_224/module_data_out[5] scanchain_224/module_data_out[6] scanchain_224/module_data_out[7]
+ scanchain_224/scan_select_in scanchain_225/scan_select_in vccd1 vssd1 scanchain
Xscanchain_213 scanchain_213/clk_in scanchain_214/clk_in scanchain_213/data_in scanchain_214/data_in
+ scanchain_213/latch_enable_in scanchain_214/latch_enable_in scanchain_213/module_data_in[0]
+ scanchain_213/module_data_in[1] scanchain_213/module_data_in[2] scanchain_213/module_data_in[3]
+ scanchain_213/module_data_in[4] scanchain_213/module_data_in[5] scanchain_213/module_data_in[6]
+ scanchain_213/module_data_in[7] scanchain_213/module_data_out[0] scanchain_213/module_data_out[1]
+ scanchain_213/module_data_out[2] scanchain_213/module_data_out[3] scanchain_213/module_data_out[4]
+ scanchain_213/module_data_out[5] scanchain_213/module_data_out[6] scanchain_213/module_data_out[7]
+ scanchain_213/scan_select_in scanchain_214/scan_select_in vccd1 vssd1 scanchain
Xscanchain_202 scanchain_202/clk_in scanchain_203/clk_in scanchain_202/data_in scanchain_203/data_in
+ scanchain_202/latch_enable_in scanchain_203/latch_enable_in scanchain_202/module_data_in[0]
+ scanchain_202/module_data_in[1] scanchain_202/module_data_in[2] scanchain_202/module_data_in[3]
+ scanchain_202/module_data_in[4] scanchain_202/module_data_in[5] scanchain_202/module_data_in[6]
+ scanchain_202/module_data_in[7] scanchain_202/module_data_out[0] scanchain_202/module_data_out[1]
+ scanchain_202/module_data_out[2] scanchain_202/module_data_out[3] scanchain_202/module_data_out[4]
+ scanchain_202/module_data_out[5] scanchain_202/module_data_out[6] scanchain_202/module_data_out[7]
+ scanchain_202/scan_select_in scanchain_203/scan_select_in vccd1 vssd1 scanchain
Xscanchain_032 scanchain_032/clk_in scanchain_033/clk_in scanchain_032/data_in scanchain_033/data_in
+ scanchain_032/latch_enable_in scanchain_033/latch_enable_in scanchain_032/module_data_in[0]
+ scanchain_032/module_data_in[1] scanchain_032/module_data_in[2] scanchain_032/module_data_in[3]
+ scanchain_032/module_data_in[4] scanchain_032/module_data_in[5] scanchain_032/module_data_in[6]
+ scanchain_032/module_data_in[7] scanchain_032/module_data_out[0] scanchain_032/module_data_out[1]
+ scanchain_032/module_data_out[2] scanchain_032/module_data_out[3] scanchain_032/module_data_out[4]
+ scanchain_032/module_data_out[5] scanchain_032/module_data_out[6] scanchain_032/module_data_out[7]
+ scanchain_032/scan_select_in scanchain_033/scan_select_in vccd1 vssd1 scanchain
Xscanchain_021 scanchain_021/clk_in scanchain_022/clk_in scanchain_021/data_in scanchain_022/data_in
+ scanchain_021/latch_enable_in scanchain_022/latch_enable_in scanchain_021/module_data_in[0]
+ scanchain_021/module_data_in[1] scanchain_021/module_data_in[2] scanchain_021/module_data_in[3]
+ scanchain_021/module_data_in[4] scanchain_021/module_data_in[5] scanchain_021/module_data_in[6]
+ scanchain_021/module_data_in[7] scanchain_021/module_data_out[0] scanchain_021/module_data_out[1]
+ scanchain_021/module_data_out[2] scanchain_021/module_data_out[3] scanchain_021/module_data_out[4]
+ scanchain_021/module_data_out[5] scanchain_021/module_data_out[6] scanchain_021/module_data_out[7]
+ scanchain_021/scan_select_in scanchain_022/scan_select_in vccd1 vssd1 scanchain
Xscanchain_010 scanchain_010/clk_in scanchain_011/clk_in scanchain_010/data_in scanchain_011/data_in
+ scanchain_010/latch_enable_in scanchain_011/latch_enable_in scanchain_010/module_data_in[0]
+ scanchain_010/module_data_in[1] scanchain_010/module_data_in[2] scanchain_010/module_data_in[3]
+ scanchain_010/module_data_in[4] scanchain_010/module_data_in[5] scanchain_010/module_data_in[6]
+ scanchain_010/module_data_in[7] scanchain_010/module_data_out[0] scanchain_010/module_data_out[1]
+ scanchain_010/module_data_out[2] scanchain_010/module_data_out[3] scanchain_010/module_data_out[4]
+ scanchain_010/module_data_out[5] scanchain_010/module_data_out[6] scanchain_010/module_data_out[7]
+ scanchain_010/scan_select_in scanchain_011/scan_select_in vccd1 vssd1 scanchain
Xscanchain_043 scanchain_043/clk_in scanchain_044/clk_in scanchain_043/data_in scanchain_044/data_in
+ scanchain_043/latch_enable_in scanchain_044/latch_enable_in rc5_top_043/io_in[0]
+ rc5_top_043/io_in[1] rc5_top_043/io_in[2] rc5_top_043/io_in[3] rc5_top_043/io_in[4]
+ rc5_top_043/io_in[5] rc5_top_043/io_in[6] rc5_top_043/io_in[7] rc5_top_043/io_out[0]
+ rc5_top_043/io_out[1] rc5_top_043/io_out[2] rc5_top_043/io_out[3] rc5_top_043/io_out[4]
+ rc5_top_043/io_out[5] rc5_top_043/io_out[6] rc5_top_043/io_out[7] scanchain_043/scan_select_in
+ scanchain_044/scan_select_in vccd1 vssd1 scanchain
Xscanchain_054 scanchain_054/clk_in scanchain_055/clk_in scanchain_054/data_in scanchain_055/data_in
+ scanchain_054/latch_enable_in scanchain_055/latch_enable_in scanchain_054/module_data_in[0]
+ scanchain_054/module_data_in[1] scanchain_054/module_data_in[2] scanchain_054/module_data_in[3]
+ scanchain_054/module_data_in[4] scanchain_054/module_data_in[5] scanchain_054/module_data_in[6]
+ scanchain_054/module_data_in[7] scanchain_054/module_data_out[0] scanchain_054/module_data_out[1]
+ scanchain_054/module_data_out[2] scanchain_054/module_data_out[3] scanchain_054/module_data_out[4]
+ scanchain_054/module_data_out[5] scanchain_054/module_data_out[6] scanchain_054/module_data_out[7]
+ scanchain_054/scan_select_in scanchain_055/scan_select_in vccd1 vssd1 scanchain
Xscanchain_065 scanchain_065/clk_in scanchain_066/clk_in scanchain_065/data_in scanchain_066/data_in
+ scanchain_065/latch_enable_in scanchain_066/latch_enable_in scanchain_065/module_data_in[0]
+ scanchain_065/module_data_in[1] scanchain_065/module_data_in[2] scanchain_065/module_data_in[3]
+ scanchain_065/module_data_in[4] scanchain_065/module_data_in[5] scanchain_065/module_data_in[6]
+ scanchain_065/module_data_in[7] scanchain_065/module_data_out[0] scanchain_065/module_data_out[1]
+ scanchain_065/module_data_out[2] scanchain_065/module_data_out[3] scanchain_065/module_data_out[4]
+ scanchain_065/module_data_out[5] scanchain_065/module_data_out[6] scanchain_065/module_data_out[7]
+ scanchain_065/scan_select_in scanchain_066/scan_select_in vccd1 vssd1 scanchain
Xscanchain_076 scanchain_076/clk_in scanchain_077/clk_in scanchain_076/data_in scanchain_077/data_in
+ scanchain_076/latch_enable_in scanchain_077/latch_enable_in scanchain_076/module_data_in[0]
+ scanchain_076/module_data_in[1] scanchain_076/module_data_in[2] scanchain_076/module_data_in[3]
+ scanchain_076/module_data_in[4] scanchain_076/module_data_in[5] scanchain_076/module_data_in[6]
+ scanchain_076/module_data_in[7] scanchain_076/module_data_out[0] scanchain_076/module_data_out[1]
+ scanchain_076/module_data_out[2] scanchain_076/module_data_out[3] scanchain_076/module_data_out[4]
+ scanchain_076/module_data_out[5] scanchain_076/module_data_out[6] scanchain_076/module_data_out[7]
+ scanchain_076/scan_select_in scanchain_077/scan_select_in vccd1 vssd1 scanchain
Xscanchain_087 scanchain_087/clk_in scanchain_088/clk_in scanchain_087/data_in scanchain_088/data_in
+ scanchain_087/latch_enable_in scanchain_088/latch_enable_in scanchain_087/module_data_in[0]
+ scanchain_087/module_data_in[1] scanchain_087/module_data_in[2] scanchain_087/module_data_in[3]
+ scanchain_087/module_data_in[4] scanchain_087/module_data_in[5] scanchain_087/module_data_in[6]
+ scanchain_087/module_data_in[7] scanchain_087/module_data_out[0] scanchain_087/module_data_out[1]
+ scanchain_087/module_data_out[2] scanchain_087/module_data_out[3] scanchain_087/module_data_out[4]
+ scanchain_087/module_data_out[5] scanchain_087/module_data_out[6] scanchain_087/module_data_out[7]
+ scanchain_087/scan_select_in scanchain_088/scan_select_in vccd1 vssd1 scanchain
Xscanchain_098 scanchain_098/clk_in scanchain_099/clk_in scanchain_098/data_in scanchain_099/data_in
+ scanchain_098/latch_enable_in scanchain_099/latch_enable_in scanchain_098/module_data_in[0]
+ scanchain_098/module_data_in[1] scanchain_098/module_data_in[2] scanchain_098/module_data_in[3]
+ scanchain_098/module_data_in[4] scanchain_098/module_data_in[5] scanchain_098/module_data_in[6]
+ scanchain_098/module_data_in[7] scanchain_098/module_data_out[0] scanchain_098/module_data_out[1]
+ scanchain_098/module_data_out[2] scanchain_098/module_data_out[3] scanchain_098/module_data_out[4]
+ scanchain_098/module_data_out[5] scanchain_098/module_data_out[6] scanchain_098/module_data_out[7]
+ scanchain_098/scan_select_in scanchain_099/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_229 scanchain_229/module_data_in[0] scanchain_229/module_data_in[1]
+ scanchain_229/module_data_in[2] scanchain_229/module_data_in[3] scanchain_229/module_data_in[4]
+ scanchain_229/module_data_in[5] scanchain_229/module_data_in[6] scanchain_229/module_data_in[7]
+ scanchain_229/module_data_out[0] scanchain_229/module_data_out[1] scanchain_229/module_data_out[2]
+ scanchain_229/module_data_out[3] scanchain_229/module_data_out[4] scanchain_229/module_data_out[5]
+ scanchain_229/module_data_out[6] scanchain_229/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_218 scanchain_218/module_data_in[0] scanchain_218/module_data_in[1]
+ scanchain_218/module_data_in[2] scanchain_218/module_data_in[3] scanchain_218/module_data_in[4]
+ scanchain_218/module_data_in[5] scanchain_218/module_data_in[6] scanchain_218/module_data_in[7]
+ scanchain_218/module_data_out[0] scanchain_218/module_data_out[1] scanchain_218/module_data_out[2]
+ scanchain_218/module_data_out[3] scanchain_218/module_data_out[4] scanchain_218/module_data_out[5]
+ scanchain_218/module_data_out[6] scanchain_218/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_207 scanchain_207/module_data_in[0] scanchain_207/module_data_in[1]
+ scanchain_207/module_data_in[2] scanchain_207/module_data_in[3] scanchain_207/module_data_in[4]
+ scanchain_207/module_data_in[5] scanchain_207/module_data_in[6] scanchain_207/module_data_in[7]
+ scanchain_207/module_data_out[0] scanchain_207/module_data_out[1] scanchain_207/module_data_out[2]
+ scanchain_207/module_data_out[3] scanchain_207/module_data_out[4] scanchain_207/module_data_out[5]
+ scanchain_207/module_data_out[6] scanchain_207/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_236 scanchain_236/clk_in scanchain_237/clk_in scanchain_236/data_in scanchain_237/data_in
+ scanchain_236/latch_enable_in scanchain_237/latch_enable_in scanchain_236/module_data_in[0]
+ scanchain_236/module_data_in[1] scanchain_236/module_data_in[2] scanchain_236/module_data_in[3]
+ scanchain_236/module_data_in[4] scanchain_236/module_data_in[5] scanchain_236/module_data_in[6]
+ scanchain_236/module_data_in[7] scanchain_236/module_data_out[0] scanchain_236/module_data_out[1]
+ scanchain_236/module_data_out[2] scanchain_236/module_data_out[3] scanchain_236/module_data_out[4]
+ scanchain_236/module_data_out[5] scanchain_236/module_data_out[6] scanchain_236/module_data_out[7]
+ scanchain_236/scan_select_in scanchain_237/scan_select_in vccd1 vssd1 scanchain
Xscanchain_247 scanchain_247/clk_in scanchain_248/clk_in scanchain_247/data_in scanchain_248/data_in
+ scanchain_247/latch_enable_in scanchain_248/latch_enable_in scanchain_247/module_data_in[0]
+ scanchain_247/module_data_in[1] scanchain_247/module_data_in[2] scanchain_247/module_data_in[3]
+ scanchain_247/module_data_in[4] scanchain_247/module_data_in[5] scanchain_247/module_data_in[6]
+ scanchain_247/module_data_in[7] scanchain_247/module_data_out[0] scanchain_247/module_data_out[1]
+ scanchain_247/module_data_out[2] scanchain_247/module_data_out[3] scanchain_247/module_data_out[4]
+ scanchain_247/module_data_out[5] scanchain_247/module_data_out[6] scanchain_247/module_data_out[7]
+ scanchain_247/scan_select_in scanchain_248/scan_select_in vccd1 vssd1 scanchain
Xscanchain_225 scanchain_225/clk_in scanchain_226/clk_in scanchain_225/data_in scanchain_226/data_in
+ scanchain_225/latch_enable_in scanchain_226/latch_enable_in scanchain_225/module_data_in[0]
+ scanchain_225/module_data_in[1] scanchain_225/module_data_in[2] scanchain_225/module_data_in[3]
+ scanchain_225/module_data_in[4] scanchain_225/module_data_in[5] scanchain_225/module_data_in[6]
+ scanchain_225/module_data_in[7] scanchain_225/module_data_out[0] scanchain_225/module_data_out[1]
+ scanchain_225/module_data_out[2] scanchain_225/module_data_out[3] scanchain_225/module_data_out[4]
+ scanchain_225/module_data_out[5] scanchain_225/module_data_out[6] scanchain_225/module_data_out[7]
+ scanchain_225/scan_select_in scanchain_226/scan_select_in vccd1 vssd1 scanchain
Xscanchain_214 scanchain_214/clk_in scanchain_215/clk_in scanchain_214/data_in scanchain_215/data_in
+ scanchain_214/latch_enable_in scanchain_215/latch_enable_in scanchain_214/module_data_in[0]
+ scanchain_214/module_data_in[1] scanchain_214/module_data_in[2] scanchain_214/module_data_in[3]
+ scanchain_214/module_data_in[4] scanchain_214/module_data_in[5] scanchain_214/module_data_in[6]
+ scanchain_214/module_data_in[7] scanchain_214/module_data_out[0] scanchain_214/module_data_out[1]
+ scanchain_214/module_data_out[2] scanchain_214/module_data_out[3] scanchain_214/module_data_out[4]
+ scanchain_214/module_data_out[5] scanchain_214/module_data_out[6] scanchain_214/module_data_out[7]
+ scanchain_214/scan_select_in scanchain_215/scan_select_in vccd1 vssd1 scanchain
Xscanchain_203 scanchain_203/clk_in scanchain_204/clk_in scanchain_203/data_in scanchain_204/data_in
+ scanchain_203/latch_enable_in scanchain_204/latch_enable_in scanchain_203/module_data_in[0]
+ scanchain_203/module_data_in[1] scanchain_203/module_data_in[2] scanchain_203/module_data_in[3]
+ scanchain_203/module_data_in[4] scanchain_203/module_data_in[5] scanchain_203/module_data_in[6]
+ scanchain_203/module_data_in[7] scanchain_203/module_data_out[0] scanchain_203/module_data_out[1]
+ scanchain_203/module_data_out[2] scanchain_203/module_data_out[3] scanchain_203/module_data_out[4]
+ scanchain_203/module_data_out[5] scanchain_203/module_data_out[6] scanchain_203/module_data_out[7]
+ scanchain_203/scan_select_in scanchain_204/scan_select_in vccd1 vssd1 scanchain
Xscanchain_033 scanchain_033/clk_in scanchain_034/clk_in scanchain_033/data_in scanchain_034/data_in
+ scanchain_033/latch_enable_in scanchain_034/latch_enable_in mbikovitsky_top_033/io_in[0]
+ mbikovitsky_top_033/io_in[1] mbikovitsky_top_033/io_in[2] mbikovitsky_top_033/io_in[3]
+ mbikovitsky_top_033/io_in[4] mbikovitsky_top_033/io_in[5] mbikovitsky_top_033/io_in[6]
+ mbikovitsky_top_033/io_in[7] mbikovitsky_top_033/io_out[0] mbikovitsky_top_033/io_out[1]
+ mbikovitsky_top_033/io_out[2] mbikovitsky_top_033/io_out[3] mbikovitsky_top_033/io_out[4]
+ mbikovitsky_top_033/io_out[5] mbikovitsky_top_033/io_out[6] mbikovitsky_top_033/io_out[7]
+ scanchain_033/scan_select_in scanchain_034/scan_select_in vccd1 vssd1 scanchain
Xscanchain_022 scanchain_022/clk_in scanchain_023/clk_in scanchain_022/data_in scanchain_023/data_in
+ scanchain_022/latch_enable_in scanchain_023/latch_enable_in scanchain_022/module_data_in[0]
+ scanchain_022/module_data_in[1] scanchain_022/module_data_in[2] scanchain_022/module_data_in[3]
+ scanchain_022/module_data_in[4] scanchain_022/module_data_in[5] scanchain_022/module_data_in[6]
+ scanchain_022/module_data_in[7] scanchain_022/module_data_out[0] scanchain_022/module_data_out[1]
+ scanchain_022/module_data_out[2] scanchain_022/module_data_out[3] scanchain_022/module_data_out[4]
+ scanchain_022/module_data_out[5] scanchain_022/module_data_out[6] scanchain_022/module_data_out[7]
+ scanchain_022/scan_select_in scanchain_023/scan_select_in vccd1 vssd1 scanchain
Xscanchain_011 scanchain_011/clk_in scanchain_012/clk_in scanchain_011/data_in scanchain_012/data_in
+ scanchain_011/latch_enable_in scanchain_012/latch_enable_in jar_sram_top_011/io_in[0]
+ jar_sram_top_011/io_in[1] jar_sram_top_011/io_in[2] jar_sram_top_011/io_in[3] jar_sram_top_011/io_in[4]
+ jar_sram_top_011/io_in[5] jar_sram_top_011/io_in[6] jar_sram_top_011/io_in[7] jar_sram_top_011/io_out[0]
+ jar_sram_top_011/io_out[1] jar_sram_top_011/io_out[2] jar_sram_top_011/io_out[3]
+ jar_sram_top_011/io_out[4] jar_sram_top_011/io_out[5] jar_sram_top_011/io_out[6]
+ jar_sram_top_011/io_out[7] scanchain_011/scan_select_in scanchain_012/scan_select_in
+ vccd1 vssd1 scanchain
Xscanchain_000 scanchain_000/clk_in scanchain_001/clk_in scanchain_000/data_in scanchain_001/data_in
+ scanchain_000/latch_enable_in scanchain_001/latch_enable_in scanchain_000/module_data_in[0]
+ scanchain_000/module_data_in[1] scanchain_000/module_data_in[2] scanchain_000/module_data_in[3]
+ scanchain_000/module_data_in[4] scanchain_000/module_data_in[5] scanchain_000/module_data_in[6]
+ scanchain_000/module_data_in[7] scanchain_000/module_data_out[0] scanchain_000/module_data_out[1]
+ scanchain_000/module_data_out[2] scanchain_000/module_data_out[3] scanchain_000/module_data_out[4]
+ scanchain_000/module_data_out[5] scanchain_000/module_data_out[6] scanchain_000/module_data_out[7]
+ scan_controller/scan_select scanchain_001/scan_select_in vccd1 vssd1 scanchain
Xscanchain_044 scanchain_044/clk_in scanchain_045/clk_in scanchain_044/data_in scanchain_045/data_in
+ scanchain_044/latch_enable_in scanchain_045/latch_enable_in scanchain_044/module_data_in[0]
+ scanchain_044/module_data_in[1] scanchain_044/module_data_in[2] scanchain_044/module_data_in[3]
+ scanchain_044/module_data_in[4] scanchain_044/module_data_in[5] scanchain_044/module_data_in[6]
+ scanchain_044/module_data_in[7] scanchain_044/module_data_out[0] scanchain_044/module_data_out[1]
+ scanchain_044/module_data_out[2] scanchain_044/module_data_out[3] scanchain_044/module_data_out[4]
+ scanchain_044/module_data_out[5] scanchain_044/module_data_out[6] scanchain_044/module_data_out[7]
+ scanchain_044/scan_select_in scanchain_045/scan_select_in vccd1 vssd1 scanchain
Xscanchain_055 scanchain_055/clk_in scanchain_056/clk_in scanchain_055/data_in scanchain_056/data_in
+ scanchain_055/latch_enable_in scanchain_056/latch_enable_in scanchain_055/module_data_in[0]
+ scanchain_055/module_data_in[1] scanchain_055/module_data_in[2] scanchain_055/module_data_in[3]
+ scanchain_055/module_data_in[4] scanchain_055/module_data_in[5] scanchain_055/module_data_in[6]
+ scanchain_055/module_data_in[7] scanchain_055/module_data_out[0] scanchain_055/module_data_out[1]
+ scanchain_055/module_data_out[2] scanchain_055/module_data_out[3] scanchain_055/module_data_out[4]
+ scanchain_055/module_data_out[5] scanchain_055/module_data_out[6] scanchain_055/module_data_out[7]
+ scanchain_055/scan_select_in scanchain_056/scan_select_in vccd1 vssd1 scanchain
Xscanchain_066 scanchain_066/clk_in scanchain_067/clk_in scanchain_066/data_in scanchain_067/data_in
+ scanchain_066/latch_enable_in scanchain_067/latch_enable_in udxs_sqrt_top_066/io_in[0]
+ udxs_sqrt_top_066/io_in[1] udxs_sqrt_top_066/io_in[2] udxs_sqrt_top_066/io_in[3]
+ udxs_sqrt_top_066/io_in[4] udxs_sqrt_top_066/io_in[5] udxs_sqrt_top_066/io_in[6]
+ udxs_sqrt_top_066/io_in[7] udxs_sqrt_top_066/io_out[0] udxs_sqrt_top_066/io_out[1]
+ udxs_sqrt_top_066/io_out[2] udxs_sqrt_top_066/io_out[3] udxs_sqrt_top_066/io_out[4]
+ udxs_sqrt_top_066/io_out[5] udxs_sqrt_top_066/io_out[6] udxs_sqrt_top_066/io_out[7]
+ scanchain_066/scan_select_in scanchain_067/scan_select_in vccd1 vssd1 scanchain
Xscanchain_077 scanchain_077/clk_in scanchain_078/clk_in scanchain_077/data_in scanchain_078/data_in
+ scanchain_077/latch_enable_in scanchain_078/latch_enable_in cpldcpu_MCPU5plus_077/io_in[0]
+ cpldcpu_MCPU5plus_077/io_in[1] cpldcpu_MCPU5plus_077/io_in[2] cpldcpu_MCPU5plus_077/io_in[3]
+ cpldcpu_MCPU5plus_077/io_in[4] cpldcpu_MCPU5plus_077/io_in[5] cpldcpu_MCPU5plus_077/io_in[6]
+ cpldcpu_MCPU5plus_077/io_in[7] cpldcpu_MCPU5plus_077/io_out[0] cpldcpu_MCPU5plus_077/io_out[1]
+ cpldcpu_MCPU5plus_077/io_out[2] cpldcpu_MCPU5plus_077/io_out[3] cpldcpu_MCPU5plus_077/io_out[4]
+ cpldcpu_MCPU5plus_077/io_out[5] cpldcpu_MCPU5plus_077/io_out[6] cpldcpu_MCPU5plus_077/io_out[7]
+ scanchain_077/scan_select_in scanchain_078/scan_select_in vccd1 vssd1 scanchain
Xscanchain_088 scanchain_088/clk_in scanchain_089/clk_in scanchain_088/data_in scanchain_089/data_in
+ scanchain_088/latch_enable_in scanchain_089/latch_enable_in scanchain_088/module_data_in[0]
+ scanchain_088/module_data_in[1] scanchain_088/module_data_in[2] scanchain_088/module_data_in[3]
+ scanchain_088/module_data_in[4] scanchain_088/module_data_in[5] scanchain_088/module_data_in[6]
+ scanchain_088/module_data_in[7] scanchain_088/module_data_out[0] scanchain_088/module_data_out[1]
+ scanchain_088/module_data_out[2] scanchain_088/module_data_out[3] scanchain_088/module_data_out[4]
+ scanchain_088/module_data_out[5] scanchain_088/module_data_out[6] scanchain_088/module_data_out[7]
+ scanchain_088/scan_select_in scanchain_089/scan_select_in vccd1 vssd1 scanchain
Xscanchain_099 scanchain_099/clk_in scanchain_100/clk_in scanchain_099/data_in scanchain_100/data_in
+ scanchain_099/latch_enable_in scanchain_100/latch_enable_in scanchain_099/module_data_in[0]
+ scanchain_099/module_data_in[1] scanchain_099/module_data_in[2] scanchain_099/module_data_in[3]
+ scanchain_099/module_data_in[4] scanchain_099/module_data_in[5] scanchain_099/module_data_in[6]
+ scanchain_099/module_data_in[7] scanchain_099/module_data_out[0] scanchain_099/module_data_out[1]
+ scanchain_099/module_data_out[2] scanchain_099/module_data_out[3] scanchain_099/module_data_out[4]
+ scanchain_099/module_data_out[5] scanchain_099/module_data_out[6] scanchain_099/module_data_out[7]
+ scanchain_099/scan_select_in scanchain_100/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_208 scanchain_208/module_data_in[0] scanchain_208/module_data_in[1]
+ scanchain_208/module_data_in[2] scanchain_208/module_data_in[3] scanchain_208/module_data_in[4]
+ scanchain_208/module_data_in[5] scanchain_208/module_data_in[6] scanchain_208/module_data_in[7]
+ scanchain_208/module_data_out[0] scanchain_208/module_data_out[1] scanchain_208/module_data_out[2]
+ scanchain_208/module_data_out[3] scanchain_208/module_data_out[4] scanchain_208/module_data_out[5]
+ scanchain_208/module_data_out[6] scanchain_208/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_219 scanchain_219/module_data_in[0] scanchain_219/module_data_in[1]
+ scanchain_219/module_data_in[2] scanchain_219/module_data_in[3] scanchain_219/module_data_in[4]
+ scanchain_219/module_data_in[5] scanchain_219/module_data_in[6] scanchain_219/module_data_in[7]
+ scanchain_219/module_data_out[0] scanchain_219/module_data_out[1] scanchain_219/module_data_out[2]
+ scanchain_219/module_data_out[3] scanchain_219/module_data_out[4] scanchain_219/module_data_out[5]
+ scanchain_219/module_data_out[6] scanchain_219/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_347894637149553236_017 scanchain_017/module_data_in[0] scanchain_017/module_data_in[1]
+ scanchain_017/module_data_in[2] scanchain_017/module_data_in[3] scanchain_017/module_data_in[4]
+ scanchain_017/module_data_in[5] scanchain_017/module_data_in[6] scanchain_017/module_data_in[7]
+ scanchain_017/module_data_out[0] scanchain_017/module_data_out[1] scanchain_017/module_data_out[2]
+ scanchain_017/module_data_out[3] scanchain_017/module_data_out[4] scanchain_017/module_data_out[5]
+ scanchain_017/module_data_out[6] scanchain_017/module_data_out[7] vccd1 vssd1 user_module_347894637149553236
Xscanchain_237 scanchain_237/clk_in scanchain_238/clk_in scanchain_237/data_in scanchain_238/data_in
+ scanchain_237/latch_enable_in scanchain_238/latch_enable_in scanchain_237/module_data_in[0]
+ scanchain_237/module_data_in[1] scanchain_237/module_data_in[2] scanchain_237/module_data_in[3]
+ scanchain_237/module_data_in[4] scanchain_237/module_data_in[5] scanchain_237/module_data_in[6]
+ scanchain_237/module_data_in[7] scanchain_237/module_data_out[0] scanchain_237/module_data_out[1]
+ scanchain_237/module_data_out[2] scanchain_237/module_data_out[3] scanchain_237/module_data_out[4]
+ scanchain_237/module_data_out[5] scanchain_237/module_data_out[6] scanchain_237/module_data_out[7]
+ scanchain_237/scan_select_in scanchain_238/scan_select_in vccd1 vssd1 scanchain
Xscanchain_248 scanchain_248/clk_in scanchain_249/clk_in scanchain_248/data_in scanchain_249/data_in
+ scanchain_248/latch_enable_in scanchain_249/latch_enable_in scanchain_248/module_data_in[0]
+ scanchain_248/module_data_in[1] scanchain_248/module_data_in[2] scanchain_248/module_data_in[3]
+ scanchain_248/module_data_in[4] scanchain_248/module_data_in[5] scanchain_248/module_data_in[6]
+ scanchain_248/module_data_in[7] scanchain_248/module_data_out[0] scanchain_248/module_data_out[1]
+ scanchain_248/module_data_out[2] scanchain_248/module_data_out[3] scanchain_248/module_data_out[4]
+ scanchain_248/module_data_out[5] scanchain_248/module_data_out[6] scanchain_248/module_data_out[7]
+ scanchain_248/scan_select_in scanchain_249/scan_select_in vccd1 vssd1 scanchain
Xscanchain_226 scanchain_226/clk_in scanchain_227/clk_in scanchain_226/data_in scanchain_227/data_in
+ scanchain_226/latch_enable_in scanchain_227/latch_enable_in scanchain_226/module_data_in[0]
+ scanchain_226/module_data_in[1] scanchain_226/module_data_in[2] scanchain_226/module_data_in[3]
+ scanchain_226/module_data_in[4] scanchain_226/module_data_in[5] scanchain_226/module_data_in[6]
+ scanchain_226/module_data_in[7] scanchain_226/module_data_out[0] scanchain_226/module_data_out[1]
+ scanchain_226/module_data_out[2] scanchain_226/module_data_out[3] scanchain_226/module_data_out[4]
+ scanchain_226/module_data_out[5] scanchain_226/module_data_out[6] scanchain_226/module_data_out[7]
+ scanchain_226/scan_select_in scanchain_227/scan_select_in vccd1 vssd1 scanchain
Xscanchain_215 scanchain_215/clk_in scanchain_216/clk_in scanchain_215/data_in scanchain_216/data_in
+ scanchain_215/latch_enable_in scanchain_216/latch_enable_in scanchain_215/module_data_in[0]
+ scanchain_215/module_data_in[1] scanchain_215/module_data_in[2] scanchain_215/module_data_in[3]
+ scanchain_215/module_data_in[4] scanchain_215/module_data_in[5] scanchain_215/module_data_in[6]
+ scanchain_215/module_data_in[7] scanchain_215/module_data_out[0] scanchain_215/module_data_out[1]
+ scanchain_215/module_data_out[2] scanchain_215/module_data_out[3] scanchain_215/module_data_out[4]
+ scanchain_215/module_data_out[5] scanchain_215/module_data_out[6] scanchain_215/module_data_out[7]
+ scanchain_215/scan_select_in scanchain_216/scan_select_in vccd1 vssd1 scanchain
Xscanchain_204 scanchain_204/clk_in scanchain_205/clk_in scanchain_204/data_in scanchain_205/data_in
+ scanchain_204/latch_enable_in scanchain_205/latch_enable_in scanchain_204/module_data_in[0]
+ scanchain_204/module_data_in[1] scanchain_204/module_data_in[2] scanchain_204/module_data_in[3]
+ scanchain_204/module_data_in[4] scanchain_204/module_data_in[5] scanchain_204/module_data_in[6]
+ scanchain_204/module_data_in[7] scanchain_204/module_data_out[0] scanchain_204/module_data_out[1]
+ scanchain_204/module_data_out[2] scanchain_204/module_data_out[3] scanchain_204/module_data_out[4]
+ scanchain_204/module_data_out[5] scanchain_204/module_data_out[6] scanchain_204/module_data_out[7]
+ scanchain_204/scan_select_in scanchain_205/scan_select_in vccd1 vssd1 scanchain
Xalu_top_007 alu_top_007/io_in[0] alu_top_007/io_in[1] alu_top_007/io_in[2] alu_top_007/io_in[3]
+ alu_top_007/io_in[4] alu_top_007/io_in[5] alu_top_007/io_in[6] alu_top_007/io_in[7]
+ alu_top_007/io_out[0] alu_top_007/io_out[1] alu_top_007/io_out[2] alu_top_007/io_out[3]
+ alu_top_007/io_out[4] alu_top_007/io_out[5] alu_top_007/io_out[6] alu_top_007/io_out[7]
+ vccd1 vssd1 alu_top
Xscanchain_034 scanchain_034/clk_in scanchain_035/clk_in scanchain_034/data_in scanchain_035/data_in
+ scanchain_034/latch_enable_in scanchain_035/latch_enable_in scanchain_034/module_data_in[0]
+ scanchain_034/module_data_in[1] scanchain_034/module_data_in[2] scanchain_034/module_data_in[3]
+ scanchain_034/module_data_in[4] scanchain_034/module_data_in[5] scanchain_034/module_data_in[6]
+ scanchain_034/module_data_in[7] scanchain_034/module_data_out[0] scanchain_034/module_data_out[1]
+ scanchain_034/module_data_out[2] scanchain_034/module_data_out[3] scanchain_034/module_data_out[4]
+ scanchain_034/module_data_out[5] scanchain_034/module_data_out[6] scanchain_034/module_data_out[7]
+ scanchain_034/scan_select_in scanchain_035/scan_select_in vccd1 vssd1 scanchain
Xscanchain_012 scanchain_012/clk_in scanchain_013/clk_in scanchain_012/data_in scanchain_013/data_in
+ scanchain_012/latch_enable_in scanchain_013/latch_enable_in scanchain_012/module_data_in[0]
+ scanchain_012/module_data_in[1] scanchain_012/module_data_in[2] scanchain_012/module_data_in[3]
+ scanchain_012/module_data_in[4] scanchain_012/module_data_in[5] scanchain_012/module_data_in[6]
+ scanchain_012/module_data_in[7] scanchain_012/module_data_out[0] scanchain_012/module_data_out[1]
+ scanchain_012/module_data_out[2] scanchain_012/module_data_out[3] scanchain_012/module_data_out[4]
+ scanchain_012/module_data_out[5] scanchain_012/module_data_out[6] scanchain_012/module_data_out[7]
+ scanchain_012/scan_select_in scanchain_013/scan_select_in vccd1 vssd1 scanchain
Xscanchain_023 scanchain_023/clk_in scanchain_024/clk_in scanchain_023/data_in scanchain_024/data_in
+ scanchain_023/latch_enable_in scanchain_024/latch_enable_in scanchain_023/module_data_in[0]
+ scanchain_023/module_data_in[1] scanchain_023/module_data_in[2] scanchain_023/module_data_in[3]
+ scanchain_023/module_data_in[4] scanchain_023/module_data_in[5] scanchain_023/module_data_in[6]
+ scanchain_023/module_data_in[7] scanchain_023/module_data_out[0] scanchain_023/module_data_out[1]
+ scanchain_023/module_data_out[2] scanchain_023/module_data_out[3] scanchain_023/module_data_out[4]
+ scanchain_023/module_data_out[5] scanchain_023/module_data_out[6] scanchain_023/module_data_out[7]
+ scanchain_023/scan_select_in scanchain_024/scan_select_in vccd1 vssd1 scanchain
Xscanchain_001 scanchain_001/clk_in scanchain_002/clk_in scanchain_001/data_in scanchain_002/data_in
+ scanchain_001/latch_enable_in scanchain_002/latch_enable_in fraserbc_simon_001/io_in[0]
+ fraserbc_simon_001/io_in[1] fraserbc_simon_001/io_in[2] fraserbc_simon_001/io_in[3]
+ fraserbc_simon_001/io_in[4] fraserbc_simon_001/io_in[5] fraserbc_simon_001/io_in[6]
+ fraserbc_simon_001/io_in[7] fraserbc_simon_001/io_out[0] fraserbc_simon_001/io_out[1]
+ fraserbc_simon_001/io_out[2] fraserbc_simon_001/io_out[3] fraserbc_simon_001/io_out[4]
+ fraserbc_simon_001/io_out[5] fraserbc_simon_001/io_out[6] fraserbc_simon_001/io_out[7]
+ scanchain_001/scan_select_in scanchain_002/scan_select_in vccd1 vssd1 scanchain
Xscanchain_045 scanchain_045/clk_in scanchain_046/clk_in scanchain_045/data_in scanchain_046/data_in
+ scanchain_045/latch_enable_in scanchain_046/latch_enable_in scanchain_045/module_data_in[0]
+ scanchain_045/module_data_in[1] scanchain_045/module_data_in[2] scanchain_045/module_data_in[3]
+ scanchain_045/module_data_in[4] scanchain_045/module_data_in[5] scanchain_045/module_data_in[6]
+ scanchain_045/module_data_in[7] scanchain_045/module_data_out[0] scanchain_045/module_data_out[1]
+ scanchain_045/module_data_out[2] scanchain_045/module_data_out[3] scanchain_045/module_data_out[4]
+ scanchain_045/module_data_out[5] scanchain_045/module_data_out[6] scanchain_045/module_data_out[7]
+ scanchain_045/scan_select_in scanchain_046/scan_select_in vccd1 vssd1 scanchain
Xscanchain_056 scanchain_056/clk_in scanchain_057/clk_in scanchain_056/data_in scanchain_057/data_in
+ scanchain_056/latch_enable_in scanchain_057/latch_enable_in scanchain_056/module_data_in[0]
+ scanchain_056/module_data_in[1] scanchain_056/module_data_in[2] scanchain_056/module_data_in[3]
+ scanchain_056/module_data_in[4] scanchain_056/module_data_in[5] scanchain_056/module_data_in[6]
+ scanchain_056/module_data_in[7] scanchain_056/module_data_out[0] scanchain_056/module_data_out[1]
+ scanchain_056/module_data_out[2] scanchain_056/module_data_out[3] scanchain_056/module_data_out[4]
+ scanchain_056/module_data_out[5] scanchain_056/module_data_out[6] scanchain_056/module_data_out[7]
+ scanchain_056/scan_select_in scanchain_057/scan_select_in vccd1 vssd1 scanchain
Xscanchain_067 scanchain_067/clk_in scanchain_068/clk_in scanchain_067/data_in scanchain_068/data_in
+ scanchain_067/latch_enable_in scanchain_068/latch_enable_in pwm_gen_067/io_in[0]
+ pwm_gen_067/io_in[1] pwm_gen_067/io_in[2] pwm_gen_067/io_in[3] pwm_gen_067/io_in[4]
+ pwm_gen_067/io_in[5] pwm_gen_067/io_in[6] pwm_gen_067/io_in[7] pwm_gen_067/io_out[0]
+ pwm_gen_067/io_out[1] pwm_gen_067/io_out[2] pwm_gen_067/io_out[3] pwm_gen_067/io_out[4]
+ pwm_gen_067/io_out[5] pwm_gen_067/io_out[6] pwm_gen_067/io_out[7] scanchain_067/scan_select_in
+ scanchain_068/scan_select_in vccd1 vssd1 scanchain
Xmoonbase_cpu_4bit_078 moonbase_cpu_4bit_078/io_in[0] moonbase_cpu_4bit_078/io_in[1]
+ moonbase_cpu_4bit_078/io_in[2] moonbase_cpu_4bit_078/io_in[3] moonbase_cpu_4bit_078/io_in[4]
+ moonbase_cpu_4bit_078/io_in[5] moonbase_cpu_4bit_078/io_in[6] moonbase_cpu_4bit_078/io_in[7]
+ moonbase_cpu_4bit_078/io_out[0] moonbase_cpu_4bit_078/io_out[1] moonbase_cpu_4bit_078/io_out[2]
+ moonbase_cpu_4bit_078/io_out[3] moonbase_cpu_4bit_078/io_out[4] moonbase_cpu_4bit_078/io_out[5]
+ moonbase_cpu_4bit_078/io_out[6] moonbase_cpu_4bit_078/io_out[7] vccd1 vssd1 moonbase_cpu_4bit
Xscanchain_078 scanchain_078/clk_in scanchain_079/clk_in scanchain_078/data_in scanchain_079/data_in
+ scanchain_078/latch_enable_in scanchain_079/latch_enable_in moonbase_cpu_4bit_078/io_in[0]
+ moonbase_cpu_4bit_078/io_in[1] moonbase_cpu_4bit_078/io_in[2] moonbase_cpu_4bit_078/io_in[3]
+ moonbase_cpu_4bit_078/io_in[4] moonbase_cpu_4bit_078/io_in[5] moonbase_cpu_4bit_078/io_in[6]
+ moonbase_cpu_4bit_078/io_in[7] moonbase_cpu_4bit_078/io_out[0] moonbase_cpu_4bit_078/io_out[1]
+ moonbase_cpu_4bit_078/io_out[2] moonbase_cpu_4bit_078/io_out[3] moonbase_cpu_4bit_078/io_out[4]
+ moonbase_cpu_4bit_078/io_out[5] moonbase_cpu_4bit_078/io_out[6] moonbase_cpu_4bit_078/io_out[7]
+ scanchain_078/scan_select_in scanchain_079/scan_select_in vccd1 vssd1 scanchain
Xscanchain_089 scanchain_089/clk_in scanchain_090/clk_in scanchain_089/data_in scanchain_090/data_in
+ scanchain_089/latch_enable_in scanchain_090/latch_enable_in gatecat_fpga_top_089/io_in[0]
+ gatecat_fpga_top_089/io_in[1] gatecat_fpga_top_089/io_in[2] gatecat_fpga_top_089/io_in[3]
+ gatecat_fpga_top_089/io_in[4] gatecat_fpga_top_089/io_in[5] gatecat_fpga_top_089/io_in[6]
+ gatecat_fpga_top_089/io_in[7] gatecat_fpga_top_089/io_out[0] gatecat_fpga_top_089/io_out[1]
+ gatecat_fpga_top_089/io_out[2] gatecat_fpga_top_089/io_out[3] gatecat_fpga_top_089/io_out[4]
+ gatecat_fpga_top_089/io_out[5] gatecat_fpga_top_089/io_out[6] gatecat_fpga_top_089/io_out[7]
+ scanchain_089/scan_select_in scanchain_090/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341164910646919762_068 scanchain_068/module_data_in[0] scanchain_068/module_data_in[1]
+ scanchain_068/module_data_in[2] scanchain_068/module_data_in[3] scanchain_068/module_data_in[4]
+ scanchain_068/module_data_in[5] scanchain_068/module_data_in[6] scanchain_068/module_data_in[7]
+ scanchain_068/module_data_out[0] scanchain_068/module_data_out[1] scanchain_068/module_data_out[2]
+ scanchain_068/module_data_out[3] scanchain_068/module_data_out[4] scanchain_068/module_data_out[5]
+ scanchain_068/module_data_out[6] scanchain_068/module_data_out[7] vccd1 vssd1 user_module_341164910646919762
Xfraserbc_simon_001 fraserbc_simon_001/io_in[0] fraserbc_simon_001/io_in[1] fraserbc_simon_001/io_in[2]
+ fraserbc_simon_001/io_in[3] fraserbc_simon_001/io_in[4] fraserbc_simon_001/io_in[5]
+ fraserbc_simon_001/io_in[6] fraserbc_simon_001/io_in[7] fraserbc_simon_001/io_out[0]
+ fraserbc_simon_001/io_out[1] fraserbc_simon_001/io_out[2] fraserbc_simon_001/io_out[3]
+ fraserbc_simon_001/io_out[4] fraserbc_simon_001/io_out[5] fraserbc_simon_001/io_out[6]
+ fraserbc_simon_001/io_out[7] vccd1 vssd1 fraserbc_simon
Xuser_module_341535056611770964_209 scanchain_209/module_data_in[0] scanchain_209/module_data_in[1]
+ scanchain_209/module_data_in[2] scanchain_209/module_data_in[3] scanchain_209/module_data_in[4]
+ scanchain_209/module_data_in[5] scanchain_209/module_data_in[6] scanchain_209/module_data_in[7]
+ scanchain_209/module_data_out[0] scanchain_209/module_data_out[1] scanchain_209/module_data_out[2]
+ scanchain_209/module_data_out[3] scanchain_209/module_data_out[4] scanchain_209/module_data_out[5]
+ scanchain_209/module_data_out[6] scanchain_209/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xdavidsiaw_stackcalc_079 scanchain_079/module_data_in[0] scanchain_079/module_data_in[1]
+ scanchain_079/module_data_in[2] scanchain_079/module_data_in[3] scanchain_079/module_data_in[4]
+ scanchain_079/module_data_in[5] scanchain_079/module_data_in[6] scanchain_079/module_data_in[7]
+ scanchain_079/module_data_out[0] scanchain_079/module_data_out[1] scanchain_079/module_data_out[2]
+ scanchain_079/module_data_out[3] scanchain_079/module_data_out[4] scanchain_079/module_data_out[5]
+ scanchain_079/module_data_out[6] scanchain_079/module_data_out[7] vccd1 vssd1 davidsiaw_stackcalc
Xtt2_tholin_multiplier_049 scanchain_049/module_data_in[0] scanchain_049/module_data_in[1]
+ scanchain_049/module_data_in[2] scanchain_049/module_data_in[3] scanchain_049/module_data_in[4]
+ scanchain_049/module_data_in[5] scanchain_049/module_data_in[6] scanchain_049/module_data_in[7]
+ scanchain_049/module_data_out[0] scanchain_049/module_data_out[1] scanchain_049/module_data_out[2]
+ scanchain_049/module_data_out[3] scanchain_049/module_data_out[4] scanchain_049/module_data_out[5]
+ scanchain_049/module_data_out[6] scanchain_049/module_data_out[7] vccd1 vssd1 tt2_tholin_multiplier
Xuser_module_341571228858843732_082 scanchain_082/module_data_in[0] scanchain_082/module_data_in[1]
+ scanchain_082/module_data_in[2] scanchain_082/module_data_in[3] scanchain_082/module_data_in[4]
+ scanchain_082/module_data_in[5] scanchain_082/module_data_in[6] scanchain_082/module_data_in[7]
+ scanchain_082/module_data_out[0] scanchain_082/module_data_out[1] scanchain_082/module_data_out[2]
+ scanchain_082/module_data_out[3] scanchain_082/module_data_out[4] scanchain_082/module_data_out[5]
+ scanchain_082/module_data_out[6] scanchain_082/module_data_out[7] vccd1 vssd1 user_module_341571228858843732
Xscanchain_238 scanchain_238/clk_in scanchain_239/clk_in scanchain_238/data_in scanchain_239/data_in
+ scanchain_238/latch_enable_in scanchain_239/latch_enable_in scanchain_238/module_data_in[0]
+ scanchain_238/module_data_in[1] scanchain_238/module_data_in[2] scanchain_238/module_data_in[3]
+ scanchain_238/module_data_in[4] scanchain_238/module_data_in[5] scanchain_238/module_data_in[6]
+ scanchain_238/module_data_in[7] scanchain_238/module_data_out[0] scanchain_238/module_data_out[1]
+ scanchain_238/module_data_out[2] scanchain_238/module_data_out[3] scanchain_238/module_data_out[4]
+ scanchain_238/module_data_out[5] scanchain_238/module_data_out[6] scanchain_238/module_data_out[7]
+ scanchain_238/scan_select_in scanchain_239/scan_select_in vccd1 vssd1 scanchain
Xscanchain_249 scanchain_249/clk_in scanchain_249/clk_out scanchain_249/data_in scanchain_249/data_out
+ scanchain_249/latch_enable_in scanchain_249/latch_enable_out scanchain_249/module_data_in[0]
+ scanchain_249/module_data_in[1] scanchain_249/module_data_in[2] scanchain_249/module_data_in[3]
+ scanchain_249/module_data_in[4] scanchain_249/module_data_in[5] scanchain_249/module_data_in[6]
+ scanchain_249/module_data_in[7] scanchain_249/module_data_out[0] scanchain_249/module_data_out[1]
+ scanchain_249/module_data_out[2] scanchain_249/module_data_out[3] scanchain_249/module_data_out[4]
+ scanchain_249/module_data_out[5] scanchain_249/module_data_out[6] scanchain_249/module_data_out[7]
+ scanchain_249/scan_select_in scanchain_249/scan_select_out vccd1 vssd1 scanchain
Xscanchain_227 scanchain_227/clk_in scanchain_228/clk_in scanchain_227/data_in scanchain_228/data_in
+ scanchain_227/latch_enable_in scanchain_228/latch_enable_in scanchain_227/module_data_in[0]
+ scanchain_227/module_data_in[1] scanchain_227/module_data_in[2] scanchain_227/module_data_in[3]
+ scanchain_227/module_data_in[4] scanchain_227/module_data_in[5] scanchain_227/module_data_in[6]
+ scanchain_227/module_data_in[7] scanchain_227/module_data_out[0] scanchain_227/module_data_out[1]
+ scanchain_227/module_data_out[2] scanchain_227/module_data_out[3] scanchain_227/module_data_out[4]
+ scanchain_227/module_data_out[5] scanchain_227/module_data_out[6] scanchain_227/module_data_out[7]
+ scanchain_227/scan_select_in scanchain_228/scan_select_in vccd1 vssd1 scanchain
Xscanchain_216 scanchain_216/clk_in scanchain_217/clk_in scanchain_216/data_in scanchain_217/data_in
+ scanchain_216/latch_enable_in scanchain_217/latch_enable_in scanchain_216/module_data_in[0]
+ scanchain_216/module_data_in[1] scanchain_216/module_data_in[2] scanchain_216/module_data_in[3]
+ scanchain_216/module_data_in[4] scanchain_216/module_data_in[5] scanchain_216/module_data_in[6]
+ scanchain_216/module_data_in[7] scanchain_216/module_data_out[0] scanchain_216/module_data_out[1]
+ scanchain_216/module_data_out[2] scanchain_216/module_data_out[3] scanchain_216/module_data_out[4]
+ scanchain_216/module_data_out[5] scanchain_216/module_data_out[6] scanchain_216/module_data_out[7]
+ scanchain_216/scan_select_in scanchain_217/scan_select_in vccd1 vssd1 scanchain
Xscanchain_205 scanchain_205/clk_in scanchain_206/clk_in scanchain_205/data_in scanchain_206/data_in
+ scanchain_205/latch_enable_in scanchain_206/latch_enable_in scanchain_205/module_data_in[0]
+ scanchain_205/module_data_in[1] scanchain_205/module_data_in[2] scanchain_205/module_data_in[3]
+ scanchain_205/module_data_in[4] scanchain_205/module_data_in[5] scanchain_205/module_data_in[6]
+ scanchain_205/module_data_in[7] scanchain_205/module_data_out[0] scanchain_205/module_data_out[1]
+ scanchain_205/module_data_out[2] scanchain_205/module_data_out[3] scanchain_205/module_data_out[4]
+ scanchain_205/module_data_out[5] scanchain_205/module_data_out[6] scanchain_205/module_data_out[7]
+ scanchain_205/scan_select_in scanchain_206/scan_select_in vccd1 vssd1 scanchain
Xscanchain_035 scanchain_035/clk_in scanchain_036/clk_in scanchain_035/data_in scanchain_036/data_in
+ scanchain_035/latch_enable_in scanchain_036/latch_enable_in scanchain_035/module_data_in[0]
+ scanchain_035/module_data_in[1] scanchain_035/module_data_in[2] scanchain_035/module_data_in[3]
+ scanchain_035/module_data_in[4] scanchain_035/module_data_in[5] scanchain_035/module_data_in[6]
+ scanchain_035/module_data_in[7] scanchain_035/module_data_out[0] scanchain_035/module_data_out[1]
+ scanchain_035/module_data_out[2] scanchain_035/module_data_out[3] scanchain_035/module_data_out[4]
+ scanchain_035/module_data_out[5] scanchain_035/module_data_out[6] scanchain_035/module_data_out[7]
+ scanchain_035/scan_select_in scanchain_036/scan_select_in vccd1 vssd1 scanchain
Xscanchain_013 scanchain_013/clk_in scanchain_014/clk_in scanchain_013/data_in scanchain_014/data_in
+ scanchain_013/latch_enable_in scanchain_014/latch_enable_in scanchain_013/module_data_in[0]
+ scanchain_013/module_data_in[1] scanchain_013/module_data_in[2] scanchain_013/module_data_in[3]
+ scanchain_013/module_data_in[4] scanchain_013/module_data_in[5] scanchain_013/module_data_in[6]
+ scanchain_013/module_data_in[7] scanchain_013/module_data_out[0] scanchain_013/module_data_out[1]
+ scanchain_013/module_data_out[2] scanchain_013/module_data_out[3] scanchain_013/module_data_out[4]
+ scanchain_013/module_data_out[5] scanchain_013/module_data_out[6] scanchain_013/module_data_out[7]
+ scanchain_013/scan_select_in scanchain_014/scan_select_in vccd1 vssd1 scanchain
Xscanchain_024 scanchain_024/clk_in scanchain_025/clk_in scanchain_024/data_in scanchain_025/data_in
+ scanchain_024/latch_enable_in scanchain_025/latch_enable_in scanchain_024/module_data_in[0]
+ scanchain_024/module_data_in[1] scanchain_024/module_data_in[2] scanchain_024/module_data_in[3]
+ scanchain_024/module_data_in[4] scanchain_024/module_data_in[5] scanchain_024/module_data_in[6]
+ scanchain_024/module_data_in[7] scanchain_024/module_data_out[0] scanchain_024/module_data_out[1]
+ scanchain_024/module_data_out[2] scanchain_024/module_data_out[3] scanchain_024/module_data_out[4]
+ scanchain_024/module_data_out[5] scanchain_024/module_data_out[6] scanchain_024/module_data_out[7]
+ scanchain_024/scan_select_in scanchain_025/scan_select_in vccd1 vssd1 scanchain
Xscanchain_002 scanchain_002/clk_in scanchain_003/clk_in scanchain_002/data_in scanchain_003/data_in
+ scanchain_002/latch_enable_in scanchain_003/latch_enable_in tomkeddie_top_tto_002/io_in[0]
+ tomkeddie_top_tto_002/io_in[1] tomkeddie_top_tto_002/io_in[2] tomkeddie_top_tto_002/io_in[3]
+ tomkeddie_top_tto_002/io_in[4] tomkeddie_top_tto_002/io_in[5] tomkeddie_top_tto_002/io_in[6]
+ tomkeddie_top_tto_002/io_in[7] tomkeddie_top_tto_002/io_out[0] tomkeddie_top_tto_002/io_out[1]
+ tomkeddie_top_tto_002/io_out[2] tomkeddie_top_tto_002/io_out[3] tomkeddie_top_tto_002/io_out[4]
+ tomkeddie_top_tto_002/io_out[5] tomkeddie_top_tto_002/io_out[6] tomkeddie_top_tto_002/io_out[7]
+ scanchain_002/scan_select_in scanchain_003/scan_select_in vccd1 vssd1 scanchain
Xscanchain_046 scanchain_046/clk_in scanchain_047/clk_in scanchain_046/data_in scanchain_047/data_in
+ scanchain_046/latch_enable_in scanchain_047/latch_enable_in scanchain_046/module_data_in[0]
+ scanchain_046/module_data_in[1] scanchain_046/module_data_in[2] scanchain_046/module_data_in[3]
+ scanchain_046/module_data_in[4] scanchain_046/module_data_in[5] scanchain_046/module_data_in[6]
+ scanchain_046/module_data_in[7] scanchain_046/module_data_out[0] scanchain_046/module_data_out[1]
+ scanchain_046/module_data_out[2] scanchain_046/module_data_out[3] scanchain_046/module_data_out[4]
+ scanchain_046/module_data_out[5] scanchain_046/module_data_out[6] scanchain_046/module_data_out[7]
+ scanchain_046/scan_select_in scanchain_047/scan_select_in vccd1 vssd1 scanchain
Xscanchain_057 scanchain_057/clk_in scanchain_058/clk_in scanchain_057/data_in scanchain_058/data_in
+ scanchain_057/latch_enable_in scanchain_058/latch_enable_in scanchain_057/module_data_in[0]
+ scanchain_057/module_data_in[1] scanchain_057/module_data_in[2] scanchain_057/module_data_in[3]
+ scanchain_057/module_data_in[4] scanchain_057/module_data_in[5] scanchain_057/module_data_in[6]
+ scanchain_057/module_data_in[7] scanchain_057/module_data_out[0] scanchain_057/module_data_out[1]
+ scanchain_057/module_data_out[2] scanchain_057/module_data_out[3] scanchain_057/module_data_out[4]
+ scanchain_057/module_data_out[5] scanchain_057/module_data_out[6] scanchain_057/module_data_out[7]
+ scanchain_057/scan_select_in scanchain_058/scan_select_in vccd1 vssd1 scanchain
Xscanchain_079 scanchain_079/clk_in scanchain_080/clk_in scanchain_079/data_in scanchain_080/data_in
+ scanchain_079/latch_enable_in scanchain_080/latch_enable_in scanchain_079/module_data_in[0]
+ scanchain_079/module_data_in[1] scanchain_079/module_data_in[2] scanchain_079/module_data_in[3]
+ scanchain_079/module_data_in[4] scanchain_079/module_data_in[5] scanchain_079/module_data_in[6]
+ scanchain_079/module_data_in[7] scanchain_079/module_data_out[0] scanchain_079/module_data_out[1]
+ scanchain_079/module_data_out[2] scanchain_079/module_data_out[3] scanchain_079/module_data_out[4]
+ scanchain_079/module_data_out[5] scanchain_079/module_data_out[6] scanchain_079/module_data_out[7]
+ scanchain_079/scan_select_in scanchain_080/scan_select_in vccd1 vssd1 scanchain
Xscanchain_068 scanchain_068/clk_in scanchain_069/clk_in scanchain_068/data_in scanchain_069/data_in
+ scanchain_068/latch_enable_in scanchain_069/latch_enable_in scanchain_068/module_data_in[0]
+ scanchain_068/module_data_in[1] scanchain_068/module_data_in[2] scanchain_068/module_data_in[3]
+ scanchain_068/module_data_in[4] scanchain_068/module_data_in[5] scanchain_068/module_data_in[6]
+ scanchain_068/module_data_in[7] scanchain_068/module_data_out[0] scanchain_068/module_data_out[1]
+ scanchain_068/module_data_out[2] scanchain_068/module_data_out[3] scanchain_068/module_data_out[4]
+ scanchain_068/module_data_out[5] scanchain_068/module_data_out[6] scanchain_068/module_data_out[7]
+ scanchain_068/scan_select_in scanchain_069/scan_select_in vccd1 vssd1 scanchain
Xxor_shift32_evango_053 xor_shift32_evango_053/io_in[0] xor_shift32_evango_053/io_in[1]
+ xor_shift32_evango_053/io_in[2] xor_shift32_evango_053/io_in[3] xor_shift32_evango_053/io_in[4]
+ xor_shift32_evango_053/io_in[5] xor_shift32_evango_053/io_in[6] xor_shift32_evango_053/io_in[7]
+ xor_shift32_evango_053/io_out[0] xor_shift32_evango_053/io_out[1] xor_shift32_evango_053/io_out[2]
+ xor_shift32_evango_053/io_out[3] xor_shift32_evango_053/io_out[4] xor_shift32_evango_053/io_out[5]
+ xor_shift32_evango_053/io_out[6] xor_shift32_evango_053/io_out[7] vccd1 vssd1 xor_shift32_evango
Xscanchain_239 scanchain_239/clk_in scanchain_240/clk_in scanchain_239/data_in scanchain_240/data_in
+ scanchain_239/latch_enable_in scanchain_240/latch_enable_in scanchain_239/module_data_in[0]
+ scanchain_239/module_data_in[1] scanchain_239/module_data_in[2] scanchain_239/module_data_in[3]
+ scanchain_239/module_data_in[4] scanchain_239/module_data_in[5] scanchain_239/module_data_in[6]
+ scanchain_239/module_data_in[7] scanchain_239/module_data_out[0] scanchain_239/module_data_out[1]
+ scanchain_239/module_data_out[2] scanchain_239/module_data_out[3] scanchain_239/module_data_out[4]
+ scanchain_239/module_data_out[5] scanchain_239/module_data_out[6] scanchain_239/module_data_out[7]
+ scanchain_239/scan_select_in scanchain_240/scan_select_in vccd1 vssd1 scanchain
Xscanchain_228 scanchain_228/clk_in scanchain_229/clk_in scanchain_228/data_in scanchain_229/data_in
+ scanchain_228/latch_enable_in scanchain_229/latch_enable_in scanchain_228/module_data_in[0]
+ scanchain_228/module_data_in[1] scanchain_228/module_data_in[2] scanchain_228/module_data_in[3]
+ scanchain_228/module_data_in[4] scanchain_228/module_data_in[5] scanchain_228/module_data_in[6]
+ scanchain_228/module_data_in[7] scanchain_228/module_data_out[0] scanchain_228/module_data_out[1]
+ scanchain_228/module_data_out[2] scanchain_228/module_data_out[3] scanchain_228/module_data_out[4]
+ scanchain_228/module_data_out[5] scanchain_228/module_data_out[6] scanchain_228/module_data_out[7]
+ scanchain_228/scan_select_in scanchain_229/scan_select_in vccd1 vssd1 scanchain
Xscanchain_217 scanchain_217/clk_in scanchain_218/clk_in scanchain_217/data_in scanchain_218/data_in
+ scanchain_217/latch_enable_in scanchain_218/latch_enable_in scanchain_217/module_data_in[0]
+ scanchain_217/module_data_in[1] scanchain_217/module_data_in[2] scanchain_217/module_data_in[3]
+ scanchain_217/module_data_in[4] scanchain_217/module_data_in[5] scanchain_217/module_data_in[6]
+ scanchain_217/module_data_in[7] scanchain_217/module_data_out[0] scanchain_217/module_data_out[1]
+ scanchain_217/module_data_out[2] scanchain_217/module_data_out[3] scanchain_217/module_data_out[4]
+ scanchain_217/module_data_out[5] scanchain_217/module_data_out[6] scanchain_217/module_data_out[7]
+ scanchain_217/scan_select_in scanchain_218/scan_select_in vccd1 vssd1 scanchain
Xscanchain_206 scanchain_206/clk_in scanchain_207/clk_in scanchain_206/data_in scanchain_207/data_in
+ scanchain_206/latch_enable_in scanchain_207/latch_enable_in scanchain_206/module_data_in[0]
+ scanchain_206/module_data_in[1] scanchain_206/module_data_in[2] scanchain_206/module_data_in[3]
+ scanchain_206/module_data_in[4] scanchain_206/module_data_in[5] scanchain_206/module_data_in[6]
+ scanchain_206/module_data_in[7] scanchain_206/module_data_out[0] scanchain_206/module_data_out[1]
+ scanchain_206/module_data_out[2] scanchain_206/module_data_out[3] scanchain_206/module_data_out[4]
+ scanchain_206/module_data_out[5] scanchain_206/module_data_out[6] scanchain_206/module_data_out[7]
+ scanchain_206/scan_select_in scanchain_207/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_190 scanchain_190/module_data_in[0] scanchain_190/module_data_in[1]
+ scanchain_190/module_data_in[2] scanchain_190/module_data_in[3] scanchain_190/module_data_in[4]
+ scanchain_190/module_data_in[5] scanchain_190/module_data_in[6] scanchain_190/module_data_in[7]
+ scanchain_190/module_data_out[0] scanchain_190/module_data_out[1] scanchain_190/module_data_out[2]
+ scanchain_190/module_data_out[3] scanchain_190/module_data_out[4] scanchain_190/module_data_out[5]
+ scanchain_190/module_data_out[6] scanchain_190/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_047 scanchain_047/clk_in scanchain_048/clk_in scanchain_047/data_in scanchain_048/data_in
+ scanchain_047/latch_enable_in scanchain_048/latch_enable_in scanchain_047/module_data_in[0]
+ scanchain_047/module_data_in[1] scanchain_047/module_data_in[2] scanchain_047/module_data_in[3]
+ scanchain_047/module_data_in[4] scanchain_047/module_data_in[5] scanchain_047/module_data_in[6]
+ scanchain_047/module_data_in[7] scanchain_047/module_data_out[0] scanchain_047/module_data_out[1]
+ scanchain_047/module_data_out[2] scanchain_047/module_data_out[3] scanchain_047/module_data_out[4]
+ scanchain_047/module_data_out[5] scanchain_047/module_data_out[6] scanchain_047/module_data_out[7]
+ scanchain_047/scan_select_in scanchain_048/scan_select_in vccd1 vssd1 scanchain
Xscanchain_036 scanchain_036/clk_in scanchain_037/clk_in scanchain_036/data_in scanchain_037/data_in
+ scanchain_036/latch_enable_in scanchain_037/latch_enable_in jar_illegal_logic_036/io_in[0]
+ jar_illegal_logic_036/io_in[1] jar_illegal_logic_036/io_in[2] jar_illegal_logic_036/io_in[3]
+ jar_illegal_logic_036/io_in[4] jar_illegal_logic_036/io_in[5] jar_illegal_logic_036/io_in[6]
+ jar_illegal_logic_036/io_in[7] jar_illegal_logic_036/io_out[0] jar_illegal_logic_036/io_out[1]
+ jar_illegal_logic_036/io_out[2] jar_illegal_logic_036/io_out[3] jar_illegal_logic_036/io_out[4]
+ jar_illegal_logic_036/io_out[5] jar_illegal_logic_036/io_out[6] jar_illegal_logic_036/io_out[7]
+ scanchain_036/scan_select_in scanchain_037/scan_select_in vccd1 vssd1 scanchain
Xscanchain_014 scanchain_014/clk_in scanchain_015/clk_in scanchain_014/data_in scanchain_015/data_in
+ scanchain_014/latch_enable_in scanchain_015/latch_enable_in scanchain_014/module_data_in[0]
+ scanchain_014/module_data_in[1] scanchain_014/module_data_in[2] scanchain_014/module_data_in[3]
+ scanchain_014/module_data_in[4] scanchain_014/module_data_in[5] scanchain_014/module_data_in[6]
+ scanchain_014/module_data_in[7] scanchain_014/module_data_out[0] scanchain_014/module_data_out[1]
+ scanchain_014/module_data_out[2] scanchain_014/module_data_out[3] scanchain_014/module_data_out[4]
+ scanchain_014/module_data_out[5] scanchain_014/module_data_out[6] scanchain_014/module_data_out[7]
+ scanchain_014/scan_select_in scanchain_015/scan_select_in vccd1 vssd1 scanchain
Xscanchain_025 scanchain_025/clk_in scanchain_026/clk_in scanchain_025/data_in scanchain_026/data_in
+ scanchain_025/latch_enable_in scanchain_026/latch_enable_in scanchain_025/module_data_in[0]
+ scanchain_025/module_data_in[1] scanchain_025/module_data_in[2] scanchain_025/module_data_in[3]
+ scanchain_025/module_data_in[4] scanchain_025/module_data_in[5] scanchain_025/module_data_in[6]
+ scanchain_025/module_data_in[7] scanchain_025/module_data_out[0] scanchain_025/module_data_out[1]
+ scanchain_025/module_data_out[2] scanchain_025/module_data_out[3] scanchain_025/module_data_out[4]
+ scanchain_025/module_data_out[5] scanchain_025/module_data_out[6] scanchain_025/module_data_out[7]
+ scanchain_025/scan_select_in scanchain_026/scan_select_in vccd1 vssd1 scanchain
Xscanchain_003 scanchain_003/clk_in scanchain_004/clk_in scanchain_003/data_in scanchain_004/data_in
+ scanchain_003/latch_enable_in scanchain_004/latch_enable_in chrisruk_matrix_003/io_in[0]
+ chrisruk_matrix_003/io_in[1] chrisruk_matrix_003/io_in[2] chrisruk_matrix_003/io_in[3]
+ chrisruk_matrix_003/io_in[4] chrisruk_matrix_003/io_in[5] chrisruk_matrix_003/io_in[6]
+ chrisruk_matrix_003/io_in[7] chrisruk_matrix_003/io_out[0] chrisruk_matrix_003/io_out[1]
+ chrisruk_matrix_003/io_out[2] chrisruk_matrix_003/io_out[3] chrisruk_matrix_003/io_out[4]
+ chrisruk_matrix_003/io_out[5] chrisruk_matrix_003/io_out[6] chrisruk_matrix_003/io_out[7]
+ scanchain_003/scan_select_in scanchain_004/scan_select_in vccd1 vssd1 scanchain
Xscanchain_058 scanchain_058/clk_in scanchain_059/clk_in scanchain_058/data_in scanchain_059/data_in
+ scanchain_058/latch_enable_in scanchain_059/latch_enable_in user_module_nickoe_058/io_in[0]
+ user_module_nickoe_058/io_in[1] user_module_nickoe_058/io_in[2] user_module_nickoe_058/io_in[3]
+ user_module_nickoe_058/io_in[4] user_module_nickoe_058/io_in[5] user_module_nickoe_058/io_in[6]
+ user_module_nickoe_058/io_in[7] user_module_nickoe_058/io_out[0] user_module_nickoe_058/io_out[1]
+ user_module_nickoe_058/io_out[2] user_module_nickoe_058/io_out[3] user_module_nickoe_058/io_out[4]
+ user_module_nickoe_058/io_out[5] user_module_nickoe_058/io_out[6] user_module_nickoe_058/io_out[7]
+ scanchain_058/scan_select_in scanchain_059/scan_select_in vccd1 vssd1 scanchain
Xscanchain_069 scanchain_069/clk_in scanchain_070/clk_in scanchain_069/data_in scanchain_070/data_in
+ scanchain_069/latch_enable_in scanchain_070/latch_enable_in scanchain_069/module_data_in[0]
+ scanchain_069/module_data_in[1] scanchain_069/module_data_in[2] scanchain_069/module_data_in[3]
+ scanchain_069/module_data_in[4] scanchain_069/module_data_in[5] scanchain_069/module_data_in[6]
+ scanchain_069/module_data_in[7] scanchain_069/module_data_out[0] scanchain_069/module_data_out[1]
+ scanchain_069/module_data_out[2] scanchain_069/module_data_out[3] scanchain_069/module_data_out[4]
+ scanchain_069/module_data_out[5] scanchain_069/module_data_out[6] scanchain_069/module_data_out[7]
+ scanchain_069/scan_select_in scanchain_070/scan_select_in vccd1 vssd1 scanchain
Xscanchain_229 scanchain_229/clk_in scanchain_230/clk_in scanchain_229/data_in scanchain_230/data_in
+ scanchain_229/latch_enable_in scanchain_230/latch_enable_in scanchain_229/module_data_in[0]
+ scanchain_229/module_data_in[1] scanchain_229/module_data_in[2] scanchain_229/module_data_in[3]
+ scanchain_229/module_data_in[4] scanchain_229/module_data_in[5] scanchain_229/module_data_in[6]
+ scanchain_229/module_data_in[7] scanchain_229/module_data_out[0] scanchain_229/module_data_out[1]
+ scanchain_229/module_data_out[2] scanchain_229/module_data_out[3] scanchain_229/module_data_out[4]
+ scanchain_229/module_data_out[5] scanchain_229/module_data_out[6] scanchain_229/module_data_out[7]
+ scanchain_229/scan_select_in scanchain_230/scan_select_in vccd1 vssd1 scanchain
Xscanchain_218 scanchain_218/clk_in scanchain_219/clk_in scanchain_218/data_in scanchain_219/data_in
+ scanchain_218/latch_enable_in scanchain_219/latch_enable_in scanchain_218/module_data_in[0]
+ scanchain_218/module_data_in[1] scanchain_218/module_data_in[2] scanchain_218/module_data_in[3]
+ scanchain_218/module_data_in[4] scanchain_218/module_data_in[5] scanchain_218/module_data_in[6]
+ scanchain_218/module_data_in[7] scanchain_218/module_data_out[0] scanchain_218/module_data_out[1]
+ scanchain_218/module_data_out[2] scanchain_218/module_data_out[3] scanchain_218/module_data_out[4]
+ scanchain_218/module_data_out[5] scanchain_218/module_data_out[6] scanchain_218/module_data_out[7]
+ scanchain_218/scan_select_in scanchain_219/scan_select_in vccd1 vssd1 scanchain
Xscanchain_207 scanchain_207/clk_in scanchain_208/clk_in scanchain_207/data_in scanchain_208/data_in
+ scanchain_207/latch_enable_in scanchain_208/latch_enable_in scanchain_207/module_data_in[0]
+ scanchain_207/module_data_in[1] scanchain_207/module_data_in[2] scanchain_207/module_data_in[3]
+ scanchain_207/module_data_in[4] scanchain_207/module_data_in[5] scanchain_207/module_data_in[6]
+ scanchain_207/module_data_in[7] scanchain_207/module_data_out[0] scanchain_207/module_data_out[1]
+ scanchain_207/module_data_out[2] scanchain_207/module_data_out[3] scanchain_207/module_data_out[4]
+ scanchain_207/module_data_out[5] scanchain_207/module_data_out[6] scanchain_207/module_data_out[7]
+ scanchain_207/scan_select_in scanchain_208/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_180 scanchain_180/module_data_in[0] scanchain_180/module_data_in[1]
+ scanchain_180/module_data_in[2] scanchain_180/module_data_in[3] scanchain_180/module_data_in[4]
+ scanchain_180/module_data_in[5] scanchain_180/module_data_in[6] scanchain_180/module_data_in[7]
+ scanchain_180/module_data_out[0] scanchain_180/module_data_out[1] scanchain_180/module_data_out[2]
+ scanchain_180/module_data_out[3] scanchain_180/module_data_out[4] scanchain_180/module_data_out[5]
+ scanchain_180/module_data_out[6] scanchain_180/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_191 scanchain_191/module_data_in[0] scanchain_191/module_data_in[1]
+ scanchain_191/module_data_in[2] scanchain_191/module_data_in[3] scanchain_191/module_data_in[4]
+ scanchain_191/module_data_in[5] scanchain_191/module_data_in[6] scanchain_191/module_data_in[7]
+ scanchain_191/module_data_out[0] scanchain_191/module_data_out[1] scanchain_191/module_data_out[2]
+ scanchain_191/module_data_out[3] scanchain_191/module_data_out[4] scanchain_191/module_data_out[5]
+ scanchain_191/module_data_out[6] scanchain_191/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_048 scanchain_048/clk_in scanchain_049/clk_in scanchain_048/data_in scanchain_049/data_in
+ scanchain_048/latch_enable_in scanchain_049/latch_enable_in scanchain_048/module_data_in[0]
+ scanchain_048/module_data_in[1] scanchain_048/module_data_in[2] scanchain_048/module_data_in[3]
+ scanchain_048/module_data_in[4] scanchain_048/module_data_in[5] scanchain_048/module_data_in[6]
+ scanchain_048/module_data_in[7] scanchain_048/module_data_out[0] scanchain_048/module_data_out[1]
+ scanchain_048/module_data_out[2] scanchain_048/module_data_out[3] scanchain_048/module_data_out[4]
+ scanchain_048/module_data_out[5] scanchain_048/module_data_out[6] scanchain_048/module_data_out[7]
+ scanchain_048/scan_select_in scanchain_049/scan_select_in vccd1 vssd1 scanchain
Xgithub_com_proppy_tt02_xls_counter_051 scanchain_051/module_data_in[0] scanchain_051/module_data_in[1]
+ scanchain_051/module_data_in[2] scanchain_051/module_data_in[3] scanchain_051/module_data_in[4]
+ scanchain_051/module_data_in[5] scanchain_051/module_data_in[6] scanchain_051/module_data_in[7]
+ scanchain_051/module_data_out[0] scanchain_051/module_data_out[1] scanchain_051/module_data_out[2]
+ scanchain_051/module_data_out[3] scanchain_051/module_data_out[4] scanchain_051/module_data_out[5]
+ scanchain_051/module_data_out[6] scanchain_051/module_data_out[7] vccd1 vssd1 github_com_proppy_tt02_xls_counter
Xscanchain_037 scanchain_037/clk_in scanchain_038/clk_in scanchain_037/data_in scanchain_038/data_in
+ scanchain_037/latch_enable_in scanchain_038/latch_enable_in scanchain_037/module_data_in[0]
+ scanchain_037/module_data_in[1] scanchain_037/module_data_in[2] scanchain_037/module_data_in[3]
+ scanchain_037/module_data_in[4] scanchain_037/module_data_in[5] scanchain_037/module_data_in[6]
+ scanchain_037/module_data_in[7] scanchain_037/module_data_out[0] scanchain_037/module_data_out[1]
+ scanchain_037/module_data_out[2] scanchain_037/module_data_out[3] scanchain_037/module_data_out[4]
+ scanchain_037/module_data_out[5] scanchain_037/module_data_out[6] scanchain_037/module_data_out[7]
+ scanchain_037/scan_select_in scanchain_038/scan_select_in vccd1 vssd1 scanchain
Xscanchain_026 scanchain_026/clk_in scanchain_027/clk_in scanchain_026/data_in scanchain_027/data_in
+ scanchain_026/latch_enable_in scanchain_027/latch_enable_in mm21_LEDMatrixTop_026/io_in[0]
+ mm21_LEDMatrixTop_026/io_in[1] mm21_LEDMatrixTop_026/io_in[2] mm21_LEDMatrixTop_026/io_in[3]
+ mm21_LEDMatrixTop_026/io_in[4] mm21_LEDMatrixTop_026/io_in[5] mm21_LEDMatrixTop_026/io_in[6]
+ mm21_LEDMatrixTop_026/io_in[7] mm21_LEDMatrixTop_026/io_out[0] mm21_LEDMatrixTop_026/io_out[1]
+ mm21_LEDMatrixTop_026/io_out[2] mm21_LEDMatrixTop_026/io_out[3] mm21_LEDMatrixTop_026/io_out[4]
+ mm21_LEDMatrixTop_026/io_out[5] mm21_LEDMatrixTop_026/io_out[6] mm21_LEDMatrixTop_026/io_out[7]
+ scanchain_026/scan_select_in scanchain_027/scan_select_in vccd1 vssd1 scanchain
Xscanchain_015 scanchain_015/clk_in scanchain_016/clk_in scanchain_015/data_in scanchain_016/data_in
+ scanchain_015/latch_enable_in scanchain_016/latch_enable_in tiny_fft_015/io_in[0]
+ tiny_fft_015/io_in[1] tiny_fft_015/io_in[2] tiny_fft_015/io_in[3] tiny_fft_015/io_in[4]
+ tiny_fft_015/io_in[5] tiny_fft_015/io_in[6] tiny_fft_015/io_in[7] tiny_fft_015/io_out[0]
+ tiny_fft_015/io_out[1] tiny_fft_015/io_out[2] tiny_fft_015/io_out[3] tiny_fft_015/io_out[4]
+ tiny_fft_015/io_out[5] tiny_fft_015/io_out[6] tiny_fft_015/io_out[7] scanchain_015/scan_select_in
+ scanchain_016/scan_select_in vccd1 vssd1 scanchain
Xscanchain_004 scanchain_004/clk_in scanchain_005/clk_in scanchain_004/data_in scanchain_005/data_in
+ scanchain_004/latch_enable_in scanchain_005/latch_enable_in loxodes_sequencer_004/io_in[0]
+ loxodes_sequencer_004/io_in[1] loxodes_sequencer_004/io_in[2] loxodes_sequencer_004/io_in[3]
+ loxodes_sequencer_004/io_in[4] loxodes_sequencer_004/io_in[5] loxodes_sequencer_004/io_in[6]
+ loxodes_sequencer_004/io_in[7] loxodes_sequencer_004/io_out[0] loxodes_sequencer_004/io_out[1]
+ loxodes_sequencer_004/io_out[2] loxodes_sequencer_004/io_out[3] loxodes_sequencer_004/io_out[4]
+ loxodes_sequencer_004/io_out[5] loxodes_sequencer_004/io_out[6] loxodes_sequencer_004/io_out[7]
+ scanchain_004/scan_select_in scanchain_005/scan_select_in vccd1 vssd1 scanchain
Xscanchain_059 scanchain_059/clk_in scanchain_060/clk_in scanchain_059/data_in scanchain_060/data_in
+ scanchain_059/latch_enable_in scanchain_060/latch_enable_in scanchain_059/module_data_in[0]
+ scanchain_059/module_data_in[1] scanchain_059/module_data_in[2] scanchain_059/module_data_in[3]
+ scanchain_059/module_data_in[4] scanchain_059/module_data_in[5] scanchain_059/module_data_in[6]
+ scanchain_059/module_data_in[7] scanchain_059/module_data_out[0] scanchain_059/module_data_out[1]
+ scanchain_059/module_data_out[2] scanchain_059/module_data_out[3] scanchain_059/module_data_out[4]
+ scanchain_059/module_data_out[5] scanchain_059/module_data_out[6] scanchain_059/module_data_out[7]
+ scanchain_059/scan_select_in scanchain_060/scan_select_in vccd1 vssd1 scanchain
Xtt2_tholin_multiplexed_counter_050 scanchain_050/module_data_in[0] scanchain_050/module_data_in[1]
+ scanchain_050/module_data_in[2] scanchain_050/module_data_in[3] scanchain_050/module_data_in[4]
+ scanchain_050/module_data_in[5] scanchain_050/module_data_in[6] scanchain_050/module_data_in[7]
+ scanchain_050/module_data_out[0] scanchain_050/module_data_out[1] scanchain_050/module_data_out[2]
+ scanchain_050/module_data_out[3] scanchain_050/module_data_out[4] scanchain_050/module_data_out[5]
+ scanchain_050/module_data_out[6] scanchain_050/module_data_out[7] vccd1 vssd1 tt2_tholin_multiplexed_counter
Xasic_multiplier_wrapper_023 scanchain_023/module_data_in[0] scanchain_023/module_data_in[1]
+ scanchain_023/module_data_in[2] scanchain_023/module_data_in[3] scanchain_023/module_data_in[4]
+ scanchain_023/module_data_in[5] scanchain_023/module_data_in[6] scanchain_023/module_data_in[7]
+ scanchain_023/module_data_out[0] scanchain_023/module_data_out[1] scanchain_023/module_data_out[2]
+ scanchain_023/module_data_out[3] scanchain_023/module_data_out[4] scanchain_023/module_data_out[5]
+ scanchain_023/module_data_out[6] scanchain_023/module_data_out[7] vccd1 vssd1 asic_multiplier_wrapper
Xuser_module_349405063877231188_061 scanchain_061/module_data_in[0] scanchain_061/module_data_in[1]
+ scanchain_061/module_data_in[2] scanchain_061/module_data_in[3] scanchain_061/module_data_in[4]
+ scanchain_061/module_data_in[5] scanchain_061/module_data_in[6] scanchain_061/module_data_in[7]
+ scanchain_061/module_data_out[0] scanchain_061/module_data_out[1] scanchain_061/module_data_out[2]
+ scanchain_061/module_data_out[3] scanchain_061/module_data_out[4] scanchain_061/module_data_out[5]
+ scanchain_061/module_data_out[6] scanchain_061/module_data_out[7] vccd1 vssd1 user_module_349405063877231188
Xpwm_gen_067 pwm_gen_067/io_in[0] pwm_gen_067/io_in[1] pwm_gen_067/io_in[2] pwm_gen_067/io_in[3]
+ pwm_gen_067/io_in[4] pwm_gen_067/io_in[5] pwm_gen_067/io_in[6] pwm_gen_067/io_in[7]
+ pwm_gen_067/io_out[0] pwm_gen_067/io_out[1] pwm_gen_067/io_out[2] pwm_gen_067/io_out[3]
+ pwm_gen_067/io_out[4] pwm_gen_067/io_out[5] pwm_gen_067/io_out[6] pwm_gen_067/io_out[7]
+ vccd1 vssd1 pwm_gen
Xscanchain_208 scanchain_208/clk_in scanchain_209/clk_in scanchain_208/data_in scanchain_209/data_in
+ scanchain_208/latch_enable_in scanchain_209/latch_enable_in scanchain_208/module_data_in[0]
+ scanchain_208/module_data_in[1] scanchain_208/module_data_in[2] scanchain_208/module_data_in[3]
+ scanchain_208/module_data_in[4] scanchain_208/module_data_in[5] scanchain_208/module_data_in[6]
+ scanchain_208/module_data_in[7] scanchain_208/module_data_out[0] scanchain_208/module_data_out[1]
+ scanchain_208/module_data_out[2] scanchain_208/module_data_out[3] scanchain_208/module_data_out[4]
+ scanchain_208/module_data_out[5] scanchain_208/module_data_out[6] scanchain_208/module_data_out[7]
+ scanchain_208/scan_select_in scanchain_209/scan_select_in vccd1 vssd1 scanchain
Xscanchain_219 scanchain_219/clk_in scanchain_220/clk_in scanchain_219/data_in scanchain_220/data_in
+ scanchain_219/latch_enable_in scanchain_220/latch_enable_in scanchain_219/module_data_in[0]
+ scanchain_219/module_data_in[1] scanchain_219/module_data_in[2] scanchain_219/module_data_in[3]
+ scanchain_219/module_data_in[4] scanchain_219/module_data_in[5] scanchain_219/module_data_in[6]
+ scanchain_219/module_data_in[7] scanchain_219/module_data_out[0] scanchain_219/module_data_out[1]
+ scanchain_219/module_data_out[2] scanchain_219/module_data_out[3] scanchain_219/module_data_out[4]
+ scanchain_219/module_data_out[5] scanchain_219/module_data_out[6] scanchain_219/module_data_out[7]
+ scanchain_219/scan_select_in scanchain_220/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_181 scanchain_181/module_data_in[0] scanchain_181/module_data_in[1]
+ scanchain_181/module_data_in[2] scanchain_181/module_data_in[3] scanchain_181/module_data_in[4]
+ scanchain_181/module_data_in[5] scanchain_181/module_data_in[6] scanchain_181/module_data_in[7]
+ scanchain_181/module_data_out[0] scanchain_181/module_data_out[1] scanchain_181/module_data_out[2]
+ scanchain_181/module_data_out[3] scanchain_181/module_data_out[4] scanchain_181/module_data_out[5]
+ scanchain_181/module_data_out[6] scanchain_181/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_049 scanchain_049/clk_in scanchain_050/clk_in scanchain_049/data_in scanchain_050/data_in
+ scanchain_049/latch_enable_in scanchain_050/latch_enable_in scanchain_049/module_data_in[0]
+ scanchain_049/module_data_in[1] scanchain_049/module_data_in[2] scanchain_049/module_data_in[3]
+ scanchain_049/module_data_in[4] scanchain_049/module_data_in[5] scanchain_049/module_data_in[6]
+ scanchain_049/module_data_in[7] scanchain_049/module_data_out[0] scanchain_049/module_data_out[1]
+ scanchain_049/module_data_out[2] scanchain_049/module_data_out[3] scanchain_049/module_data_out[4]
+ scanchain_049/module_data_out[5] scanchain_049/module_data_out[6] scanchain_049/module_data_out[7]
+ scanchain_049/scan_select_in scanchain_050/scan_select_in vccd1 vssd1 scanchain
Xscanchain_038 scanchain_038/clk_in scanchain_039/clk_in scanchain_038/data_in scanchain_039/data_in
+ scanchain_038/latch_enable_in scanchain_039/latch_enable_in thezoq2_yafpga_038/io_in[0]
+ thezoq2_yafpga_038/io_in[1] thezoq2_yafpga_038/io_in[2] thezoq2_yafpga_038/io_in[3]
+ thezoq2_yafpga_038/io_in[4] thezoq2_yafpga_038/io_in[5] thezoq2_yafpga_038/io_in[6]
+ thezoq2_yafpga_038/io_in[7] thezoq2_yafpga_038/io_out[0] thezoq2_yafpga_038/io_out[1]
+ thezoq2_yafpga_038/io_out[2] thezoq2_yafpga_038/io_out[3] thezoq2_yafpga_038/io_out[4]
+ thezoq2_yafpga_038/io_out[5] thezoq2_yafpga_038/io_out[6] thezoq2_yafpga_038/io_out[7]
+ scanchain_038/scan_select_in scanchain_039/scan_select_in vccd1 vssd1 scanchain
Xscanchain_027 scanchain_027/clk_in scanchain_028/clk_in scanchain_027/data_in scanchain_028/data_in
+ scanchain_027/latch_enable_in scanchain_028/latch_enable_in scanchain_027/module_data_in[0]
+ scanchain_027/module_data_in[1] scanchain_027/module_data_in[2] scanchain_027/module_data_in[3]
+ scanchain_027/module_data_in[4] scanchain_027/module_data_in[5] scanchain_027/module_data_in[6]
+ scanchain_027/module_data_in[7] scanchain_027/module_data_out[0] scanchain_027/module_data_out[1]
+ scanchain_027/module_data_out[2] scanchain_027/module_data_out[3] scanchain_027/module_data_out[4]
+ scanchain_027/module_data_out[5] scanchain_027/module_data_out[6] scanchain_027/module_data_out[7]
+ scanchain_027/scan_select_in scanchain_028/scan_select_in vccd1 vssd1 scanchain
Xscanchain_016 scanchain_016/clk_in scanchain_017/clk_in scanchain_016/data_in scanchain_017/data_in
+ scanchain_016/latch_enable_in scanchain_017/latch_enable_in scanchain_016/module_data_in[0]
+ scanchain_016/module_data_in[1] scanchain_016/module_data_in[2] scanchain_016/module_data_in[3]
+ scanchain_016/module_data_in[4] scanchain_016/module_data_in[5] scanchain_016/module_data_in[6]
+ scanchain_016/module_data_in[7] scanchain_016/module_data_out[0] scanchain_016/module_data_out[1]
+ scanchain_016/module_data_out[2] scanchain_016/module_data_out[3] scanchain_016/module_data_out[4]
+ scanchain_016/module_data_out[5] scanchain_016/module_data_out[6] scanchain_016/module_data_out[7]
+ scanchain_016/scan_select_in scanchain_017/scan_select_in vccd1 vssd1 scanchain
Xscanchain_005 scanchain_005/clk_in scanchain_006/clk_in scanchain_005/data_in scanchain_006/data_in
+ scanchain_005/latch_enable_in scanchain_006/latch_enable_in migcorre_pwm_005/io_in[0]
+ migcorre_pwm_005/io_in[1] migcorre_pwm_005/io_in[2] migcorre_pwm_005/io_in[3] migcorre_pwm_005/io_in[4]
+ migcorre_pwm_005/io_in[5] migcorre_pwm_005/io_in[6] migcorre_pwm_005/io_in[7] migcorre_pwm_005/io_out[0]
+ migcorre_pwm_005/io_out[1] migcorre_pwm_005/io_out[2] migcorre_pwm_005/io_out[3]
+ migcorre_pwm_005/io_out[4] migcorre_pwm_005/io_out[5] migcorre_pwm_005/io_out[6]
+ migcorre_pwm_005/io_out[7] scanchain_005/scan_select_in scanchain_006/scan_select_in
+ vccd1 vssd1 scanchain
Xuser_module_341535056611770964_170 scanchain_170/module_data_in[0] scanchain_170/module_data_in[1]
+ scanchain_170/module_data_in[2] scanchain_170/module_data_in[3] scanchain_170/module_data_in[4]
+ scanchain_170/module_data_in[5] scanchain_170/module_data_in[6] scanchain_170/module_data_in[7]
+ scanchain_170/module_data_out[0] scanchain_170/module_data_out[1] scanchain_170/module_data_out[2]
+ scanchain_170/module_data_out[3] scanchain_170/module_data_out[4] scanchain_170/module_data_out[5]
+ scanchain_170/module_data_out[6] scanchain_170/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_192 scanchain_192/module_data_in[0] scanchain_192/module_data_in[1]
+ scanchain_192/module_data_in[2] scanchain_192/module_data_in[3] scanchain_192/module_data_in[4]
+ scanchain_192/module_data_in[5] scanchain_192/module_data_in[6] scanchain_192/module_data_in[7]
+ scanchain_192/module_data_out[0] scanchain_192/module_data_out[1] scanchain_192/module_data_out[2]
+ scanchain_192/module_data_out[3] scanchain_192/module_data_out[4] scanchain_192/module_data_out[5]
+ scanchain_192/module_data_out[6] scanchain_192/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_209 scanchain_209/clk_in scanchain_210/clk_in scanchain_209/data_in scanchain_210/data_in
+ scanchain_209/latch_enable_in scanchain_210/latch_enable_in scanchain_209/module_data_in[0]
+ scanchain_209/module_data_in[1] scanchain_209/module_data_in[2] scanchain_209/module_data_in[3]
+ scanchain_209/module_data_in[4] scanchain_209/module_data_in[5] scanchain_209/module_data_in[6]
+ scanchain_209/module_data_in[7] scanchain_209/module_data_out[0] scanchain_209/module_data_out[1]
+ scanchain_209/module_data_out[2] scanchain_209/module_data_out[3] scanchain_209/module_data_out[4]
+ scanchain_209/module_data_out[5] scanchain_209/module_data_out[6] scanchain_209/module_data_out[7]
+ scanchain_209/scan_select_in scanchain_210/scan_select_in vccd1 vssd1 scanchain
Xscanchain_039 scanchain_039/clk_in scanchain_040/clk_in scanchain_039/data_in scanchain_040/data_in
+ scanchain_039/latch_enable_in scanchain_040/latch_enable_in moyes0_top_module_039/io_in[0]
+ moyes0_top_module_039/io_in[1] moyes0_top_module_039/io_in[2] moyes0_top_module_039/io_in[3]
+ moyes0_top_module_039/io_in[4] moyes0_top_module_039/io_in[5] moyes0_top_module_039/io_in[6]
+ moyes0_top_module_039/io_in[7] moyes0_top_module_039/io_out[0] moyes0_top_module_039/io_out[1]
+ moyes0_top_module_039/io_out[2] moyes0_top_module_039/io_out[3] moyes0_top_module_039/io_out[4]
+ moyes0_top_module_039/io_out[5] moyes0_top_module_039/io_out[6] moyes0_top_module_039/io_out[7]
+ scanchain_039/scan_select_in scanchain_040/scan_select_in vccd1 vssd1 scanchain
Xscanchain_028 scanchain_028/clk_in scanchain_029/clk_in scanchain_028/data_in scanchain_029/data_in
+ scanchain_028/latch_enable_in scanchain_029/latch_enable_in scanchain_028/module_data_in[0]
+ scanchain_028/module_data_in[1] scanchain_028/module_data_in[2] scanchain_028/module_data_in[3]
+ scanchain_028/module_data_in[4] scanchain_028/module_data_in[5] scanchain_028/module_data_in[6]
+ scanchain_028/module_data_in[7] scanchain_028/module_data_out[0] scanchain_028/module_data_out[1]
+ scanchain_028/module_data_out[2] scanchain_028/module_data_out[3] scanchain_028/module_data_out[4]
+ scanchain_028/module_data_out[5] scanchain_028/module_data_out[6] scanchain_028/module_data_out[7]
+ scanchain_028/scan_select_in scanchain_029/scan_select_in vccd1 vssd1 scanchain
Xscanchain_017 scanchain_017/clk_in scanchain_018/clk_in scanchain_017/data_in scanchain_018/data_in
+ scanchain_017/latch_enable_in scanchain_018/latch_enable_in scanchain_017/module_data_in[0]
+ scanchain_017/module_data_in[1] scanchain_017/module_data_in[2] scanchain_017/module_data_in[3]
+ scanchain_017/module_data_in[4] scanchain_017/module_data_in[5] scanchain_017/module_data_in[6]
+ scanchain_017/module_data_in[7] scanchain_017/module_data_out[0] scanchain_017/module_data_out[1]
+ scanchain_017/module_data_out[2] scanchain_017/module_data_out[3] scanchain_017/module_data_out[4]
+ scanchain_017/module_data_out[5] scanchain_017/module_data_out[6] scanchain_017/module_data_out[7]
+ scanchain_017/scan_select_in scanchain_018/scan_select_in vccd1 vssd1 scanchain
Xscanchain_006 scanchain_006/clk_in scanchain_007/clk_in scanchain_006/data_in scanchain_007/data_in
+ scanchain_006/latch_enable_in scanchain_007/latch_enable_in s4ga_006/io_in[0] s4ga_006/io_in[1]
+ s4ga_006/io_in[2] s4ga_006/io_in[3] s4ga_006/io_in[4] s4ga_006/io_in[5] s4ga_006/io_in[6]
+ s4ga_006/io_in[7] s4ga_006/io_out[0] s4ga_006/io_out[1] s4ga_006/io_out[2] s4ga_006/io_out[3]
+ s4ga_006/io_out[4] s4ga_006/io_out[5] s4ga_006/io_out[6] s4ga_006/io_out[7] scanchain_006/scan_select_in
+ scanchain_007/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_160 scanchain_160/module_data_in[0] scanchain_160/module_data_in[1]
+ scanchain_160/module_data_in[2] scanchain_160/module_data_in[3] scanchain_160/module_data_in[4]
+ scanchain_160/module_data_in[5] scanchain_160/module_data_in[6] scanchain_160/module_data_in[7]
+ scanchain_160/module_data_out[0] scanchain_160/module_data_out[1] scanchain_160/module_data_out[2]
+ scanchain_160/module_data_out[3] scanchain_160/module_data_out[4] scanchain_160/module_data_out[5]
+ scanchain_160/module_data_out[6] scanchain_160/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_171 scanchain_171/module_data_in[0] scanchain_171/module_data_in[1]
+ scanchain_171/module_data_in[2] scanchain_171/module_data_in[3] scanchain_171/module_data_in[4]
+ scanchain_171/module_data_in[5] scanchain_171/module_data_in[6] scanchain_171/module_data_in[7]
+ scanchain_171/module_data_out[0] scanchain_171/module_data_out[1] scanchain_171/module_data_out[2]
+ scanchain_171/module_data_out[3] scanchain_171/module_data_out[4] scanchain_171/module_data_out[5]
+ scanchain_171/module_data_out[6] scanchain_171/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_193 scanchain_193/module_data_in[0] scanchain_193/module_data_in[1]
+ scanchain_193/module_data_in[2] scanchain_193/module_data_in[3] scanchain_193/module_data_in[4]
+ scanchain_193/module_data_in[5] scanchain_193/module_data_in[6] scanchain_193/module_data_in[7]
+ scanchain_193/module_data_out[0] scanchain_193/module_data_out[1] scanchain_193/module_data_out[2]
+ scanchain_193/module_data_out[3] scanchain_193/module_data_out[4] scanchain_193/module_data_out[5]
+ scanchain_193/module_data_out[6] scanchain_193/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_182 scanchain_182/module_data_in[0] scanchain_182/module_data_in[1]
+ scanchain_182/module_data_in[2] scanchain_182/module_data_in[3] scanchain_182/module_data_in[4]
+ scanchain_182/module_data_in[5] scanchain_182/module_data_in[6] scanchain_182/module_data_in[7]
+ scanchain_182/module_data_out[0] scanchain_182/module_data_out[1] scanchain_182/module_data_out[2]
+ scanchain_182/module_data_out[3] scanchain_182/module_data_out[4] scanchain_182/module_data_out[5]
+ scanchain_182/module_data_out[6] scanchain_182/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_348195845106041428_027 scanchain_027/module_data_in[0] scanchain_027/module_data_in[1]
+ scanchain_027/module_data_in[2] scanchain_027/module_data_in[3] scanchain_027/module_data_in[4]
+ scanchain_027/module_data_in[5] scanchain_027/module_data_in[6] scanchain_027/module_data_in[7]
+ scanchain_027/module_data_out[0] scanchain_027/module_data_out[1] scanchain_027/module_data_out[2]
+ scanchain_027/module_data_out[3] scanchain_027/module_data_out[4] scanchain_027/module_data_out[5]
+ scanchain_027/module_data_out[6] scanchain_027/module_data_out[7] vccd1 vssd1 user_module_348195845106041428
Xaidan_McCoy_008 aidan_McCoy_008/io_in[0] aidan_McCoy_008/io_in[1] aidan_McCoy_008/io_in[2]
+ aidan_McCoy_008/io_in[3] aidan_McCoy_008/io_in[4] aidan_McCoy_008/io_in[5] aidan_McCoy_008/io_in[6]
+ aidan_McCoy_008/io_in[7] aidan_McCoy_008/io_out[0] aidan_McCoy_008/io_out[1] aidan_McCoy_008/io_out[2]
+ aidan_McCoy_008/io_out[3] aidan_McCoy_008/io_out[4] aidan_McCoy_008/io_out[5] aidan_McCoy_008/io_out[6]
+ aidan_McCoy_008/io_out[7] vccd1 vssd1 aidan_McCoy
Xuser_module_341609034095264340_069 scanchain_069/module_data_in[0] scanchain_069/module_data_in[1]
+ scanchain_069/module_data_in[2] scanchain_069/module_data_in[3] scanchain_069/module_data_in[4]
+ scanchain_069/module_data_in[5] scanchain_069/module_data_in[6] scanchain_069/module_data_in[7]
+ scanchain_069/module_data_out[0] scanchain_069/module_data_out[1] scanchain_069/module_data_out[2]
+ scanchain_069/module_data_out[3] scanchain_069/module_data_out[4] scanchain_069/module_data_out[5]
+ scanchain_069/module_data_out[6] scanchain_069/module_data_out[7] vccd1 vssd1 user_module_341609034095264340
Xuser_module_341535056611770964_194 scanchain_194/module_data_in[0] scanchain_194/module_data_in[1]
+ scanchain_194/module_data_in[2] scanchain_194/module_data_in[3] scanchain_194/module_data_in[4]
+ scanchain_194/module_data_in[5] scanchain_194/module_data_in[6] scanchain_194/module_data_in[7]
+ scanchain_194/module_data_out[0] scanchain_194/module_data_out[1] scanchain_194/module_data_out[2]
+ scanchain_194/module_data_out[3] scanchain_194/module_data_out[4] scanchain_194/module_data_out[5]
+ scanchain_194/module_data_out[6] scanchain_194/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_029 scanchain_029/clk_in scanchain_030/clk_in scanchain_029/data_in scanchain_030/data_in
+ scanchain_029/latch_enable_in scanchain_030/latch_enable_in yubex_egg_timer_029/io_in[0]
+ yubex_egg_timer_029/io_in[1] yubex_egg_timer_029/io_in[2] yubex_egg_timer_029/io_in[3]
+ yubex_egg_timer_029/io_in[4] yubex_egg_timer_029/io_in[5] yubex_egg_timer_029/io_in[6]
+ yubex_egg_timer_029/io_in[7] yubex_egg_timer_029/io_out[0] yubex_egg_timer_029/io_out[1]
+ yubex_egg_timer_029/io_out[2] yubex_egg_timer_029/io_out[3] yubex_egg_timer_029/io_out[4]
+ yubex_egg_timer_029/io_out[5] yubex_egg_timer_029/io_out[6] yubex_egg_timer_029/io_out[7]
+ scanchain_029/scan_select_in scanchain_030/scan_select_in vccd1 vssd1 scanchain
Xscanchain_018 scanchain_018/clk_in scanchain_019/clk_in scanchain_018/data_in scanchain_019/data_in
+ scanchain_018/latch_enable_in scanchain_019/latch_enable_in scanchain_018/module_data_in[0]
+ scanchain_018/module_data_in[1] scanchain_018/module_data_in[2] scanchain_018/module_data_in[3]
+ scanchain_018/module_data_in[4] scanchain_018/module_data_in[5] scanchain_018/module_data_in[6]
+ scanchain_018/module_data_in[7] scanchain_018/module_data_out[0] scanchain_018/module_data_out[1]
+ scanchain_018/module_data_out[2] scanchain_018/module_data_out[3] scanchain_018/module_data_out[4]
+ scanchain_018/module_data_out[5] scanchain_018/module_data_out[6] scanchain_018/module_data_out[7]
+ scanchain_018/scan_select_in scanchain_019/scan_select_in vccd1 vssd1 scanchain
Xscanchain_007 scanchain_007/clk_in scanchain_008/clk_in scanchain_007/data_in scanchain_008/data_in
+ scanchain_007/latch_enable_in scanchain_008/latch_enable_in alu_top_007/io_in[0]
+ alu_top_007/io_in[1] alu_top_007/io_in[2] alu_top_007/io_in[3] alu_top_007/io_in[4]
+ alu_top_007/io_in[5] alu_top_007/io_in[6] alu_top_007/io_in[7] alu_top_007/io_out[0]
+ alu_top_007/io_out[1] alu_top_007/io_out[2] alu_top_007/io_out[3] alu_top_007/io_out[4]
+ alu_top_007/io_out[5] alu_top_007/io_out[6] alu_top_007/io_out[7] scanchain_007/scan_select_in
+ scanchain_008/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_150 scanchain_150/module_data_in[0] scanchain_150/module_data_in[1]
+ scanchain_150/module_data_in[2] scanchain_150/module_data_in[3] scanchain_150/module_data_in[4]
+ scanchain_150/module_data_in[5] scanchain_150/module_data_in[6] scanchain_150/module_data_in[7]
+ scanchain_150/module_data_out[0] scanchain_150/module_data_out[1] scanchain_150/module_data_out[2]
+ scanchain_150/module_data_out[3] scanchain_150/module_data_out[4] scanchain_150/module_data_out[5]
+ scanchain_150/module_data_out[6] scanchain_150/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_161 scanchain_161/module_data_in[0] scanchain_161/module_data_in[1]
+ scanchain_161/module_data_in[2] scanchain_161/module_data_in[3] scanchain_161/module_data_in[4]
+ scanchain_161/module_data_in[5] scanchain_161/module_data_in[6] scanchain_161/module_data_in[7]
+ scanchain_161/module_data_out[0] scanchain_161/module_data_out[1] scanchain_161/module_data_out[2]
+ scanchain_161/module_data_out[3] scanchain_161/module_data_out[4] scanchain_161/module_data_out[5]
+ scanchain_161/module_data_out[6] scanchain_161/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_172 scanchain_172/module_data_in[0] scanchain_172/module_data_in[1]
+ scanchain_172/module_data_in[2] scanchain_172/module_data_in[3] scanchain_172/module_data_in[4]
+ scanchain_172/module_data_in[5] scanchain_172/module_data_in[6] scanchain_172/module_data_in[7]
+ scanchain_172/module_data_out[0] scanchain_172/module_data_out[1] scanchain_172/module_data_out[2]
+ scanchain_172/module_data_out[3] scanchain_172/module_data_out[4] scanchain_172/module_data_out[5]
+ scanchain_172/module_data_out[6] scanchain_172/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_183 scanchain_183/module_data_in[0] scanchain_183/module_data_in[1]
+ scanchain_183/module_data_in[2] scanchain_183/module_data_in[3] scanchain_183/module_data_in[4]
+ scanchain_183/module_data_in[5] scanchain_183/module_data_in[6] scanchain_183/module_data_in[7]
+ scanchain_183/module_data_out[0] scanchain_183/module_data_out[1] scanchain_183/module_data_out[2]
+ scanchain_183/module_data_out[3] scanchain_183/module_data_out[4] scanchain_183/module_data_out[5]
+ scanchain_183/module_data_out[6] scanchain_183/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscan_controller io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18]
+ io_in[19] io_in[20] wb_clk_i io_in[8] io_in[9] io_in[21] io_in[22] io_in[23] io_in[24]
+ io_in[25] io_in[26] io_in[27] io_in[28] la_data_in[0] la_data_in[1] la_data_out[0]
+ la_data_in[3] la_data_in[2] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13]
+ io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20]
+ io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28]
+ io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[29] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35]
+ io_out[36] io_out[37] wb_rst_i scanchain_249/clk_out scanchain_000/clk_in scanchain_249/data_out
+ scanchain_000/data_in scanchain_000/latch_enable_in scan_controller/scan_select
+ io_in[11] io_out[10] vccd1 vssd1 scan_controller
Xscanchain_190 scanchain_190/clk_in scanchain_191/clk_in scanchain_190/data_in scanchain_191/data_in
+ scanchain_190/latch_enable_in scanchain_191/latch_enable_in scanchain_190/module_data_in[0]
+ scanchain_190/module_data_in[1] scanchain_190/module_data_in[2] scanchain_190/module_data_in[3]
+ scanchain_190/module_data_in[4] scanchain_190/module_data_in[5] scanchain_190/module_data_in[6]
+ scanchain_190/module_data_in[7] scanchain_190/module_data_out[0] scanchain_190/module_data_out[1]
+ scanchain_190/module_data_out[2] scanchain_190/module_data_out[3] scanchain_190/module_data_out[4]
+ scanchain_190/module_data_out[5] scanchain_190/module_data_out[6] scanchain_190/module_data_out[7]
+ scanchain_190/scan_select_in scanchain_191/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_195 scanchain_195/module_data_in[0] scanchain_195/module_data_in[1]
+ scanchain_195/module_data_in[2] scanchain_195/module_data_in[3] scanchain_195/module_data_in[4]
+ scanchain_195/module_data_in[5] scanchain_195/module_data_in[6] scanchain_195/module_data_in[7]
+ scanchain_195/module_data_out[0] scanchain_195/module_data_out[1] scanchain_195/module_data_out[2]
+ scanchain_195/module_data_out[3] scanchain_195/module_data_out[4] scanchain_195/module_data_out[5]
+ scanchain_195/module_data_out[6] scanchain_195/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_140 scanchain_140/module_data_in[0] scanchain_140/module_data_in[1]
+ scanchain_140/module_data_in[2] scanchain_140/module_data_in[3] scanchain_140/module_data_in[4]
+ scanchain_140/module_data_in[5] scanchain_140/module_data_in[6] scanchain_140/module_data_in[7]
+ scanchain_140/module_data_out[0] scanchain_140/module_data_out[1] scanchain_140/module_data_out[2]
+ scanchain_140/module_data_out[3] scanchain_140/module_data_out[4] scanchain_140/module_data_out[5]
+ scanchain_140/module_data_out[6] scanchain_140/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_151 scanchain_151/module_data_in[0] scanchain_151/module_data_in[1]
+ scanchain_151/module_data_in[2] scanchain_151/module_data_in[3] scanchain_151/module_data_in[4]
+ scanchain_151/module_data_in[5] scanchain_151/module_data_in[6] scanchain_151/module_data_in[7]
+ scanchain_151/module_data_out[0] scanchain_151/module_data_out[1] scanchain_151/module_data_out[2]
+ scanchain_151/module_data_out[3] scanchain_151/module_data_out[4] scanchain_151/module_data_out[5]
+ scanchain_151/module_data_out[6] scanchain_151/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_162 scanchain_162/module_data_in[0] scanchain_162/module_data_in[1]
+ scanchain_162/module_data_in[2] scanchain_162/module_data_in[3] scanchain_162/module_data_in[4]
+ scanchain_162/module_data_in[5] scanchain_162/module_data_in[6] scanchain_162/module_data_in[7]
+ scanchain_162/module_data_out[0] scanchain_162/module_data_out[1] scanchain_162/module_data_out[2]
+ scanchain_162/module_data_out[3] scanchain_162/module_data_out[4] scanchain_162/module_data_out[5]
+ scanchain_162/module_data_out[6] scanchain_162/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_173 scanchain_173/module_data_in[0] scanchain_173/module_data_in[1]
+ scanchain_173/module_data_in[2] scanchain_173/module_data_in[3] scanchain_173/module_data_in[4]
+ scanchain_173/module_data_in[5] scanchain_173/module_data_in[6] scanchain_173/module_data_in[7]
+ scanchain_173/module_data_out[0] scanchain_173/module_data_out[1] scanchain_173/module_data_out[2]
+ scanchain_173/module_data_out[3] scanchain_173/module_data_out[4] scanchain_173/module_data_out[5]
+ scanchain_173/module_data_out[6] scanchain_173/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_184 scanchain_184/module_data_in[0] scanchain_184/module_data_in[1]
+ scanchain_184/module_data_in[2] scanchain_184/module_data_in[3] scanchain_184/module_data_in[4]
+ scanchain_184/module_data_in[5] scanchain_184/module_data_in[6] scanchain_184/module_data_in[7]
+ scanchain_184/module_data_out[0] scanchain_184/module_data_out[1] scanchain_184/module_data_out[2]
+ scanchain_184/module_data_out[3] scanchain_184/module_data_out[4] scanchain_184/module_data_out[5]
+ scanchain_184/module_data_out[6] scanchain_184/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_019 scanchain_019/clk_in scanchain_020/clk_in scanchain_019/data_in scanchain_020/data_in
+ scanchain_019/latch_enable_in scanchain_020/latch_enable_in scanchain_019/module_data_in[0]
+ scanchain_019/module_data_in[1] scanchain_019/module_data_in[2] scanchain_019/module_data_in[3]
+ scanchain_019/module_data_in[4] scanchain_019/module_data_in[5] scanchain_019/module_data_in[6]
+ scanchain_019/module_data_in[7] scanchain_019/module_data_out[0] scanchain_019/module_data_out[1]
+ scanchain_019/module_data_out[2] scanchain_019/module_data_out[3] scanchain_019/module_data_out[4]
+ scanchain_019/module_data_out[5] scanchain_019/module_data_out[6] scanchain_019/module_data_out[7]
+ scanchain_019/scan_select_in scanchain_020/scan_select_in vccd1 vssd1 scanchain
Xscanchain_008 scanchain_008/clk_in scanchain_009/clk_in scanchain_008/data_in scanchain_009/data_in
+ scanchain_008/latch_enable_in scanchain_009/latch_enable_in aidan_McCoy_008/io_in[0]
+ aidan_McCoy_008/io_in[1] aidan_McCoy_008/io_in[2] aidan_McCoy_008/io_in[3] aidan_McCoy_008/io_in[4]
+ aidan_McCoy_008/io_in[5] aidan_McCoy_008/io_in[6] aidan_McCoy_008/io_in[7] aidan_McCoy_008/io_out[0]
+ aidan_McCoy_008/io_out[1] aidan_McCoy_008/io_out[2] aidan_McCoy_008/io_out[3] aidan_McCoy_008/io_out[4]
+ aidan_McCoy_008/io_out[5] aidan_McCoy_008/io_out[6] aidan_McCoy_008/io_out[7] scanchain_008/scan_select_in
+ scanchain_009/scan_select_in vccd1 vssd1 scanchain
Xuser_module_347688030570545747_021 scanchain_021/module_data_in[0] scanchain_021/module_data_in[1]
+ scanchain_021/module_data_in[2] scanchain_021/module_data_in[3] scanchain_021/module_data_in[4]
+ scanchain_021/module_data_in[5] scanchain_021/module_data_in[6] scanchain_021/module_data_in[7]
+ scanchain_021/module_data_out[0] scanchain_021/module_data_out[1] scanchain_021/module_data_out[2]
+ scanchain_021/module_data_out[3] scanchain_021/module_data_out[4] scanchain_021/module_data_out[5]
+ scanchain_021/module_data_out[6] scanchain_021/module_data_out[7] vccd1 vssd1 user_module_347688030570545747
Xscanchain_180 scanchain_180/clk_in scanchain_181/clk_in scanchain_180/data_in scanchain_181/data_in
+ scanchain_180/latch_enable_in scanchain_181/latch_enable_in scanchain_180/module_data_in[0]
+ scanchain_180/module_data_in[1] scanchain_180/module_data_in[2] scanchain_180/module_data_in[3]
+ scanchain_180/module_data_in[4] scanchain_180/module_data_in[5] scanchain_180/module_data_in[6]
+ scanchain_180/module_data_in[7] scanchain_180/module_data_out[0] scanchain_180/module_data_out[1]
+ scanchain_180/module_data_out[2] scanchain_180/module_data_out[3] scanchain_180/module_data_out[4]
+ scanchain_180/module_data_out[5] scanchain_180/module_data_out[6] scanchain_180/module_data_out[7]
+ scanchain_180/scan_select_in scanchain_181/scan_select_in vccd1 vssd1 scanchain
Xscanchain_191 scanchain_191/clk_in scanchain_192/clk_in scanchain_191/data_in scanchain_192/data_in
+ scanchain_191/latch_enable_in scanchain_192/latch_enable_in scanchain_191/module_data_in[0]
+ scanchain_191/module_data_in[1] scanchain_191/module_data_in[2] scanchain_191/module_data_in[3]
+ scanchain_191/module_data_in[4] scanchain_191/module_data_in[5] scanchain_191/module_data_in[6]
+ scanchain_191/module_data_in[7] scanchain_191/module_data_out[0] scanchain_191/module_data_out[1]
+ scanchain_191/module_data_out[2] scanchain_191/module_data_out[3] scanchain_191/module_data_out[4]
+ scanchain_191/module_data_out[5] scanchain_191/module_data_out[6] scanchain_191/module_data_out[7]
+ scanchain_191/scan_select_in scanchain_192/scan_select_in vccd1 vssd1 scanchain
Xuser_module_341535056611770964_196 scanchain_196/module_data_in[0] scanchain_196/module_data_in[1]
+ scanchain_196/module_data_in[2] scanchain_196/module_data_in[3] scanchain_196/module_data_in[4]
+ scanchain_196/module_data_in[5] scanchain_196/module_data_in[6] scanchain_196/module_data_in[7]
+ scanchain_196/module_data_out[0] scanchain_196/module_data_out[1] scanchain_196/module_data_out[2]
+ scanchain_196/module_data_out[3] scanchain_196/module_data_out[4] scanchain_196/module_data_out[5]
+ scanchain_196/module_data_out[6] scanchain_196/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xchase_the_beat_020 chase_the_beat_020/io_in[0] chase_the_beat_020/io_in[1] chase_the_beat_020/io_in[2]
+ chase_the_beat_020/io_in[3] chase_the_beat_020/io_in[4] chase_the_beat_020/io_in[5]
+ chase_the_beat_020/io_in[6] chase_the_beat_020/io_in[7] chase_the_beat_020/io_out[0]
+ chase_the_beat_020/io_out[1] chase_the_beat_020/io_out[2] chase_the_beat_020/io_out[3]
+ chase_the_beat_020/io_out[4] chase_the_beat_020/io_out[5] chase_the_beat_020/io_out[6]
+ chase_the_beat_020/io_out[7] vccd1 vssd1 chase_the_beat
Xuser_module_349047610915422802_065 scanchain_065/module_data_in[0] scanchain_065/module_data_in[1]
+ scanchain_065/module_data_in[2] scanchain_065/module_data_in[3] scanchain_065/module_data_in[4]
+ scanchain_065/module_data_in[5] scanchain_065/module_data_in[6] scanchain_065/module_data_in[7]
+ scanchain_065/module_data_out[0] scanchain_065/module_data_out[1] scanchain_065/module_data_out[2]
+ scanchain_065/module_data_out[3] scanchain_065/module_data_out[4] scanchain_065/module_data_out[5]
+ scanchain_065/module_data_out[6] scanchain_065/module_data_out[7] vccd1 vssd1 user_module_349047610915422802
Xuser_module_341535056611770964_130 scanchain_130/module_data_in[0] scanchain_130/module_data_in[1]
+ scanchain_130/module_data_in[2] scanchain_130/module_data_in[3] scanchain_130/module_data_in[4]
+ scanchain_130/module_data_in[5] scanchain_130/module_data_in[6] scanchain_130/module_data_in[7]
+ scanchain_130/module_data_out[0] scanchain_130/module_data_out[1] scanchain_130/module_data_out[2]
+ scanchain_130/module_data_out[3] scanchain_130/module_data_out[4] scanchain_130/module_data_out[5]
+ scanchain_130/module_data_out[6] scanchain_130/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_141 scanchain_141/module_data_in[0] scanchain_141/module_data_in[1]
+ scanchain_141/module_data_in[2] scanchain_141/module_data_in[3] scanchain_141/module_data_in[4]
+ scanchain_141/module_data_in[5] scanchain_141/module_data_in[6] scanchain_141/module_data_in[7]
+ scanchain_141/module_data_out[0] scanchain_141/module_data_out[1] scanchain_141/module_data_out[2]
+ scanchain_141/module_data_out[3] scanchain_141/module_data_out[4] scanchain_141/module_data_out[5]
+ scanchain_141/module_data_out[6] scanchain_141/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_163 scanchain_163/module_data_in[0] scanchain_163/module_data_in[1]
+ scanchain_163/module_data_in[2] scanchain_163/module_data_in[3] scanchain_163/module_data_in[4]
+ scanchain_163/module_data_in[5] scanchain_163/module_data_in[6] scanchain_163/module_data_in[7]
+ scanchain_163/module_data_out[0] scanchain_163/module_data_out[1] scanchain_163/module_data_out[2]
+ scanchain_163/module_data_out[3] scanchain_163/module_data_out[4] scanchain_163/module_data_out[5]
+ scanchain_163/module_data_out[6] scanchain_163/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_152 scanchain_152/module_data_in[0] scanchain_152/module_data_in[1]
+ scanchain_152/module_data_in[2] scanchain_152/module_data_in[3] scanchain_152/module_data_in[4]
+ scanchain_152/module_data_in[5] scanchain_152/module_data_in[6] scanchain_152/module_data_in[7]
+ scanchain_152/module_data_out[0] scanchain_152/module_data_out[1] scanchain_152/module_data_out[2]
+ scanchain_152/module_data_out[3] scanchain_152/module_data_out[4] scanchain_152/module_data_out[5]
+ scanchain_152/module_data_out[6] scanchain_152/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_174 scanchain_174/module_data_in[0] scanchain_174/module_data_in[1]
+ scanchain_174/module_data_in[2] scanchain_174/module_data_in[3] scanchain_174/module_data_in[4]
+ scanchain_174/module_data_in[5] scanchain_174/module_data_in[6] scanchain_174/module_data_in[7]
+ scanchain_174/module_data_out[0] scanchain_174/module_data_out[1] scanchain_174/module_data_out[2]
+ scanchain_174/module_data_out[3] scanchain_174/module_data_out[4] scanchain_174/module_data_out[5]
+ scanchain_174/module_data_out[6] scanchain_174/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_185 scanchain_185/module_data_in[0] scanchain_185/module_data_in[1]
+ scanchain_185/module_data_in[2] scanchain_185/module_data_in[3] scanchain_185/module_data_in[4]
+ scanchain_185/module_data_in[5] scanchain_185/module_data_in[6] scanchain_185/module_data_in[7]
+ scanchain_185/module_data_out[0] scanchain_185/module_data_out[1] scanchain_185/module_data_out[2]
+ scanchain_185/module_data_out[3] scanchain_185/module_data_out[4] scanchain_185/module_data_out[5]
+ scanchain_185/module_data_out[6] scanchain_185/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xscanchain_009 scanchain_009/clk_in scanchain_010/clk_in scanchain_009/data_in scanchain_010/data_in
+ scanchain_009/latch_enable_in scanchain_010/latch_enable_in scanchain_009/module_data_in[0]
+ scanchain_009/module_data_in[1] scanchain_009/module_data_in[2] scanchain_009/module_data_in[3]
+ scanchain_009/module_data_in[4] scanchain_009/module_data_in[5] scanchain_009/module_data_in[6]
+ scanchain_009/module_data_in[7] scanchain_009/module_data_out[0] scanchain_009/module_data_out[1]
+ scanchain_009/module_data_out[2] scanchain_009/module_data_out[3] scanchain_009/module_data_out[4]
+ scanchain_009/module_data_out[5] scanchain_009/module_data_out[6] scanchain_009/module_data_out[7]
+ scanchain_009/scan_select_in scanchain_010/scan_select_in vccd1 vssd1 scanchain
Xnavray_top_070 navray_top_070/io_in[0] navray_top_070/io_in[1] navray_top_070/io_in[2]
+ navray_top_070/io_in[3] navray_top_070/io_in[4] navray_top_070/io_in[5] navray_top_070/io_in[6]
+ navray_top_070/io_in[7] navray_top_070/io_out[0] navray_top_070/io_out[1] navray_top_070/io_out[2]
+ navray_top_070/io_out[3] navray_top_070/io_out[4] navray_top_070/io_out[5] navray_top_070/io_out[6]
+ navray_top_070/io_out[7] vccd1 vssd1 navray_top
Xgatecat_fpga_top_089 gatecat_fpga_top_089/io_in[0] gatecat_fpga_top_089/io_in[1]
+ gatecat_fpga_top_089/io_in[2] gatecat_fpga_top_089/io_in[3] gatecat_fpga_top_089/io_in[4]
+ gatecat_fpga_top_089/io_in[5] gatecat_fpga_top_089/io_in[6] gatecat_fpga_top_089/io_in[7]
+ gatecat_fpga_top_089/io_out[0] gatecat_fpga_top_089/io_out[1] gatecat_fpga_top_089/io_out[2]
+ gatecat_fpga_top_089/io_out[3] gatecat_fpga_top_089/io_out[4] gatecat_fpga_top_089/io_out[5]
+ gatecat_fpga_top_089/io_out[6] gatecat_fpga_top_089/io_out[7] vccd1 vssd1 gatecat_fpga_top
Xscanchain_181 scanchain_181/clk_in scanchain_182/clk_in scanchain_181/data_in scanchain_182/data_in
+ scanchain_181/latch_enable_in scanchain_182/latch_enable_in scanchain_181/module_data_in[0]
+ scanchain_181/module_data_in[1] scanchain_181/module_data_in[2] scanchain_181/module_data_in[3]
+ scanchain_181/module_data_in[4] scanchain_181/module_data_in[5] scanchain_181/module_data_in[6]
+ scanchain_181/module_data_in[7] scanchain_181/module_data_out[0] scanchain_181/module_data_out[1]
+ scanchain_181/module_data_out[2] scanchain_181/module_data_out[3] scanchain_181/module_data_out[4]
+ scanchain_181/module_data_out[5] scanchain_181/module_data_out[6] scanchain_181/module_data_out[7]
+ scanchain_181/scan_select_in scanchain_182/scan_select_in vccd1 vssd1 scanchain
Xscanchain_170 scanchain_170/clk_in scanchain_171/clk_in scanchain_170/data_in scanchain_171/data_in
+ scanchain_170/latch_enable_in scanchain_171/latch_enable_in scanchain_170/module_data_in[0]
+ scanchain_170/module_data_in[1] scanchain_170/module_data_in[2] scanchain_170/module_data_in[3]
+ scanchain_170/module_data_in[4] scanchain_170/module_data_in[5] scanchain_170/module_data_in[6]
+ scanchain_170/module_data_in[7] scanchain_170/module_data_out[0] scanchain_170/module_data_out[1]
+ scanchain_170/module_data_out[2] scanchain_170/module_data_out[3] scanchain_170/module_data_out[4]
+ scanchain_170/module_data_out[5] scanchain_170/module_data_out[6] scanchain_170/module_data_out[7]
+ scanchain_170/scan_select_in scanchain_171/scan_select_in vccd1 vssd1 scanchain
Xscanchain_192 scanchain_192/clk_in scanchain_193/clk_in scanchain_192/data_in scanchain_193/data_in
+ scanchain_192/latch_enable_in scanchain_193/latch_enable_in scanchain_192/module_data_in[0]
+ scanchain_192/module_data_in[1] scanchain_192/module_data_in[2] scanchain_192/module_data_in[3]
+ scanchain_192/module_data_in[4] scanchain_192/module_data_in[5] scanchain_192/module_data_in[6]
+ scanchain_192/module_data_in[7] scanchain_192/module_data_out[0] scanchain_192/module_data_out[1]
+ scanchain_192/module_data_out[2] scanchain_192/module_data_out[3] scanchain_192/module_data_out[4]
+ scanchain_192/module_data_out[5] scanchain_192/module_data_out[6] scanchain_192/module_data_out[7]
+ scanchain_192/scan_select_in scanchain_193/scan_select_in vccd1 vssd1 scanchain
Xthezoq2_yafpga_038 thezoq2_yafpga_038/io_in[0] thezoq2_yafpga_038/io_in[1] thezoq2_yafpga_038/io_in[2]
+ thezoq2_yafpga_038/io_in[3] thezoq2_yafpga_038/io_in[4] thezoq2_yafpga_038/io_in[5]
+ thezoq2_yafpga_038/io_in[6] thezoq2_yafpga_038/io_in[7] thezoq2_yafpga_038/io_out[0]
+ thezoq2_yafpga_038/io_out[1] thezoq2_yafpga_038/io_out[2] thezoq2_yafpga_038/io_out[3]
+ thezoq2_yafpga_038/io_out[4] thezoq2_yafpga_038/io_out[5] thezoq2_yafpga_038/io_out[6]
+ thezoq2_yafpga_038/io_out[7] vccd1 vssd1 thezoq2_yafpga
Xuser_module_340318610245288530_080 scanchain_080/module_data_in[0] scanchain_080/module_data_in[1]
+ scanchain_080/module_data_in[2] scanchain_080/module_data_in[3] scanchain_080/module_data_in[4]
+ scanchain_080/module_data_in[5] scanchain_080/module_data_in[6] scanchain_080/module_data_in[7]
+ scanchain_080/module_data_out[0] scanchain_080/module_data_out[1] scanchain_080/module_data_out[2]
+ scanchain_080/module_data_out[3] scanchain_080/module_data_out[4] scanchain_080/module_data_out[5]
+ scanchain_080/module_data_out[6] scanchain_080/module_data_out[7] vccd1 vssd1 user_module_340318610245288530
Xchrisruk_matrix_003 chrisruk_matrix_003/io_in[0] chrisruk_matrix_003/io_in[1] chrisruk_matrix_003/io_in[2]
+ chrisruk_matrix_003/io_in[3] chrisruk_matrix_003/io_in[4] chrisruk_matrix_003/io_in[5]
+ chrisruk_matrix_003/io_in[6] chrisruk_matrix_003/io_in[7] chrisruk_matrix_003/io_out[0]
+ chrisruk_matrix_003/io_out[1] chrisruk_matrix_003/io_out[2] chrisruk_matrix_003/io_out[3]
+ chrisruk_matrix_003/io_out[4] chrisruk_matrix_003/io_out[5] chrisruk_matrix_003/io_out[6]
+ chrisruk_matrix_003/io_out[7] vccd1 vssd1 chrisruk_matrix
Xuser_module_348540666182107731_063 scanchain_063/module_data_in[0] scanchain_063/module_data_in[1]
+ scanchain_063/module_data_in[2] scanchain_063/module_data_in[3] scanchain_063/module_data_in[4]
+ scanchain_063/module_data_in[5] scanchain_063/module_data_in[6] scanchain_063/module_data_in[7]
+ scanchain_063/module_data_out[0] scanchain_063/module_data_out[1] scanchain_063/module_data_out[2]
+ scanchain_063/module_data_out[3] scanchain_063/module_data_out[4] scanchain_063/module_data_out[5]
+ scanchain_063/module_data_out[6] scanchain_063/module_data_out[7] vccd1 vssd1 user_module_348540666182107731
Xuser_module_347787021138264660_010 scanchain_010/module_data_in[0] scanchain_010/module_data_in[1]
+ scanchain_010/module_data_in[2] scanchain_010/module_data_in[3] scanchain_010/module_data_in[4]
+ scanchain_010/module_data_in[5] scanchain_010/module_data_in[6] scanchain_010/module_data_in[7]
+ scanchain_010/module_data_out[0] scanchain_010/module_data_out[1] scanchain_010/module_data_out[2]
+ scanchain_010/module_data_out[3] scanchain_010/module_data_out[4] scanchain_010/module_data_out[5]
+ scanchain_010/module_data_out[6] scanchain_010/module_data_out[7] vccd1 vssd1 user_module_347787021138264660
Xuser_module_341535056611770964_120 scanchain_120/module_data_in[0] scanchain_120/module_data_in[1]
+ scanchain_120/module_data_in[2] scanchain_120/module_data_in[3] scanchain_120/module_data_in[4]
+ scanchain_120/module_data_in[5] scanchain_120/module_data_in[6] scanchain_120/module_data_in[7]
+ scanchain_120/module_data_out[0] scanchain_120/module_data_out[1] scanchain_120/module_data_out[2]
+ scanchain_120/module_data_out[3] scanchain_120/module_data_out[4] scanchain_120/module_data_out[5]
+ scanchain_120/module_data_out[6] scanchain_120/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_131 scanchain_131/module_data_in[0] scanchain_131/module_data_in[1]
+ scanchain_131/module_data_in[2] scanchain_131/module_data_in[3] scanchain_131/module_data_in[4]
+ scanchain_131/module_data_in[5] scanchain_131/module_data_in[6] scanchain_131/module_data_in[7]
+ scanchain_131/module_data_out[0] scanchain_131/module_data_out[1] scanchain_131/module_data_out[2]
+ scanchain_131/module_data_out[3] scanchain_131/module_data_out[4] scanchain_131/module_data_out[5]
+ scanchain_131/module_data_out[6] scanchain_131/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_197 scanchain_197/module_data_in[0] scanchain_197/module_data_in[1]
+ scanchain_197/module_data_in[2] scanchain_197/module_data_in[3] scanchain_197/module_data_in[4]
+ scanchain_197/module_data_in[5] scanchain_197/module_data_in[6] scanchain_197/module_data_in[7]
+ scanchain_197/module_data_out[0] scanchain_197/module_data_out[1] scanchain_197/module_data_out[2]
+ scanchain_197/module_data_out[3] scanchain_197/module_data_out[4] scanchain_197/module_data_out[5]
+ scanchain_197/module_data_out[6] scanchain_197/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xcpldcpu_TrainLED2top_076 scanchain_076/module_data_in[0] scanchain_076/module_data_in[1]
+ scanchain_076/module_data_in[2] scanchain_076/module_data_in[3] scanchain_076/module_data_in[4]
+ scanchain_076/module_data_in[5] scanchain_076/module_data_in[6] scanchain_076/module_data_in[7]
+ scanchain_076/module_data_out[0] scanchain_076/module_data_out[1] scanchain_076/module_data_out[2]
+ scanchain_076/module_data_out[3] scanchain_076/module_data_out[4] scanchain_076/module_data_out[5]
+ scanchain_076/module_data_out[6] scanchain_076/module_data_out[7] vccd1 vssd1 cpldcpu_TrainLED2top
Xuser_module_341535056611770964_142 scanchain_142/module_data_in[0] scanchain_142/module_data_in[1]
+ scanchain_142/module_data_in[2] scanchain_142/module_data_in[3] scanchain_142/module_data_in[4]
+ scanchain_142/module_data_in[5] scanchain_142/module_data_in[6] scanchain_142/module_data_in[7]
+ scanchain_142/module_data_out[0] scanchain_142/module_data_out[1] scanchain_142/module_data_out[2]
+ scanchain_142/module_data_out[3] scanchain_142/module_data_out[4] scanchain_142/module_data_out[5]
+ scanchain_142/module_data_out[6] scanchain_142/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_164 scanchain_164/module_data_in[0] scanchain_164/module_data_in[1]
+ scanchain_164/module_data_in[2] scanchain_164/module_data_in[3] scanchain_164/module_data_in[4]
+ scanchain_164/module_data_in[5] scanchain_164/module_data_in[6] scanchain_164/module_data_in[7]
+ scanchain_164/module_data_out[0] scanchain_164/module_data_out[1] scanchain_164/module_data_out[2]
+ scanchain_164/module_data_out[3] scanchain_164/module_data_out[4] scanchain_164/module_data_out[5]
+ scanchain_164/module_data_out[6] scanchain_164/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_153 scanchain_153/module_data_in[0] scanchain_153/module_data_in[1]
+ scanchain_153/module_data_in[2] scanchain_153/module_data_in[3] scanchain_153/module_data_in[4]
+ scanchain_153/module_data_in[5] scanchain_153/module_data_in[6] scanchain_153/module_data_in[7]
+ scanchain_153/module_data_out[0] scanchain_153/module_data_out[1] scanchain_153/module_data_out[2]
+ scanchain_153/module_data_out[3] scanchain_153/module_data_out[4] scanchain_153/module_data_out[5]
+ scanchain_153/module_data_out[6] scanchain_153/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_175 scanchain_175/module_data_in[0] scanchain_175/module_data_in[1]
+ scanchain_175/module_data_in[2] scanchain_175/module_data_in[3] scanchain_175/module_data_in[4]
+ scanchain_175/module_data_in[5] scanchain_175/module_data_in[6] scanchain_175/module_data_in[7]
+ scanchain_175/module_data_out[0] scanchain_175/module_data_out[1] scanchain_175/module_data_out[2]
+ scanchain_175/module_data_out[3] scanchain_175/module_data_out[4] scanchain_175/module_data_out[5]
+ scanchain_175/module_data_out[6] scanchain_175/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_186 scanchain_186/module_data_in[0] scanchain_186/module_data_in[1]
+ scanchain_186/module_data_in[2] scanchain_186/module_data_in[3] scanchain_186/module_data_in[4]
+ scanchain_186/module_data_in[5] scanchain_186/module_data_in[6] scanchain_186/module_data_in[7]
+ scanchain_186/module_data_out[0] scanchain_186/module_data_out[1] scanchain_186/module_data_out[2]
+ scanchain_186/module_data_out[3] scanchain_186/module_data_out[4] scanchain_186/module_data_out[5]
+ scanchain_186/module_data_out[6] scanchain_186/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_347690870424732244_012 scanchain_012/module_data_in[0] scanchain_012/module_data_in[1]
+ scanchain_012/module_data_in[2] scanchain_012/module_data_in[3] scanchain_012/module_data_in[4]
+ scanchain_012/module_data_in[5] scanchain_012/module_data_in[6] scanchain_012/module_data_in[7]
+ scanchain_012/module_data_out[0] scanchain_012/module_data_out[1] scanchain_012/module_data_out[2]
+ scanchain_012/module_data_out[3] scanchain_012/module_data_out[4] scanchain_012/module_data_out[5]
+ scanchain_012/module_data_out[6] scanchain_012/module_data_out[7] vccd1 vssd1 user_module_347690870424732244
Xuser_module_348787952842703444_095 scanchain_095/module_data_in[0] scanchain_095/module_data_in[1]
+ scanchain_095/module_data_in[2] scanchain_095/module_data_in[3] scanchain_095/module_data_in[4]
+ scanchain_095/module_data_in[5] scanchain_095/module_data_in[6] scanchain_095/module_data_in[7]
+ scanchain_095/module_data_out[0] scanchain_095/module_data_out[1] scanchain_095/module_data_out[2]
+ scanchain_095/module_data_out[3] scanchain_095/module_data_out[4] scanchain_095/module_data_out[5]
+ scanchain_095/module_data_out[6] scanchain_095/module_data_out[7] vccd1 vssd1 user_module_348787952842703444
Xscanchain_182 scanchain_182/clk_in scanchain_183/clk_in scanchain_182/data_in scanchain_183/data_in
+ scanchain_182/latch_enable_in scanchain_183/latch_enable_in scanchain_182/module_data_in[0]
+ scanchain_182/module_data_in[1] scanchain_182/module_data_in[2] scanchain_182/module_data_in[3]
+ scanchain_182/module_data_in[4] scanchain_182/module_data_in[5] scanchain_182/module_data_in[6]
+ scanchain_182/module_data_in[7] scanchain_182/module_data_out[0] scanchain_182/module_data_out[1]
+ scanchain_182/module_data_out[2] scanchain_182/module_data_out[3] scanchain_182/module_data_out[4]
+ scanchain_182/module_data_out[5] scanchain_182/module_data_out[6] scanchain_182/module_data_out[7]
+ scanchain_182/scan_select_in scanchain_183/scan_select_in vccd1 vssd1 scanchain
Xscanchain_160 scanchain_160/clk_in scanchain_161/clk_in scanchain_160/data_in scanchain_161/data_in
+ scanchain_160/latch_enable_in scanchain_161/latch_enable_in scanchain_160/module_data_in[0]
+ scanchain_160/module_data_in[1] scanchain_160/module_data_in[2] scanchain_160/module_data_in[3]
+ scanchain_160/module_data_in[4] scanchain_160/module_data_in[5] scanchain_160/module_data_in[6]
+ scanchain_160/module_data_in[7] scanchain_160/module_data_out[0] scanchain_160/module_data_out[1]
+ scanchain_160/module_data_out[2] scanchain_160/module_data_out[3] scanchain_160/module_data_out[4]
+ scanchain_160/module_data_out[5] scanchain_160/module_data_out[6] scanchain_160/module_data_out[7]
+ scanchain_160/scan_select_in scanchain_161/scan_select_in vccd1 vssd1 scanchain
Xscanchain_171 scanchain_171/clk_in scanchain_172/clk_in scanchain_171/data_in scanchain_172/data_in
+ scanchain_171/latch_enable_in scanchain_172/latch_enable_in scanchain_171/module_data_in[0]
+ scanchain_171/module_data_in[1] scanchain_171/module_data_in[2] scanchain_171/module_data_in[3]
+ scanchain_171/module_data_in[4] scanchain_171/module_data_in[5] scanchain_171/module_data_in[6]
+ scanchain_171/module_data_in[7] scanchain_171/module_data_out[0] scanchain_171/module_data_out[1]
+ scanchain_171/module_data_out[2] scanchain_171/module_data_out[3] scanchain_171/module_data_out[4]
+ scanchain_171/module_data_out[5] scanchain_171/module_data_out[6] scanchain_171/module_data_out[7]
+ scanchain_171/scan_select_in scanchain_172/scan_select_in vccd1 vssd1 scanchain
Xscanchain_193 scanchain_193/clk_in scanchain_194/clk_in scanchain_193/data_in scanchain_194/data_in
+ scanchain_193/latch_enable_in scanchain_194/latch_enable_in scanchain_193/module_data_in[0]
+ scanchain_193/module_data_in[1] scanchain_193/module_data_in[2] scanchain_193/module_data_in[3]
+ scanchain_193/module_data_in[4] scanchain_193/module_data_in[5] scanchain_193/module_data_in[6]
+ scanchain_193/module_data_in[7] scanchain_193/module_data_out[0] scanchain_193/module_data_out[1]
+ scanchain_193/module_data_out[2] scanchain_193/module_data_out[3] scanchain_193/module_data_out[4]
+ scanchain_193/module_data_out[5] scanchain_193/module_data_out[6] scanchain_193/module_data_out[7]
+ scanchain_193/scan_select_in scanchain_194/scan_select_in vccd1 vssd1 scanchain
Xuser_module_348242239268323922_037 scanchain_037/module_data_in[0] scanchain_037/module_data_in[1]
+ scanchain_037/module_data_in[2] scanchain_037/module_data_in[3] scanchain_037/module_data_in[4]
+ scanchain_037/module_data_in[5] scanchain_037/module_data_in[6] scanchain_037/module_data_in[7]
+ scanchain_037/module_data_out[0] scanchain_037/module_data_out[1] scanchain_037/module_data_out[2]
+ scanchain_037/module_data_out[3] scanchain_037/module_data_out[4] scanchain_037/module_data_out[5]
+ scanchain_037/module_data_out[6] scanchain_037/module_data_out[7] vccd1 vssd1 user_module_348242239268323922
Xuser_module_341535056611770964_198 scanchain_198/module_data_in[0] scanchain_198/module_data_in[1]
+ scanchain_198/module_data_in[2] scanchain_198/module_data_in[3] scanchain_198/module_data_in[4]
+ scanchain_198/module_data_in[5] scanchain_198/module_data_in[6] scanchain_198/module_data_in[7]
+ scanchain_198/module_data_out[0] scanchain_198/module_data_out[1] scanchain_198/module_data_out[2]
+ scanchain_198/module_data_out[3] scanchain_198/module_data_out[4] scanchain_198/module_data_out[5]
+ scanchain_198/module_data_out[6] scanchain_198/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_110 scanchain_110/module_data_in[0] scanchain_110/module_data_in[1]
+ scanchain_110/module_data_in[2] scanchain_110/module_data_in[3] scanchain_110/module_data_in[4]
+ scanchain_110/module_data_in[5] scanchain_110/module_data_in[6] scanchain_110/module_data_in[7]
+ scanchain_110/module_data_out[0] scanchain_110/module_data_out[1] scanchain_110/module_data_out[2]
+ scanchain_110/module_data_out[3] scanchain_110/module_data_out[4] scanchain_110/module_data_out[5]
+ scanchain_110/module_data_out[6] scanchain_110/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_121 scanchain_121/module_data_in[0] scanchain_121/module_data_in[1]
+ scanchain_121/module_data_in[2] scanchain_121/module_data_in[3] scanchain_121/module_data_in[4]
+ scanchain_121/module_data_in[5] scanchain_121/module_data_in[6] scanchain_121/module_data_in[7]
+ scanchain_121/module_data_out[0] scanchain_121/module_data_out[1] scanchain_121/module_data_out[2]
+ scanchain_121/module_data_out[3] scanchain_121/module_data_out[4] scanchain_121/module_data_out[5]
+ scanchain_121/module_data_out[6] scanchain_121/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_132 scanchain_132/module_data_in[0] scanchain_132/module_data_in[1]
+ scanchain_132/module_data_in[2] scanchain_132/module_data_in[3] scanchain_132/module_data_in[4]
+ scanchain_132/module_data_in[5] scanchain_132/module_data_in[6] scanchain_132/module_data_in[7]
+ scanchain_132/module_data_out[0] scanchain_132/module_data_out[1] scanchain_132/module_data_out[2]
+ scanchain_132/module_data_out[3] scanchain_132/module_data_out[4] scanchain_132/module_data_out[5]
+ scanchain_132/module_data_out[6] scanchain_132/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_143 scanchain_143/module_data_in[0] scanchain_143/module_data_in[1]
+ scanchain_143/module_data_in[2] scanchain_143/module_data_in[3] scanchain_143/module_data_in[4]
+ scanchain_143/module_data_in[5] scanchain_143/module_data_in[6] scanchain_143/module_data_in[7]
+ scanchain_143/module_data_out[0] scanchain_143/module_data_out[1] scanchain_143/module_data_out[2]
+ scanchain_143/module_data_out[3] scanchain_143/module_data_out[4] scanchain_143/module_data_out[5]
+ scanchain_143/module_data_out[6] scanchain_143/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_165 scanchain_165/module_data_in[0] scanchain_165/module_data_in[1]
+ scanchain_165/module_data_in[2] scanchain_165/module_data_in[3] scanchain_165/module_data_in[4]
+ scanchain_165/module_data_in[5] scanchain_165/module_data_in[6] scanchain_165/module_data_in[7]
+ scanchain_165/module_data_out[0] scanchain_165/module_data_out[1] scanchain_165/module_data_out[2]
+ scanchain_165/module_data_out[3] scanchain_165/module_data_out[4] scanchain_165/module_data_out[5]
+ scanchain_165/module_data_out[6] scanchain_165/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_154 scanchain_154/module_data_in[0] scanchain_154/module_data_in[1]
+ scanchain_154/module_data_in[2] scanchain_154/module_data_in[3] scanchain_154/module_data_in[4]
+ scanchain_154/module_data_in[5] scanchain_154/module_data_in[6] scanchain_154/module_data_in[7]
+ scanchain_154/module_data_out[0] scanchain_154/module_data_out[1] scanchain_154/module_data_out[2]
+ scanchain_154/module_data_out[3] scanchain_154/module_data_out[4] scanchain_154/module_data_out[5]
+ scanchain_154/module_data_out[6] scanchain_154/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_176 scanchain_176/module_data_in[0] scanchain_176/module_data_in[1]
+ scanchain_176/module_data_in[2] scanchain_176/module_data_in[3] scanchain_176/module_data_in[4]
+ scanchain_176/module_data_in[5] scanchain_176/module_data_in[6] scanchain_176/module_data_in[7]
+ scanchain_176/module_data_out[0] scanchain_176/module_data_out[1] scanchain_176/module_data_out[2]
+ scanchain_176/module_data_out[3] scanchain_176/module_data_out[4] scanchain_176/module_data_out[5]
+ scanchain_176/module_data_out[6] scanchain_176/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
Xuser_module_341535056611770964_187 scanchain_187/module_data_in[0] scanchain_187/module_data_in[1]
+ scanchain_187/module_data_in[2] scanchain_187/module_data_in[3] scanchain_187/module_data_in[4]
+ scanchain_187/module_data_in[5] scanchain_187/module_data_in[6] scanchain_187/module_data_in[7]
+ scanchain_187/module_data_out[0] scanchain_187/module_data_out[1] scanchain_187/module_data_out[2]
+ scanchain_187/module_data_out[3] scanchain_187/module_data_out[4] scanchain_187/module_data_out[5]
+ scanchain_187/module_data_out[6] scanchain_187/module_data_out[7] vccd1 vssd1 user_module_341535056611770964
.ends

