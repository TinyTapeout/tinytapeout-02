VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tomkeddie_top_tto
  CLASS BLOCK ;
  FOREIGN tomkeddie_top_tto ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 120.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 2.000 4.040 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 2.000 11.520 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.000 19.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.000 26.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.000 33.960 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.000 41.440 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.000 48.920 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.000 56.400 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 2.000 63.880 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 2.000 71.360 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.000 78.840 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.000 86.320 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.000 93.800 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.000 101.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 2.000 108.760 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.000 116.240 ;
    END
  END io_out[7]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.590 5.200 16.190 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.330 5.200 35.930 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.070 5.200 55.670 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.810 5.200 75.410 114.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.460 5.200 26.060 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.200 5.200 45.800 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.940 5.200 65.540 114.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 84.180 114.325 ;
      LAYER met1 ;
        RECT 2.830 1.060 85.490 114.480 ;
      LAYER met2 ;
        RECT 2.850 0.835 85.470 116.125 ;
      LAYER met3 ;
        RECT 2.400 115.240 85.495 116.105 ;
        RECT 2.000 109.160 85.495 115.240 ;
        RECT 2.400 107.760 85.495 109.160 ;
        RECT 2.000 101.680 85.495 107.760 ;
        RECT 2.400 100.280 85.495 101.680 ;
        RECT 2.000 94.200 85.495 100.280 ;
        RECT 2.400 92.800 85.495 94.200 ;
        RECT 2.000 86.720 85.495 92.800 ;
        RECT 2.400 85.320 85.495 86.720 ;
        RECT 2.000 79.240 85.495 85.320 ;
        RECT 2.400 77.840 85.495 79.240 ;
        RECT 2.000 71.760 85.495 77.840 ;
        RECT 2.400 70.360 85.495 71.760 ;
        RECT 2.000 64.280 85.495 70.360 ;
        RECT 2.400 62.880 85.495 64.280 ;
        RECT 2.000 56.800 85.495 62.880 ;
        RECT 2.400 55.400 85.495 56.800 ;
        RECT 2.000 49.320 85.495 55.400 ;
        RECT 2.400 47.920 85.495 49.320 ;
        RECT 2.000 41.840 85.495 47.920 ;
        RECT 2.400 40.440 85.495 41.840 ;
        RECT 2.000 34.360 85.495 40.440 ;
        RECT 2.400 32.960 85.495 34.360 ;
        RECT 2.000 26.880 85.495 32.960 ;
        RECT 2.400 25.480 85.495 26.880 ;
        RECT 2.000 19.400 85.495 25.480 ;
        RECT 2.400 18.000 85.495 19.400 ;
        RECT 2.000 11.920 85.495 18.000 ;
        RECT 2.400 10.520 85.495 11.920 ;
        RECT 2.000 4.440 85.495 10.520 ;
        RECT 2.400 3.040 85.495 4.440 ;
        RECT 2.000 0.855 85.495 3.040 ;
      LAYER met4 ;
        RECT 5.815 4.800 14.190 110.665 ;
        RECT 16.590 4.800 24.060 110.665 ;
        RECT 26.460 4.800 33.930 110.665 ;
        RECT 36.330 4.800 43.800 110.665 ;
        RECT 46.200 4.800 53.670 110.665 ;
        RECT 56.070 4.800 63.540 110.665 ;
        RECT 65.940 4.800 73.410 110.665 ;
        RECT 75.810 4.800 80.665 110.665 ;
        RECT 5.815 0.855 80.665 4.800 ;
  END
END tomkeddie_top_tto
END LIBRARY

