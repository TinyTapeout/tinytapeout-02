VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 120.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 118.000 1.290 120.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 118.000 24.290 120.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 118.000 26.590 120.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 118.000 28.890 120.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 118.000 31.190 120.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 118.000 33.490 120.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 118.000 35.790 120.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 118.000 38.090 120.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 118.000 40.390 120.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 118.000 42.690 120.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 118.000 44.990 120.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 118.000 3.590 120.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 118.000 47.290 120.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 118.000 49.590 120.000 ;
    END
  END io_in[21]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 118.000 5.890 120.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 118.000 8.190 120.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 118.000 10.490 120.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 118.000 12.790 120.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 118.000 15.090 120.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 118.000 17.390 120.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 118.000 19.690 120.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 118.000 21.990 120.000 ;
    END
  END io_in[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 118.000 51.890 120.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 118.000 74.890 120.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 118.000 77.190 120.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 118.000 79.490 120.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 118.000 81.790 120.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 118.000 84.090 120.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 118.000 86.390 120.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 118.000 88.690 120.000 ;
    END
  END io_out[16]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 118.000 54.190 120.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 118.000 56.490 120.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 118.000 58.790 120.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 118.000 61.090 120.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 118.000 63.390 120.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 118.000 65.690 120.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 118.000 67.990 120.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 118.000 70.290 120.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 118.000 72.590 120.000 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.590 5.200 16.190 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.330 5.200 35.930 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.070 5.200 55.670 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.810 5.200 75.410 114.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.460 5.200 26.060 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.200 5.200 45.800 114.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.940 5.200 65.540 114.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 84.180 114.325 ;
      LAYER met1 ;
        RECT 0.070 5.200 88.710 117.940 ;
      LAYER met2 ;
        RECT 0.100 117.720 0.730 119.525 ;
        RECT 1.570 117.720 3.030 119.525 ;
        RECT 3.870 117.720 5.330 119.525 ;
        RECT 6.170 117.720 7.630 119.525 ;
        RECT 8.470 117.720 9.930 119.525 ;
        RECT 10.770 117.720 12.230 119.525 ;
        RECT 13.070 117.720 14.530 119.525 ;
        RECT 15.370 117.720 16.830 119.525 ;
        RECT 17.670 117.720 19.130 119.525 ;
        RECT 19.970 117.720 21.430 119.525 ;
        RECT 22.270 117.720 23.730 119.525 ;
        RECT 24.570 117.720 26.030 119.525 ;
        RECT 26.870 117.720 28.330 119.525 ;
        RECT 29.170 117.720 30.630 119.525 ;
        RECT 31.470 117.720 32.930 119.525 ;
        RECT 33.770 117.720 35.230 119.525 ;
        RECT 36.070 117.720 37.530 119.525 ;
        RECT 38.370 117.720 39.830 119.525 ;
        RECT 40.670 117.720 42.130 119.525 ;
        RECT 42.970 117.720 44.430 119.525 ;
        RECT 45.270 117.720 46.730 119.525 ;
        RECT 47.570 117.720 49.030 119.525 ;
        RECT 49.870 117.720 51.330 119.525 ;
        RECT 52.170 117.720 53.630 119.525 ;
        RECT 54.470 117.720 55.930 119.525 ;
        RECT 56.770 117.720 58.230 119.525 ;
        RECT 59.070 117.720 60.530 119.525 ;
        RECT 61.370 117.720 62.830 119.525 ;
        RECT 63.670 117.720 65.130 119.525 ;
        RECT 65.970 117.720 67.430 119.525 ;
        RECT 68.270 117.720 69.730 119.525 ;
        RECT 70.570 117.720 72.030 119.525 ;
        RECT 72.870 117.720 74.330 119.525 ;
        RECT 75.170 117.720 76.630 119.525 ;
        RECT 77.470 117.720 78.930 119.525 ;
        RECT 79.770 117.720 81.230 119.525 ;
        RECT 82.070 117.720 83.530 119.525 ;
        RECT 84.370 117.720 85.830 119.525 ;
        RECT 86.670 117.720 88.130 119.525 ;
        RECT 0.100 5.255 88.680 117.720 ;
      LAYER met3 ;
        RECT 0.525 5.275 85.290 119.505 ;
      LAYER met4 ;
        RECT 1.215 114.880 85.265 119.505 ;
        RECT 1.215 55.935 14.190 114.880 ;
        RECT 16.590 55.935 24.060 114.880 ;
        RECT 26.460 55.935 33.930 114.880 ;
        RECT 36.330 55.935 43.800 114.880 ;
        RECT 46.200 55.935 53.670 114.880 ;
        RECT 56.070 55.935 63.540 114.880 ;
        RECT 65.940 55.935 73.410 114.880 ;
        RECT 75.810 55.935 85.265 114.880 ;
  END
END top
END LIBRARY

